
module fpu_add ( inq_op, inq_rnd_mode, inq_id, inq_fcc, inq_in1, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2, inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, 
        inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_add, add_dest_rdy, 
        fadd_clken_l, arst_l, grst_l, rclk, add_pipe_active, a1stg_step, 
        a6stg_fadd_in, add_id_out_in, a6stg_fcmpop, add_exc_out, a6stg_dbl_dst, 
        a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst, add_sign_out, 
        add_exp_out, add_frac_out, add_cc_out, add_fcc_out, se_add_exp, 
        se_add_frac, si, so );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [1:0] inq_fcc;
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  output [9:0] add_id_out_in;
  output [4:0] add_exc_out;
  output [10:0] add_exp_out;
  output [63:0] add_frac_out;
  output [1:0] add_cc_out;
  output [1:0] add_fcc_out;
  input inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0,
         inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0, inq_in2_53_32_neq_0,
         inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_add, add_dest_rdy,
         fadd_clken_l, arst_l, grst_l, rclk, se_add_exp, se_add_frac, si;
  output add_pipe_active, a1stg_step, a6stg_fadd_in, a6stg_fcmpop,
         a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst,
         add_sign_out, so;
  wire   a1stg_fsdtoix, a1stg_faddsubs, a1stg_fdtos, a3stg_fdtos_inv,
         \a4stg_shl_cnt[5] , \fpu_add_ctl/n941 , \fpu_add_ctl/n940 ,
         \fpu_add_ctl/n939 , \fpu_add_ctl/n938 , \fpu_add_ctl/n937 ,
         \fpu_add_ctl/n936 , \fpu_add_ctl/n470 , \fpu_add_ctl/n49 ,
         \fpu_add_ctl/n47 , \fpu_add_ctl/n338 , \fpu_add_ctl/n337 ,
         \fpu_add_ctl/n336 , \fpu_add_ctl/n335 , \fpu_add_ctl/n334 ,
         \fpu_add_ctl/n333 , \fpu_add_ctl/n332 , \fpu_add_ctl/n330 ,
         \fpu_add_ctl/n329 , \fpu_add_ctl/n328 , \fpu_add_ctl/n327 ,
         \fpu_add_ctl/n326 , \fpu_add_ctl/n325 , \fpu_add_ctl/n324 ,
         \fpu_add_ctl/n323 , \fpu_add_ctl/n322 , \fpu_add_ctl/n321 ,
         \fpu_add_ctl/n320 , \fpu_add_ctl/n319 , \fpu_add_ctl/n318 ,
         \fpu_add_ctl/n317 , \fpu_add_ctl/n316 , \fpu_add_ctl/n315 ,
         \fpu_add_ctl/n314 , \fpu_add_ctl/n313 , \fpu_add_ctl/n312 ,
         \fpu_add_ctl/n311 , \fpu_add_ctl/n310 , \fpu_add_ctl/n309 ,
         \fpu_add_ctl/n308 , \fpu_add_ctl/n307 , \fpu_add_ctl/n303 ,
         \fpu_add_ctl/n752 , \fpu_add_ctl/n751 , \fpu_add_ctl/n750 ,
         \fpu_add_ctl/n749 , \fpu_add_ctl/n748 , \fpu_add_ctl/n747 ,
         \fpu_add_ctl/n746 , \fpu_add_ctl/n745 , \fpu_add_ctl/n744 ,
         \fpu_add_ctl/n743 , \fpu_add_ctl/n742 , \fpu_add_ctl/n741 ,
         \fpu_add_ctl/n740 , \fpu_add_ctl/n739 , \fpu_add_ctl/n738 ,
         \fpu_add_ctl/n737 , \fpu_add_ctl/n736 , \fpu_add_ctl/n735 ,
         \fpu_add_ctl/n734 , \fpu_add_ctl/n733 , \fpu_add_ctl/n732 ,
         \fpu_add_ctl/n731 , \fpu_add_ctl/n730 , \fpu_add_ctl/n729 ,
         \fpu_add_ctl/n728 , \fpu_add_ctl/n727 , \fpu_add_ctl/n726 ,
         \fpu_add_ctl/n725 , \fpu_add_ctl/n724 , \fpu_add_ctl/n723 ,
         \fpu_add_ctl/n722 , \fpu_add_ctl/n721 , \fpu_add_ctl/n720 ,
         \fpu_add_ctl/n719 , \fpu_add_ctl/n718 , \fpu_add_ctl/n717 ,
         \fpu_add_ctl/n716 , \fpu_add_ctl/n715 , \fpu_add_ctl/n714 ,
         \fpu_add_ctl/n713 , \fpu_add_ctl/n712 , \fpu_add_ctl/n711 ,
         \fpu_add_ctl/n710 , \fpu_add_ctl/n709 , \fpu_add_ctl/n708 ,
         \fpu_add_ctl/n707 , \fpu_add_ctl/n706 , \fpu_add_ctl/n705 ,
         \fpu_add_ctl/n704 , \fpu_add_ctl/n703 , \fpu_add_ctl/n702 ,
         \fpu_add_ctl/n701 , \fpu_add_ctl/n700 , \fpu_add_ctl/n699 ,
         \fpu_add_ctl/n698 , \fpu_add_ctl/n697 , \fpu_add_ctl/n696 ,
         \fpu_add_ctl/n695 , \fpu_add_ctl/n694 , \fpu_add_ctl/n693 ,
         \fpu_add_ctl/n692 , \fpu_add_ctl/n691 , \fpu_add_ctl/n690 ,
         \fpu_add_ctl/n689 , \fpu_add_ctl/n688 , \fpu_add_ctl/n687 ,
         \fpu_add_ctl/n686 , \fpu_add_ctl/n685 , \fpu_add_ctl/n684 ,
         \fpu_add_ctl/n683 , \fpu_add_ctl/n682 , \fpu_add_ctl/n681 ,
         \fpu_add_ctl/n680 , \fpu_add_ctl/n679 , \fpu_add_ctl/n678 ,
         \fpu_add_ctl/n677 , \fpu_add_ctl/n676 , \fpu_add_ctl/n675 ,
         \fpu_add_ctl/n674 , \fpu_add_ctl/n673 , \fpu_add_ctl/n672 ,
         \fpu_add_ctl/n671 , \fpu_add_ctl/n670 , \fpu_add_ctl/n669 ,
         \fpu_add_ctl/n668 , \fpu_add_ctl/n667 , \fpu_add_ctl/n666 ,
         \fpu_add_ctl/n665 , \fpu_add_ctl/n664 , \fpu_add_ctl/n663 ,
         \fpu_add_ctl/n662 , \fpu_add_ctl/n661 , \fpu_add_ctl/n660 ,
         \fpu_add_ctl/n659 , \fpu_add_ctl/n658 , \fpu_add_ctl/n657 ,
         \fpu_add_ctl/n656 , \fpu_add_ctl/n655 , \fpu_add_ctl/n654 ,
         \fpu_add_ctl/n653 , \fpu_add_ctl/n652 , \fpu_add_ctl/n651 ,
         \fpu_add_ctl/n650 , \fpu_add_ctl/n649 , \fpu_add_ctl/n648 ,
         \fpu_add_ctl/n647 , \fpu_add_ctl/n646 , \fpu_add_ctl/n645 ,
         \fpu_add_ctl/n644 , \fpu_add_ctl/n643 , \fpu_add_ctl/n642 ,
         \fpu_add_ctl/n641 , \fpu_add_ctl/n640 , \fpu_add_ctl/n639 ,
         \fpu_add_ctl/n638 , \fpu_add_ctl/n637 , \fpu_add_ctl/n636 ,
         \fpu_add_ctl/n635 , \fpu_add_ctl/n634 , \fpu_add_ctl/n633 ,
         \fpu_add_ctl/n632 , \fpu_add_ctl/n631 , \fpu_add_ctl/n630 ,
         \fpu_add_ctl/n629 , \fpu_add_ctl/n628 , \fpu_add_ctl/n627 ,
         \fpu_add_ctl/n626 , \fpu_add_ctl/n625 , \fpu_add_ctl/n624 ,
         \fpu_add_ctl/n623 , \fpu_add_ctl/n622 , \fpu_add_ctl/n621 ,
         \fpu_add_ctl/n620 , \fpu_add_ctl/n619 , \fpu_add_ctl/n618 ,
         \fpu_add_ctl/n617 , \fpu_add_ctl/n616 , \fpu_add_ctl/n615 ,
         \fpu_add_ctl/n614 , \fpu_add_ctl/n613 , \fpu_add_ctl/n612 ,
         \fpu_add_ctl/n611 , \fpu_add_ctl/n610 , \fpu_add_ctl/n609 ,
         \fpu_add_ctl/n608 , \fpu_add_ctl/n607 , \fpu_add_ctl/n606 ,
         \fpu_add_ctl/n605 , \fpu_add_ctl/n604 , \fpu_add_ctl/n603 ,
         \fpu_add_ctl/n602 , \fpu_add_ctl/n601 , \fpu_add_ctl/n600 ,
         \fpu_add_ctl/n599 , \fpu_add_ctl/n598 , \fpu_add_ctl/n597 ,
         \fpu_add_ctl/n596 , \fpu_add_ctl/n595 , \fpu_add_ctl/n594 ,
         \fpu_add_ctl/n593 , \fpu_add_ctl/n592 , \fpu_add_ctl/n591 ,
         \fpu_add_ctl/n590 , \fpu_add_ctl/n589 , \fpu_add_ctl/n588 ,
         \fpu_add_ctl/n587 , \fpu_add_ctl/n586 , \fpu_add_ctl/n585 ,
         \fpu_add_ctl/n584 , \fpu_add_ctl/n583 , \fpu_add_ctl/n582 ,
         \fpu_add_ctl/n581 , \fpu_add_ctl/n580 , \fpu_add_ctl/n579 ,
         \fpu_add_ctl/n578 , \fpu_add_ctl/n577 , \fpu_add_ctl/n576 ,
         \fpu_add_ctl/n575 , \fpu_add_ctl/n574 , \fpu_add_ctl/n573 ,
         \fpu_add_ctl/n572 , \fpu_add_ctl/n571 , \fpu_add_ctl/n570 ,
         \fpu_add_ctl/n569 , \fpu_add_ctl/n568 , \fpu_add_ctl/n567 ,
         \fpu_add_ctl/n566 , \fpu_add_ctl/n565 , \fpu_add_ctl/n564 ,
         \fpu_add_ctl/n563 , \fpu_add_ctl/n562 , \fpu_add_ctl/n561 ,
         \fpu_add_ctl/n560 , \fpu_add_ctl/n559 , \fpu_add_ctl/n558 ,
         \fpu_add_ctl/n557 , \fpu_add_ctl/n556 , \fpu_add_ctl/n555 ,
         \fpu_add_ctl/n554 , \fpu_add_ctl/n553 , \fpu_add_ctl/n552 ,
         \fpu_add_ctl/n551 , \fpu_add_ctl/n550 , \fpu_add_ctl/n549 ,
         \fpu_add_ctl/n548 , \fpu_add_ctl/n547 , \fpu_add_ctl/n546 ,
         \fpu_add_ctl/n545 , \fpu_add_ctl/n544 , \fpu_add_ctl/n543 ,
         \fpu_add_ctl/n542 , \fpu_add_ctl/n541 , \fpu_add_ctl/n540 ,
         \fpu_add_ctl/n441 , \fpu_add_ctl/n426 , \fpu_add_ctl/n425 ,
         \fpu_add_ctl/n416 , \fpu_add_ctl/n269 , \fpu_add_ctl/n255 ,
         \fpu_add_ctl/n252 , \fpu_add_ctl/n210 , \fpu_add_ctl/n207 ,
         \fpu_add_ctl/n205 , \fpu_add_ctl/n203 , \fpu_add_ctl/n202 ,
         \fpu_add_ctl/n200 , \fpu_add_ctl/n196 , \fpu_add_ctl/n183 ,
         \fpu_add_ctl/n182 , \fpu_add_ctl/n177 , \fpu_add_ctl/n150 ,
         \fpu_add_ctl/n147 , \fpu_add_ctl/n144 , \fpu_add_ctl/n143 ,
         \fpu_add_ctl/n142 , \fpu_add_ctl/n141 , \fpu_add_ctl/n140 ,
         \fpu_add_ctl/n139 , \fpu_add_ctl/n138 , \fpu_add_ctl/n133 ,
         \fpu_add_ctl/n130 , \fpu_add_ctl/n129 , \fpu_add_ctl/n127 ,
         \fpu_add_ctl/n125 , \fpu_add_ctl/n124 , \fpu_add_ctl/n123 ,
         \fpu_add_ctl/n122 , \fpu_add_ctl/n121 , \fpu_add_ctl/n119 ,
         \fpu_add_ctl/n118 , \fpu_add_ctl/n117 , \fpu_add_ctl/n116 ,
         \fpu_add_ctl/n113 , \fpu_add_ctl/n110 , \fpu_add_ctl/n109 ,
         \fpu_add_ctl/n102 , \fpu_add_ctl/n101 , \fpu_add_ctl/n97 ,
         \fpu_add_ctl/n90 , \fpu_add_ctl/n89 , \fpu_add_ctl/n86 ,
         \fpu_add_ctl/n85 , \fpu_add_ctl/n79 , \fpu_add_ctl/n78 ,
         \fpu_add_ctl/n77 , \fpu_add_ctl/n66 , \fpu_add_ctl/n65 ,
         \fpu_add_ctl/n41 , \fpu_add_ctl/n40 , \fpu_add_ctl/n39 ,
         \fpu_add_ctl/n38 , \fpu_add_ctl/n37 , \fpu_add_ctl/n34 ,
         \fpu_add_ctl/n32 , \fpu_add_ctl/n31 , \fpu_add_ctl/n16 ,
         \fpu_add_ctl/n15 , \fpu_add_ctl/n14 , \fpu_add_ctl/n13 ,
         \fpu_add_ctl/n9 , \fpu_add_ctl/n7 , \fpu_add_ctl/n5 ,
         \fpu_add_ctl/n4 , \fpu_add_ctl/n3 , \fpu_add_ctl/n2 ,
         \fpu_add_ctl/n1 , \fpu_add_ctl/i_add_pipe_active/N7 ,
         \fpu_add_ctl/dffrl_add_ctl/N4 , \fpu_add_ctl/add_nx_out ,
         \fpu_add_ctl/add_of_out_tmp2 , \fpu_add_ctl/a3stg_a2_expadd_11 ,
         \fpu_add_ctl/a2stg_nan_in2 , \fpu_add_ctl/a2stg_in2_gt_in1_exp ,
         \fpu_add_ctl/add_id_out[9] , \fpu_add_ctl/add_id_out[8] ,
         \fpu_add_ctl/add_id_out[7] , \fpu_add_ctl/add_id_out[6] ,
         \fpu_add_ctl/add_id_out[5] , \fpu_add_ctl/add_id_out[4] ,
         \fpu_add_ctl/add_id_out[3] , \fpu_add_ctl/add_id_out[2] ,
         \fpu_add_ctl/add_id_out[1] , \fpu_add_ctl/add_id_out[0] ,
         \fpu_add_ctl/a3stg_id[2] , \fpu_add_ctl/a3stg_opdec_9_0[3] ,
         \fpu_add_ctl/a2stg_id[2] , \fpu_add_ctl/add_ctl_rst_l ,
         \fpu_add_exp_dp/n452 , \fpu_add_exp_dp/n451 , \fpu_add_exp_dp/n450 ,
         \fpu_add_exp_dp/n448 , \fpu_add_exp_dp/n447 , \fpu_add_exp_dp/n446 ,
         \fpu_add_exp_dp/n445 , \fpu_add_exp_dp/n444 , \fpu_add_exp_dp/n443 ,
         \fpu_add_exp_dp/n442 , \fpu_add_exp_dp/n441 , \fpu_add_exp_dp/n440 ,
         \fpu_add_exp_dp/n439 , \fpu_add_exp_dp/n438 , \fpu_add_exp_dp/n437 ,
         \fpu_add_exp_dp/n436 , \fpu_add_exp_dp/n435 , \fpu_add_exp_dp/n434 ,
         \fpu_add_exp_dp/n433 , \fpu_add_exp_dp/n432 , \fpu_add_exp_dp/n431 ,
         \fpu_add_exp_dp/n47 , \fpu_add_exp_dp/n45 , \fpu_add_exp_dp/n722 ,
         \fpu_add_exp_dp/n721 , \fpu_add_exp_dp/n720 , \fpu_add_exp_dp/n719 ,
         \fpu_add_exp_dp/n718 , \fpu_add_exp_dp/n717 , \fpu_add_exp_dp/n716 ,
         \fpu_add_exp_dp/n715 , \fpu_add_exp_dp/n714 , \fpu_add_exp_dp/n713 ,
         \fpu_add_exp_dp/n712 , \fpu_add_exp_dp/n711 , \fpu_add_exp_dp/n710 ,
         \fpu_add_exp_dp/n709 , \fpu_add_exp_dp/n708 , \fpu_add_exp_dp/n707 ,
         \fpu_add_exp_dp/n706 , \fpu_add_exp_dp/n705 , \fpu_add_exp_dp/n704 ,
         \fpu_add_exp_dp/n703 , \fpu_add_exp_dp/n702 , \fpu_add_exp_dp/n701 ,
         \fpu_add_exp_dp/n700 , \fpu_add_exp_dp/n699 , \fpu_add_exp_dp/n698 ,
         \fpu_add_exp_dp/n697 , \fpu_add_exp_dp/n696 , \fpu_add_exp_dp/n695 ,
         \fpu_add_exp_dp/n694 , \fpu_add_exp_dp/n693 , \fpu_add_exp_dp/n692 ,
         \fpu_add_exp_dp/n691 , \fpu_add_exp_dp/n690 , \fpu_add_exp_dp/n689 ,
         \fpu_add_exp_dp/n688 , \fpu_add_exp_dp/n687 , \fpu_add_exp_dp/n686 ,
         \fpu_add_exp_dp/n685 , \fpu_add_exp_dp/n684 , \fpu_add_exp_dp/n683 ,
         \fpu_add_exp_dp/n682 , \fpu_add_exp_dp/n681 , \fpu_add_exp_dp/n680 ,
         \fpu_add_exp_dp/n679 , \fpu_add_exp_dp/n678 , \fpu_add_exp_dp/n677 ,
         \fpu_add_exp_dp/n676 , \fpu_add_exp_dp/n675 , \fpu_add_exp_dp/n674 ,
         \fpu_add_exp_dp/n673 , \fpu_add_exp_dp/n672 , \fpu_add_exp_dp/n671 ,
         \fpu_add_exp_dp/n670 , \fpu_add_exp_dp/n669 , \fpu_add_exp_dp/n668 ,
         \fpu_add_exp_dp/n667 , \fpu_add_exp_dp/n666 , \fpu_add_exp_dp/n665 ,
         \fpu_add_exp_dp/n664 , \fpu_add_exp_dp/n663 , \fpu_add_exp_dp/n662 ,
         \fpu_add_exp_dp/n661 , \fpu_add_exp_dp/n660 , \fpu_add_exp_dp/n659 ,
         \fpu_add_exp_dp/n658 , \fpu_add_exp_dp/n657 , \fpu_add_exp_dp/n656 ,
         \fpu_add_exp_dp/n655 , \fpu_add_exp_dp/n654 , \fpu_add_exp_dp/n653 ,
         \fpu_add_exp_dp/n652 , \fpu_add_exp_dp/n651 , \fpu_add_exp_dp/n650 ,
         \fpu_add_exp_dp/n649 , \fpu_add_exp_dp/n648 , \fpu_add_exp_dp/n647 ,
         \fpu_add_exp_dp/n646 , \fpu_add_exp_dp/n645 , \fpu_add_exp_dp/n644 ,
         \fpu_add_exp_dp/n643 , \fpu_add_exp_dp/n642 , \fpu_add_exp_dp/n641 ,
         \fpu_add_exp_dp/n640 , \fpu_add_exp_dp/n639 , \fpu_add_exp_dp/n638 ,
         \fpu_add_exp_dp/n637 , \fpu_add_exp_dp/n636 , \fpu_add_exp_dp/n635 ,
         \fpu_add_exp_dp/n634 , \fpu_add_exp_dp/n633 , \fpu_add_exp_dp/n632 ,
         \fpu_add_exp_dp/n631 , \fpu_add_exp_dp/n630 , \fpu_add_exp_dp/n629 ,
         \fpu_add_exp_dp/n628 , \fpu_add_exp_dp/n627 , \fpu_add_exp_dp/n626 ,
         \fpu_add_exp_dp/n625 , \fpu_add_exp_dp/n624 , \fpu_add_exp_dp/n623 ,
         \fpu_add_exp_dp/n622 , \fpu_add_exp_dp/n621 , \fpu_add_exp_dp/n620 ,
         \fpu_add_exp_dp/n619 , \fpu_add_exp_dp/n618 , \fpu_add_exp_dp/n617 ,
         \fpu_add_exp_dp/n616 , \fpu_add_exp_dp/n615 , \fpu_add_exp_dp/n614 ,
         \fpu_add_exp_dp/n613 , \fpu_add_exp_dp/n612 , \fpu_add_exp_dp/n611 ,
         \fpu_add_exp_dp/n610 , \fpu_add_exp_dp/n609 , \fpu_add_exp_dp/n608 ,
         \fpu_add_exp_dp/n607 , \fpu_add_exp_dp/n606 , \fpu_add_exp_dp/n605 ,
         \fpu_add_exp_dp/n604 , \fpu_add_exp_dp/n603 , \fpu_add_exp_dp/n602 ,
         \fpu_add_exp_dp/n601 , \fpu_add_exp_dp/n600 , \fpu_add_exp_dp/n599 ,
         \fpu_add_exp_dp/n598 , \fpu_add_exp_dp/n597 , \fpu_add_exp_dp/n596 ,
         \fpu_add_exp_dp/n595 , \fpu_add_exp_dp/n594 , \fpu_add_exp_dp/n593 ,
         \fpu_add_exp_dp/n592 , \fpu_add_exp_dp/n591 , \fpu_add_exp_dp/n589 ,
         \fpu_add_exp_dp/n588 , \fpu_add_exp_dp/n587 , \fpu_add_exp_dp/n586 ,
         \fpu_add_exp_dp/n585 , \fpu_add_exp_dp/n584 , \fpu_add_exp_dp/n583 ,
         \fpu_add_exp_dp/n582 , \fpu_add_exp_dp/n581 , \fpu_add_exp_dp/n580 ,
         \fpu_add_exp_dp/n579 , \fpu_add_exp_dp/n578 , \fpu_add_exp_dp/n577 ,
         \fpu_add_exp_dp/n576 , \fpu_add_exp_dp/n575 , \fpu_add_exp_dp/n574 ,
         \fpu_add_exp_dp/n573 , \fpu_add_exp_dp/n572 , \fpu_add_exp_dp/n571 ,
         \fpu_add_exp_dp/n570 , \fpu_add_exp_dp/n569 , \fpu_add_exp_dp/n568 ,
         \fpu_add_exp_dp/n567 , \fpu_add_exp_dp/n566 , \fpu_add_exp_dp/n565 ,
         \fpu_add_exp_dp/n563 , \fpu_add_exp_dp/n562 , \fpu_add_exp_dp/n561 ,
         \fpu_add_exp_dp/n560 , \fpu_add_exp_dp/n559 , \fpu_add_exp_dp/n558 ,
         \fpu_add_exp_dp/n557 , \fpu_add_exp_dp/n556 , \fpu_add_exp_dp/n555 ,
         \fpu_add_exp_dp/n554 , \fpu_add_exp_dp/n553 , \fpu_add_exp_dp/n552 ,
         \fpu_add_exp_dp/n550 , \fpu_add_exp_dp/n549 , \fpu_add_exp_dp/n548 ,
         \fpu_add_exp_dp/n547 , \fpu_add_exp_dp/n546 , \fpu_add_exp_dp/n545 ,
         \fpu_add_exp_dp/n544 , \fpu_add_exp_dp/n543 , \fpu_add_exp_dp/n542 ,
         \fpu_add_exp_dp/n541 , \fpu_add_exp_dp/n540 , \fpu_add_exp_dp/n539 ,
         \fpu_add_exp_dp/n538 , \fpu_add_exp_dp/n537 , \fpu_add_exp_dp/n536 ,
         \fpu_add_exp_dp/n535 , \fpu_add_exp_dp/n534 , \fpu_add_exp_dp/n533 ,
         \fpu_add_exp_dp/n532 , \fpu_add_exp_dp/n531 , \fpu_add_exp_dp/n530 ,
         \fpu_add_exp_dp/n529 , \fpu_add_exp_dp/n528 , \fpu_add_exp_dp/n527 ,
         \fpu_add_exp_dp/n526 , \fpu_add_exp_dp/n525 , \fpu_add_exp_dp/n524 ,
         \fpu_add_exp_dp/n523 , \fpu_add_exp_dp/n522 , \fpu_add_exp_dp/n521 ,
         \fpu_add_exp_dp/n520 , \fpu_add_exp_dp/n519 , \fpu_add_exp_dp/n518 ,
         \fpu_add_exp_dp/n517 , \fpu_add_exp_dp/n516 , \fpu_add_exp_dp/n515 ,
         \fpu_add_exp_dp/n514 , \fpu_add_exp_dp/n513 , \fpu_add_exp_dp/n512 ,
         \fpu_add_exp_dp/n511 , \fpu_add_exp_dp/n510 , \fpu_add_exp_dp/n509 ,
         \fpu_add_exp_dp/n508 , \fpu_add_exp_dp/n507 , \fpu_add_exp_dp/n256 ,
         \fpu_add_exp_dp/n253 , \fpu_add_exp_dp/n252 , \fpu_add_exp_dp/n251 ,
         \fpu_add_exp_dp/n250 , \fpu_add_exp_dp/n249 , \fpu_add_exp_dp/n248 ,
         \fpu_add_exp_dp/n247 , \fpu_add_exp_dp/n246 , \fpu_add_exp_dp/n245 ,
         \fpu_add_exp_dp/n244 , \fpu_add_exp_dp/n243 , \fpu_add_exp_dp/n242 ,
         \fpu_add_exp_dp/n241 , \fpu_add_exp_dp/n240 , \fpu_add_exp_dp/n239 ,
         \fpu_add_exp_dp/n238 , \fpu_add_exp_dp/n237 , \fpu_add_exp_dp/n236 ,
         \fpu_add_exp_dp/n235 , \fpu_add_exp_dp/n234 , \fpu_add_exp_dp/n233 ,
         \fpu_add_exp_dp/n232 , \fpu_add_exp_dp/n231 , \fpu_add_exp_dp/n230 ,
         \fpu_add_exp_dp/n229 , \fpu_add_exp_dp/n228 , \fpu_add_exp_dp/n225 ,
         \fpu_add_exp_dp/n224 , \fpu_add_exp_dp/n222 , \fpu_add_exp_dp/n221 ,
         \fpu_add_exp_dp/n220 , \fpu_add_exp_dp/n219 , \fpu_add_exp_dp/n218 ,
         \fpu_add_exp_dp/n217 , \fpu_add_exp_dp/n216 , \fpu_add_exp_dp/n215 ,
         \fpu_add_exp_dp/n214 , \fpu_add_exp_dp/n213 , \fpu_add_exp_dp/n212 ,
         \fpu_add_exp_dp/n211 , \fpu_add_exp_dp/n210 , \fpu_add_exp_dp/n209 ,
         \fpu_add_exp_dp/n208 , \fpu_add_exp_dp/n207 , \fpu_add_exp_dp/n206 ,
         \fpu_add_exp_dp/n205 , \fpu_add_exp_dp/n204 , \fpu_add_exp_dp/n203 ,
         \fpu_add_exp_dp/n202 , \fpu_add_exp_dp/n201 , \fpu_add_exp_dp/n200 ,
         \fpu_add_exp_dp/n199 , \fpu_add_exp_dp/n198 , \fpu_add_exp_dp/n197 ,
         \fpu_add_exp_dp/n196 , \fpu_add_exp_dp/n195 , \fpu_add_exp_dp/n194 ,
         \fpu_add_exp_dp/n193 , \fpu_add_exp_dp/n192 , \fpu_add_exp_dp/n191 ,
         \fpu_add_exp_dp/n190 , \fpu_add_exp_dp/n189 , \fpu_add_exp_dp/n188 ,
         \fpu_add_exp_dp/n187 , \fpu_add_exp_dp/n186 , \fpu_add_exp_dp/n185 ,
         \fpu_add_exp_dp/n184 , \fpu_add_exp_dp/n183 , \fpu_add_exp_dp/n182 ,
         \fpu_add_exp_dp/n181 , \fpu_add_exp_dp/n180 , \fpu_add_exp_dp/n179 ,
         \fpu_add_exp_dp/n178 , \fpu_add_exp_dp/n177 , \fpu_add_exp_dp/n176 ,
         \fpu_add_exp_dp/n175 , \fpu_add_exp_dp/n174 , \fpu_add_exp_dp/n172 ,
         \fpu_add_exp_dp/n171 , \fpu_add_exp_dp/n170 , \fpu_add_exp_dp/n150 ,
         \fpu_add_exp_dp/n149 , \fpu_add_exp_dp/n147 , \fpu_add_exp_dp/n146 ,
         \fpu_add_exp_dp/n145 , \fpu_add_exp_dp/n144 , \fpu_add_exp_dp/n143 ,
         \fpu_add_exp_dp/n142 , \fpu_add_exp_dp/n141 , \fpu_add_exp_dp/n137 ,
         \fpu_add_exp_dp/n136 , \fpu_add_exp_dp/n135 , \fpu_add_exp_dp/n134 ,
         \fpu_add_exp_dp/n133 , \fpu_add_exp_dp/n132 , \fpu_add_exp_dp/n131 ,
         \fpu_add_exp_dp/n130 , \fpu_add_exp_dp/n129 , \fpu_add_exp_dp/n128 ,
         \fpu_add_exp_dp/n127 , \fpu_add_exp_dp/n126 , \fpu_add_exp_dp/n125 ,
         \fpu_add_exp_dp/n124 , \fpu_add_exp_dp/n122 , \fpu_add_exp_dp/n121 ,
         \fpu_add_exp_dp/n120 , \fpu_add_exp_dp/n119 , \fpu_add_exp_dp/n118 ,
         \fpu_add_exp_dp/n117 , \fpu_add_exp_dp/n116 , \fpu_add_exp_dp/n115 ,
         \fpu_add_exp_dp/n114 , \fpu_add_exp_dp/n113 , \fpu_add_exp_dp/n112 ,
         \fpu_add_exp_dp/n111 , \fpu_add_exp_dp/n109 , \fpu_add_exp_dp/n108 ,
         \fpu_add_exp_dp/n107 , \fpu_add_exp_dp/n106 , \fpu_add_exp_dp/n105 ,
         \fpu_add_exp_dp/n104 , \fpu_add_exp_dp/n103 , \fpu_add_exp_dp/n102 ,
         \fpu_add_exp_dp/n101 , \fpu_add_exp_dp/n100 , \fpu_add_exp_dp/n99 ,
         \fpu_add_exp_dp/n98 , \fpu_add_exp_dp/n96 , \fpu_add_exp_dp/n95 ,
         \fpu_add_exp_dp/n94 , \fpu_add_exp_dp/n93 , \fpu_add_exp_dp/n92 ,
         \fpu_add_exp_dp/n91 , \fpu_add_exp_dp/n90 , \fpu_add_exp_dp/n89 ,
         \fpu_add_exp_dp/n88 , \fpu_add_exp_dp/n87 , \fpu_add_exp_dp/n86 ,
         \fpu_add_exp_dp/n85 , \fpu_add_exp_dp/n83 , \fpu_add_exp_dp/n82 ,
         \fpu_add_exp_dp/n81 , \fpu_add_exp_dp/n80 , \fpu_add_exp_dp/n79 ,
         \fpu_add_exp_dp/n78 , \fpu_add_exp_dp/n77 , \fpu_add_exp_dp/n76 ,
         \fpu_add_exp_dp/n75 , \fpu_add_exp_dp/n74 , \fpu_add_exp_dp/n73 ,
         \fpu_add_exp_dp/n72 , \fpu_add_exp_dp/n71 , \fpu_add_exp_dp/n70 ,
         \fpu_add_exp_dp/n69 , \fpu_add_exp_dp/n68 , \fpu_add_exp_dp/n67 ,
         \fpu_add_exp_dp/n66 , \fpu_add_exp_dp/n65 , \fpu_add_exp_dp/n64 ,
         \fpu_add_exp_dp/n63 , \fpu_add_exp_dp/n62 , \fpu_add_exp_dp/n61 ,
         \fpu_add_exp_dp/n60 , \fpu_add_exp_dp/n57 , \fpu_add_exp_dp/n50 ,
         \fpu_add_exp_dp/n48 , \fpu_add_exp_dp/n46 , \fpu_add_exp_dp/n22 ,
         \fpu_add_exp_dp/n21 , \fpu_add_exp_dp/n20 , \fpu_add_exp_dp/n19 ,
         \fpu_add_exp_dp/n18 , \fpu_add_exp_dp/n17 , \fpu_add_exp_dp/n16 ,
         \fpu_add_exp_dp/n15 , \fpu_add_exp_dp/n14 , \fpu_add_exp_dp/n13 ,
         \fpu_add_exp_dp/n12 , \fpu_add_exp_dp/n11 , \fpu_add_exp_dp/n10 ,
         \fpu_add_exp_dp/n9 , \fpu_add_exp_dp/n8 , \fpu_add_exp_dp/n7 ,
         \fpu_add_exp_dp/n6 , \fpu_add_exp_dp/n5 , \fpu_add_exp_dp/n4 ,
         \fpu_add_exp_dp/n3 , \fpu_add_exp_dp/n2 , \fpu_add_exp_dp/n1 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N3 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N4 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N5 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N6 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N7 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N8 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N9 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N10 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N11 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N12 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N13 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre4/N14 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N3 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N4 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N5 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N6 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N7 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N8 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N9 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N10 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N11 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N12 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N13 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre2/N14 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N3 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N4 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N5 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N6 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N7 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N8 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N9 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N10 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N11 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N12 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N13 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre3/N14 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N3 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N4 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N5 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N6 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N7 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N8 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N9 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N10 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N11 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N12 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N13 ,
         \fpu_add_exp_dp/i_a4stg_exp_pre1/N14 ,
         \fpu_add_exp_dp/ckbuf_add_exp_dp/N1 ,
         \fpu_add_exp_dp/ckbuf_add_exp_dp/clken ,
         \fpu_add_exp_dp/add_exp_out3[10] , \fpu_add_exp_dp/add_exp_out3[9] ,
         \fpu_add_exp_dp/add_exp_out3[8] , \fpu_add_exp_dp/add_exp_out3[7] ,
         \fpu_add_exp_dp/add_exp_out3[6] , \fpu_add_exp_dp/add_exp_out3[5] ,
         \fpu_add_exp_dp/add_exp_out3[4] , \fpu_add_exp_dp/add_exp_out3[3] ,
         \fpu_add_exp_dp/add_exp_out3[2] , \fpu_add_exp_dp/add_exp_out3[1] ,
         \fpu_add_exp_dp/add_exp_out3[0] , \fpu_add_exp_dp/a4stg_exp2[11] ,
         \fpu_add_exp_dp/a4stg_exp2[9] , \fpu_add_exp_dp/a4stg_exp2[8] ,
         \fpu_add_exp_dp/a4stg_exp2[7] , \fpu_add_exp_dp/a4stg_exp2[4] ,
         \fpu_add_exp_dp/a4stg_exp2[3] , \fpu_add_exp_dp/a4stg_exp2[2] ,
         \fpu_add_exp_dp/a4stg_exp2[0] , \fpu_add_exp_dp/a4stg_exp_pre4[11] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[10] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[9] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[8] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[7] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[6] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[5] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[4] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[3] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[2] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[1] ,
         \fpu_add_exp_dp/a4stg_exp_pre4[0] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[11] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[10] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[9] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[8] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[7] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[6] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[5] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[4] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[3] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[2] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[1] ,
         \fpu_add_exp_dp/a4stg_exp_pre2[0] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[11] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[10] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[9] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[8] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[7] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[6] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[5] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[4] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[3] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[2] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[1] ,
         \fpu_add_exp_dp/a4stg_exp_pre3[0] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[11] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[10] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[9] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[8] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[7] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[6] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[5] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[4] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[3] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[2] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[1] ,
         \fpu_add_exp_dp/a4stg_exp_pre1[0] ,
         \fpu_add_exp_dp/a1stg_expadd3_in2[10] ,
         \fpu_add_exp_dp/a1stg_in2a[59] , \fpu_add_exp_dp/a1stg_in2a[58] ,
         \fpu_add_exp_dp/a1stg_in2a[57] , \fpu_add_exp_dp/a1stg_in2a[56] ,
         \fpu_add_exp_dp/a1stg_in2a[55] , \fpu_add_exp_dp/a1stg_in2a[54] ,
         \fpu_add_exp_dp/a1stg_in2a[53] , \fpu_add_exp_dp/a1stg_in2a[52] ,
         \fpu_add_frac_dp/n5644 , \fpu_add_frac_dp/n5643 ,
         \fpu_add_frac_dp/n5642 , \fpu_add_frac_dp/n5641 ,
         \fpu_add_frac_dp/n5640 , \fpu_add_frac_dp/n5635 ,
         \fpu_add_frac_dp/n5634 , \fpu_add_frac_dp/n5633 ,
         \fpu_add_frac_dp/n5632 , \fpu_add_frac_dp/n5631 ,
         \fpu_add_frac_dp/n5630 , \fpu_add_frac_dp/n5629 ,
         \fpu_add_frac_dp/n5627 , \fpu_add_frac_dp/n5626 ,
         \fpu_add_frac_dp/n5625 , \fpu_add_frac_dp/n5624 ,
         \fpu_add_frac_dp/n5623 , \fpu_add_frac_dp/n5622 ,
         \fpu_add_frac_dp/n5621 , \fpu_add_frac_dp/n5620 ,
         \fpu_add_frac_dp/n5619 , \fpu_add_frac_dp/n5618 ,
         \fpu_add_frac_dp/n5617 , \fpu_add_frac_dp/n5616 ,
         \fpu_add_frac_dp/n5614 , \fpu_add_frac_dp/n5613 ,
         \fpu_add_frac_dp/n5612 , \fpu_add_frac_dp/n5611 ,
         \fpu_add_frac_dp/n5610 , \fpu_add_frac_dp/n5609 ,
         \fpu_add_frac_dp/n5608 , \fpu_add_frac_dp/n5605 ,
         \fpu_add_frac_dp/n2189 , \fpu_add_frac_dp/n1574 ,
         \fpu_add_frac_dp/n1573 , \fpu_add_frac_dp/n1572 ,
         \fpu_add_frac_dp/n1571 , \fpu_add_frac_dp/n1570 ,
         \fpu_add_frac_dp/n1569 , \fpu_add_frac_dp/n1568 ,
         \fpu_add_frac_dp/n1567 , \fpu_add_frac_dp/n1566 ,
         \fpu_add_frac_dp/n1565 , \fpu_add_frac_dp/n1564 ,
         \fpu_add_frac_dp/n1563 , \fpu_add_frac_dp/n1562 ,
         \fpu_add_frac_dp/n1561 , \fpu_add_frac_dp/n1560 ,
         \fpu_add_frac_dp/n1559 , \fpu_add_frac_dp/n1558 ,
         \fpu_add_frac_dp/n1557 , \fpu_add_frac_dp/n1556 ,
         \fpu_add_frac_dp/n1555 , \fpu_add_frac_dp/n1554 ,
         \fpu_add_frac_dp/n1553 , \fpu_add_frac_dp/n1552 ,
         \fpu_add_frac_dp/n1551 , \fpu_add_frac_dp/n1550 ,
         \fpu_add_frac_dp/n1549 , \fpu_add_frac_dp/n1548 ,
         \fpu_add_frac_dp/n1547 , \fpu_add_frac_dp/n1546 ,
         \fpu_add_frac_dp/n1545 , \fpu_add_frac_dp/n1544 ,
         \fpu_add_frac_dp/n1543 , \fpu_add_frac_dp/n1542 ,
         \fpu_add_frac_dp/n1541 , \fpu_add_frac_dp/n1540 ,
         \fpu_add_frac_dp/n1539 , \fpu_add_frac_dp/n1538 ,
         \fpu_add_frac_dp/n1537 , \fpu_add_frac_dp/n1536 ,
         \fpu_add_frac_dp/n1535 , \fpu_add_frac_dp/n1534 ,
         \fpu_add_frac_dp/n1533 , \fpu_add_frac_dp/n1532 ,
         \fpu_add_frac_dp/n1531 , \fpu_add_frac_dp/n1530 ,
         \fpu_add_frac_dp/n1529 , \fpu_add_frac_dp/n1528 ,
         \fpu_add_frac_dp/n1527 , \fpu_add_frac_dp/n1526 ,
         \fpu_add_frac_dp/n1525 , \fpu_add_frac_dp/n1524 ,
         \fpu_add_frac_dp/n1523 , \fpu_add_frac_dp/n1522 ,
         \fpu_add_frac_dp/n1521 , \fpu_add_frac_dp/n1520 ,
         \fpu_add_frac_dp/n1519 , \fpu_add_frac_dp/n1518 ,
         \fpu_add_frac_dp/n1517 , \fpu_add_frac_dp/n1516 ,
         \fpu_add_frac_dp/n1515 , \fpu_add_frac_dp/n1509 ,
         \fpu_add_frac_dp/n2544 , \fpu_add_frac_dp/n2543 ,
         \fpu_add_frac_dp/n2540 , \fpu_add_frac_dp/n2539 ,
         \fpu_add_frac_dp/n2538 , \fpu_add_frac_dp/n2537 ,
         \fpu_add_frac_dp/n2536 , \fpu_add_frac_dp/n2535 ,
         \fpu_add_frac_dp/n2534 , \fpu_add_frac_dp/n2533 ,
         \fpu_add_frac_dp/n2532 , \fpu_add_frac_dp/n2531 ,
         \fpu_add_frac_dp/n2530 , \fpu_add_frac_dp/n2529 ,
         \fpu_add_frac_dp/n2528 , \fpu_add_frac_dp/n2527 ,
         \fpu_add_frac_dp/n2526 , \fpu_add_frac_dp/n2525 ,
         \fpu_add_frac_dp/n2524 , \fpu_add_frac_dp/n2523 ,
         \fpu_add_frac_dp/n2522 , \fpu_add_frac_dp/n2521 ,
         \fpu_add_frac_dp/n2520 , \fpu_add_frac_dp/n2519 ,
         \fpu_add_frac_dp/n2518 , \fpu_add_frac_dp/n2517 ,
         \fpu_add_frac_dp/n2516 , \fpu_add_frac_dp/n2515 ,
         \fpu_add_frac_dp/n2514 , \fpu_add_frac_dp/n2513 ,
         \fpu_add_frac_dp/n2512 , \fpu_add_frac_dp/n2511 ,
         \fpu_add_frac_dp/n2510 , \fpu_add_frac_dp/n2509 ,
         \fpu_add_frac_dp/n2508 , \fpu_add_frac_dp/n2507 ,
         \fpu_add_frac_dp/n2506 , \fpu_add_frac_dp/n2505 ,
         \fpu_add_frac_dp/n2504 , \fpu_add_frac_dp/n2503 ,
         \fpu_add_frac_dp/n2502 , \fpu_add_frac_dp/n2501 ,
         \fpu_add_frac_dp/n2500 , \fpu_add_frac_dp/n2499 ,
         \fpu_add_frac_dp/n2498 , \fpu_add_frac_dp/n2497 ,
         \fpu_add_frac_dp/n2496 , \fpu_add_frac_dp/n2495 ,
         \fpu_add_frac_dp/n2494 , \fpu_add_frac_dp/n2493 ,
         \fpu_add_frac_dp/n2492 , \fpu_add_frac_dp/n2491 ,
         \fpu_add_frac_dp/n2490 , \fpu_add_frac_dp/n2489 ,
         \fpu_add_frac_dp/n2488 , \fpu_add_frac_dp/n2487 ,
         \fpu_add_frac_dp/n2486 , \fpu_add_frac_dp/n2485 ,
         \fpu_add_frac_dp/n2484 , \fpu_add_frac_dp/n2483 ,
         \fpu_add_frac_dp/n2482 , \fpu_add_frac_dp/n2481 ,
         \fpu_add_frac_dp/n2480 , \fpu_add_frac_dp/n2479 ,
         \fpu_add_frac_dp/n2478 , \fpu_add_frac_dp/n2477 ,
         \fpu_add_frac_dp/n2476 , \fpu_add_frac_dp/n2475 ,
         \fpu_add_frac_dp/n2474 , \fpu_add_frac_dp/n2473 ,
         \fpu_add_frac_dp/n2472 , \fpu_add_frac_dp/n2471 ,
         \fpu_add_frac_dp/n2470 , \fpu_add_frac_dp/n2469 ,
         \fpu_add_frac_dp/n2468 , \fpu_add_frac_dp/n2467 ,
         \fpu_add_frac_dp/n2466 , \fpu_add_frac_dp/n2465 ,
         \fpu_add_frac_dp/n2462 , \fpu_add_frac_dp/n2460 ,
         \fpu_add_frac_dp/n2459 , \fpu_add_frac_dp/n2458 ,
         \fpu_add_frac_dp/n2457 , \fpu_add_frac_dp/n2455 ,
         \fpu_add_frac_dp/n2454 , \fpu_add_frac_dp/n2453 ,
         \fpu_add_frac_dp/n2452 , \fpu_add_frac_dp/n2449 ,
         \fpu_add_frac_dp/n2448 , \fpu_add_frac_dp/n2447 ,
         \fpu_add_frac_dp/n2446 , \fpu_add_frac_dp/n2445 ,
         \fpu_add_frac_dp/n2444 , \fpu_add_frac_dp/n2442 ,
         \fpu_add_frac_dp/n2441 , \fpu_add_frac_dp/n2440 ,
         \fpu_add_frac_dp/n2439 , \fpu_add_frac_dp/n2438 ,
         \fpu_add_frac_dp/n2437 , \fpu_add_frac_dp/n2436 ,
         \fpu_add_frac_dp/n2435 , \fpu_add_frac_dp/n2434 ,
         \fpu_add_frac_dp/n2433 , \fpu_add_frac_dp/n2432 ,
         \fpu_add_frac_dp/n2431 , \fpu_add_frac_dp/n2430 ,
         \fpu_add_frac_dp/n2429 , \fpu_add_frac_dp/n2428 ,
         \fpu_add_frac_dp/n2427 , \fpu_add_frac_dp/n2426 ,
         \fpu_add_frac_dp/n2425 , \fpu_add_frac_dp/n2424 ,
         \fpu_add_frac_dp/n2423 , \fpu_add_frac_dp/n2422 ,
         \fpu_add_frac_dp/n2421 , \fpu_add_frac_dp/n2420 ,
         \fpu_add_frac_dp/n2419 , \fpu_add_frac_dp/n2418 ,
         \fpu_add_frac_dp/n2417 , \fpu_add_frac_dp/n2416 ,
         \fpu_add_frac_dp/n2415 , \fpu_add_frac_dp/n2414 ,
         \fpu_add_frac_dp/n2413 , \fpu_add_frac_dp/n2412 ,
         \fpu_add_frac_dp/n2411 , \fpu_add_frac_dp/n2410 ,
         \fpu_add_frac_dp/n2409 , \fpu_add_frac_dp/n2408 ,
         \fpu_add_frac_dp/n2407 , \fpu_add_frac_dp/n2406 ,
         \fpu_add_frac_dp/n2405 , \fpu_add_frac_dp/n2404 ,
         \fpu_add_frac_dp/n2403 , \fpu_add_frac_dp/n2402 ,
         \fpu_add_frac_dp/n2401 , \fpu_add_frac_dp/n2400 ,
         \fpu_add_frac_dp/n2399 , \fpu_add_frac_dp/n2398 ,
         \fpu_add_frac_dp/n2397 , \fpu_add_frac_dp/n2396 ,
         \fpu_add_frac_dp/n2395 , \fpu_add_frac_dp/n2394 ,
         \fpu_add_frac_dp/n2393 , \fpu_add_frac_dp/n2392 ,
         \fpu_add_frac_dp/n2391 , \fpu_add_frac_dp/n2390 ,
         \fpu_add_frac_dp/n2389 , \fpu_add_frac_dp/n2388 ,
         \fpu_add_frac_dp/n2387 , \fpu_add_frac_dp/n2386 ,
         \fpu_add_frac_dp/n2385 , \fpu_add_frac_dp/n2384 ,
         \fpu_add_frac_dp/n2382 , \fpu_add_frac_dp/n2381 ,
         \fpu_add_frac_dp/n2380 , \fpu_add_frac_dp/n2379 ,
         \fpu_add_frac_dp/n2378 , \fpu_add_frac_dp/n2377 ,
         \fpu_add_frac_dp/n2376 , \fpu_add_frac_dp/n2375 ,
         \fpu_add_frac_dp/n2374 , \fpu_add_frac_dp/n2373 ,
         \fpu_add_frac_dp/n2372 , \fpu_add_frac_dp/n2370 ,
         \fpu_add_frac_dp/n2369 , \fpu_add_frac_dp/n2368 ,
         \fpu_add_frac_dp/n2367 , \fpu_add_frac_dp/n2366 ,
         \fpu_add_frac_dp/n2365 , \fpu_add_frac_dp/n2364 ,
         \fpu_add_frac_dp/n2363 , \fpu_add_frac_dp/n2362 ,
         \fpu_add_frac_dp/n2361 , \fpu_add_frac_dp/n2360 ,
         \fpu_add_frac_dp/n2359 , \fpu_add_frac_dp/n2358 ,
         \fpu_add_frac_dp/n2357 , \fpu_add_frac_dp/n2356 ,
         \fpu_add_frac_dp/n2355 , \fpu_add_frac_dp/n2354 ,
         \fpu_add_frac_dp/n2353 , \fpu_add_frac_dp/n2352 ,
         \fpu_add_frac_dp/n2351 , \fpu_add_frac_dp/n2350 ,
         \fpu_add_frac_dp/n2349 , \fpu_add_frac_dp/n2348 ,
         \fpu_add_frac_dp/n2347 , \fpu_add_frac_dp/n2346 ,
         \fpu_add_frac_dp/n2345 , \fpu_add_frac_dp/n2344 ,
         \fpu_add_frac_dp/n2343 , \fpu_add_frac_dp/n2342 ,
         \fpu_add_frac_dp/n2341 , \fpu_add_frac_dp/n2340 ,
         \fpu_add_frac_dp/n2339 , \fpu_add_frac_dp/n2338 ,
         \fpu_add_frac_dp/n2337 , \fpu_add_frac_dp/n2336 ,
         \fpu_add_frac_dp/n2335 , \fpu_add_frac_dp/n2334 ,
         \fpu_add_frac_dp/n2333 , \fpu_add_frac_dp/n2332 ,
         \fpu_add_frac_dp/n2331 , \fpu_add_frac_dp/n2330 ,
         \fpu_add_frac_dp/n2325 , \fpu_add_frac_dp/n2322 ,
         \fpu_add_frac_dp/n2320 , \fpu_add_frac_dp/n2317 ,
         \fpu_add_frac_dp/n2316 , \fpu_add_frac_dp/n2314 ,
         \fpu_add_frac_dp/n2313 , \fpu_add_frac_dp/n2310 ,
         \fpu_add_frac_dp/n2309 , \fpu_add_frac_dp/n2308 ,
         \fpu_add_frac_dp/n2307 , \fpu_add_frac_dp/n2306 ,
         \fpu_add_frac_dp/n2305 , \fpu_add_frac_dp/n2304 ,
         \fpu_add_frac_dp/n2303 , \fpu_add_frac_dp/n2302 ,
         \fpu_add_frac_dp/n2301 , \fpu_add_frac_dp/n2300 ,
         \fpu_add_frac_dp/n2299 , \fpu_add_frac_dp/n2298 ,
         \fpu_add_frac_dp/n2297 , \fpu_add_frac_dp/n2296 ,
         \fpu_add_frac_dp/n2295 , \fpu_add_frac_dp/n2294 ,
         \fpu_add_frac_dp/n2293 , \fpu_add_frac_dp/n2292 ,
         \fpu_add_frac_dp/n2291 , \fpu_add_frac_dp/n2290 ,
         \fpu_add_frac_dp/n2289 , \fpu_add_frac_dp/n2288 ,
         \fpu_add_frac_dp/n2287 , \fpu_add_frac_dp/n2285 ,
         \fpu_add_frac_dp/n2282 , \fpu_add_frac_dp/n2281 ,
         \fpu_add_frac_dp/n2280 , \fpu_add_frac_dp/n2279 ,
         \fpu_add_frac_dp/n2278 , \fpu_add_frac_dp/n2277 ,
         \fpu_add_frac_dp/n2276 , \fpu_add_frac_dp/n2275 ,
         \fpu_add_frac_dp/n2274 , \fpu_add_frac_dp/n2273 ,
         \fpu_add_frac_dp/n2272 , \fpu_add_frac_dp/n2271 ,
         \fpu_add_frac_dp/n2270 , \fpu_add_frac_dp/n2269 ,
         \fpu_add_frac_dp/n2262 , \fpu_add_frac_dp/n4285 ,
         \fpu_add_frac_dp/n4284 , \fpu_add_frac_dp/n4283 ,
         \fpu_add_frac_dp/n4282 , \fpu_add_frac_dp/n4281 ,
         \fpu_add_frac_dp/n4280 , \fpu_add_frac_dp/n4279 ,
         \fpu_add_frac_dp/n4278 , \fpu_add_frac_dp/n4277 ,
         \fpu_add_frac_dp/n4276 , \fpu_add_frac_dp/n4275 ,
         \fpu_add_frac_dp/n4274 , \fpu_add_frac_dp/n4273 ,
         \fpu_add_frac_dp/n4272 , \fpu_add_frac_dp/n4271 ,
         \fpu_add_frac_dp/n4270 , \fpu_add_frac_dp/n4269 ,
         \fpu_add_frac_dp/n4268 , \fpu_add_frac_dp/n4267 ,
         \fpu_add_frac_dp/n4266 , \fpu_add_frac_dp/n4265 ,
         \fpu_add_frac_dp/n4264 , \fpu_add_frac_dp/n4263 ,
         \fpu_add_frac_dp/n4262 , \fpu_add_frac_dp/n4261 ,
         \fpu_add_frac_dp/n4260 , \fpu_add_frac_dp/n4259 ,
         \fpu_add_frac_dp/n4258 , \fpu_add_frac_dp/n4257 ,
         \fpu_add_frac_dp/n4256 , \fpu_add_frac_dp/n4255 ,
         \fpu_add_frac_dp/n4254 , \fpu_add_frac_dp/n4253 ,
         \fpu_add_frac_dp/n4252 , \fpu_add_frac_dp/n4251 ,
         \fpu_add_frac_dp/n4250 , \fpu_add_frac_dp/n4249 ,
         \fpu_add_frac_dp/n4248 , \fpu_add_frac_dp/n4247 ,
         \fpu_add_frac_dp/n4246 , \fpu_add_frac_dp/n4245 ,
         \fpu_add_frac_dp/n4244 , \fpu_add_frac_dp/n4243 ,
         \fpu_add_frac_dp/n4242 , \fpu_add_frac_dp/n4241 ,
         \fpu_add_frac_dp/n4240 , \fpu_add_frac_dp/n4239 ,
         \fpu_add_frac_dp/n4238 , \fpu_add_frac_dp/n4237 ,
         \fpu_add_frac_dp/n4236 , \fpu_add_frac_dp/n4235 ,
         \fpu_add_frac_dp/n4234 , \fpu_add_frac_dp/n4233 ,
         \fpu_add_frac_dp/n4232 , \fpu_add_frac_dp/n4231 ,
         \fpu_add_frac_dp/n4230 , \fpu_add_frac_dp/n4229 ,
         \fpu_add_frac_dp/n4228 , \fpu_add_frac_dp/n4227 ,
         \fpu_add_frac_dp/n4226 , \fpu_add_frac_dp/n4225 ,
         \fpu_add_frac_dp/n4224 , \fpu_add_frac_dp/n4223 ,
         \fpu_add_frac_dp/n4222 , \fpu_add_frac_dp/n4221 ,
         \fpu_add_frac_dp/n4220 , \fpu_add_frac_dp/n4219 ,
         \fpu_add_frac_dp/n4218 , \fpu_add_frac_dp/n4217 ,
         \fpu_add_frac_dp/n4216 , \fpu_add_frac_dp/n4215 ,
         \fpu_add_frac_dp/n4214 , \fpu_add_frac_dp/n4213 ,
         \fpu_add_frac_dp/n4212 , \fpu_add_frac_dp/n4211 ,
         \fpu_add_frac_dp/n4210 , \fpu_add_frac_dp/n4209 ,
         \fpu_add_frac_dp/n4208 , \fpu_add_frac_dp/n4207 ,
         \fpu_add_frac_dp/n4206 , \fpu_add_frac_dp/n4205 ,
         \fpu_add_frac_dp/n4204 , \fpu_add_frac_dp/n4203 ,
         \fpu_add_frac_dp/n4202 , \fpu_add_frac_dp/n4201 ,
         \fpu_add_frac_dp/n4200 , \fpu_add_frac_dp/n4199 ,
         \fpu_add_frac_dp/n4198 , \fpu_add_frac_dp/n4197 ,
         \fpu_add_frac_dp/n4196 , \fpu_add_frac_dp/n4195 ,
         \fpu_add_frac_dp/n4194 , \fpu_add_frac_dp/n4193 ,
         \fpu_add_frac_dp/n4192 , \fpu_add_frac_dp/n4191 ,
         \fpu_add_frac_dp/n4190 , \fpu_add_frac_dp/n4189 ,
         \fpu_add_frac_dp/n4188 , \fpu_add_frac_dp/n4187 ,
         \fpu_add_frac_dp/n4186 , \fpu_add_frac_dp/n4185 ,
         \fpu_add_frac_dp/n4184 , \fpu_add_frac_dp/n4183 ,
         \fpu_add_frac_dp/n4182 , \fpu_add_frac_dp/n4181 ,
         \fpu_add_frac_dp/n4180 , \fpu_add_frac_dp/n4179 ,
         \fpu_add_frac_dp/n4178 , \fpu_add_frac_dp/n4177 ,
         \fpu_add_frac_dp/n4176 , \fpu_add_frac_dp/n4175 ,
         \fpu_add_frac_dp/n4174 , \fpu_add_frac_dp/n4173 ,
         \fpu_add_frac_dp/n4172 , \fpu_add_frac_dp/n4171 ,
         \fpu_add_frac_dp/n4170 , \fpu_add_frac_dp/n4169 ,
         \fpu_add_frac_dp/n4168 , \fpu_add_frac_dp/n4167 ,
         \fpu_add_frac_dp/n4166 , \fpu_add_frac_dp/n4165 ,
         \fpu_add_frac_dp/n4164 , \fpu_add_frac_dp/n4163 ,
         \fpu_add_frac_dp/n4162 , \fpu_add_frac_dp/n4161 ,
         \fpu_add_frac_dp/n4160 , \fpu_add_frac_dp/n4159 ,
         \fpu_add_frac_dp/n4158 , \fpu_add_frac_dp/n4157 ,
         \fpu_add_frac_dp/n4156 , \fpu_add_frac_dp/n4155 ,
         \fpu_add_frac_dp/n4154 , \fpu_add_frac_dp/n4153 ,
         \fpu_add_frac_dp/n4152 , \fpu_add_frac_dp/n4151 ,
         \fpu_add_frac_dp/n4150 , \fpu_add_frac_dp/n4149 ,
         \fpu_add_frac_dp/n4148 , \fpu_add_frac_dp/n4147 ,
         \fpu_add_frac_dp/n4146 , \fpu_add_frac_dp/n4145 ,
         \fpu_add_frac_dp/n4144 , \fpu_add_frac_dp/n4143 ,
         \fpu_add_frac_dp/n4142 , \fpu_add_frac_dp/n4141 ,
         \fpu_add_frac_dp/n4140 , \fpu_add_frac_dp/n4139 ,
         \fpu_add_frac_dp/n4138 , \fpu_add_frac_dp/n4137 ,
         \fpu_add_frac_dp/n4136 , \fpu_add_frac_dp/n4135 ,
         \fpu_add_frac_dp/n4134 , \fpu_add_frac_dp/n4133 ,
         \fpu_add_frac_dp/n4132 , \fpu_add_frac_dp/n4131 ,
         \fpu_add_frac_dp/n4130 , \fpu_add_frac_dp/n4129 ,
         \fpu_add_frac_dp/n4128 , \fpu_add_frac_dp/n4127 ,
         \fpu_add_frac_dp/n4126 , \fpu_add_frac_dp/n4125 ,
         \fpu_add_frac_dp/n4124 , \fpu_add_frac_dp/n4123 ,
         \fpu_add_frac_dp/n4122 , \fpu_add_frac_dp/n4121 ,
         \fpu_add_frac_dp/n4120 , \fpu_add_frac_dp/n4119 ,
         \fpu_add_frac_dp/n4118 , \fpu_add_frac_dp/n4117 ,
         \fpu_add_frac_dp/n4116 , \fpu_add_frac_dp/n4115 ,
         \fpu_add_frac_dp/n4114 , \fpu_add_frac_dp/n4113 ,
         \fpu_add_frac_dp/n4112 , \fpu_add_frac_dp/n4111 ,
         \fpu_add_frac_dp/n4110 , \fpu_add_frac_dp/n4109 ,
         \fpu_add_frac_dp/n4108 , \fpu_add_frac_dp/n4107 ,
         \fpu_add_frac_dp/n4106 , \fpu_add_frac_dp/n4105 ,
         \fpu_add_frac_dp/n4104 , \fpu_add_frac_dp/n4103 ,
         \fpu_add_frac_dp/n4102 , \fpu_add_frac_dp/n4101 ,
         \fpu_add_frac_dp/n4100 , \fpu_add_frac_dp/n4099 ,
         \fpu_add_frac_dp/n4098 , \fpu_add_frac_dp/n4097 ,
         \fpu_add_frac_dp/n4096 , \fpu_add_frac_dp/n4095 ,
         \fpu_add_frac_dp/n4094 , \fpu_add_frac_dp/n4093 ,
         \fpu_add_frac_dp/n4092 , \fpu_add_frac_dp/n4091 ,
         \fpu_add_frac_dp/n4090 , \fpu_add_frac_dp/n4089 ,
         \fpu_add_frac_dp/n4088 , \fpu_add_frac_dp/n4087 ,
         \fpu_add_frac_dp/n4086 , \fpu_add_frac_dp/n4085 ,
         \fpu_add_frac_dp/n4084 , \fpu_add_frac_dp/n4083 ,
         \fpu_add_frac_dp/n4082 , \fpu_add_frac_dp/n4081 ,
         \fpu_add_frac_dp/n4080 , \fpu_add_frac_dp/n4079 ,
         \fpu_add_frac_dp/n4078 , \fpu_add_frac_dp/n4077 ,
         \fpu_add_frac_dp/n4076 , \fpu_add_frac_dp/n4075 ,
         \fpu_add_frac_dp/n4074 , \fpu_add_frac_dp/n4073 ,
         \fpu_add_frac_dp/n4072 , \fpu_add_frac_dp/n4071 ,
         \fpu_add_frac_dp/n4070 , \fpu_add_frac_dp/n4069 ,
         \fpu_add_frac_dp/n4068 , \fpu_add_frac_dp/n4067 ,
         \fpu_add_frac_dp/n4066 , \fpu_add_frac_dp/n4065 ,
         \fpu_add_frac_dp/n4064 , \fpu_add_frac_dp/n4063 ,
         \fpu_add_frac_dp/n4062 , \fpu_add_frac_dp/n4061 ,
         \fpu_add_frac_dp/n4060 , \fpu_add_frac_dp/n4059 ,
         \fpu_add_frac_dp/n4058 , \fpu_add_frac_dp/n4057 ,
         \fpu_add_frac_dp/n4056 , \fpu_add_frac_dp/n4055 ,
         \fpu_add_frac_dp/n4054 , \fpu_add_frac_dp/n4053 ,
         \fpu_add_frac_dp/n4052 , \fpu_add_frac_dp/n4051 ,
         \fpu_add_frac_dp/n4050 , \fpu_add_frac_dp/n4049 ,
         \fpu_add_frac_dp/n4048 , \fpu_add_frac_dp/n4047 ,
         \fpu_add_frac_dp/n4046 , \fpu_add_frac_dp/n4045 ,
         \fpu_add_frac_dp/n4044 , \fpu_add_frac_dp/n4043 ,
         \fpu_add_frac_dp/n4042 , \fpu_add_frac_dp/n4041 ,
         \fpu_add_frac_dp/n4040 , \fpu_add_frac_dp/n4039 ,
         \fpu_add_frac_dp/n4038 , \fpu_add_frac_dp/n4037 ,
         \fpu_add_frac_dp/n4036 , \fpu_add_frac_dp/n4035 ,
         \fpu_add_frac_dp/n4034 , \fpu_add_frac_dp/n4033 ,
         \fpu_add_frac_dp/n4032 , \fpu_add_frac_dp/n4031 ,
         \fpu_add_frac_dp/n4030 , \fpu_add_frac_dp/n4029 ,
         \fpu_add_frac_dp/n4028 , \fpu_add_frac_dp/n4027 ,
         \fpu_add_frac_dp/n4026 , \fpu_add_frac_dp/n4025 ,
         \fpu_add_frac_dp/n4024 , \fpu_add_frac_dp/n4023 ,
         \fpu_add_frac_dp/n4022 , \fpu_add_frac_dp/n4021 ,
         \fpu_add_frac_dp/n4020 , \fpu_add_frac_dp/n4019 ,
         \fpu_add_frac_dp/n4018 , \fpu_add_frac_dp/n4017 ,
         \fpu_add_frac_dp/n4016 , \fpu_add_frac_dp/n4015 ,
         \fpu_add_frac_dp/n4014 , \fpu_add_frac_dp/n4013 ,
         \fpu_add_frac_dp/n4012 , \fpu_add_frac_dp/n4011 ,
         \fpu_add_frac_dp/n4010 , \fpu_add_frac_dp/n4009 ,
         \fpu_add_frac_dp/n4008 , \fpu_add_frac_dp/n4007 ,
         \fpu_add_frac_dp/n4006 , \fpu_add_frac_dp/n4005 ,
         \fpu_add_frac_dp/n4004 , \fpu_add_frac_dp/n4003 ,
         \fpu_add_frac_dp/n4002 , \fpu_add_frac_dp/n4001 ,
         \fpu_add_frac_dp/n4000 , \fpu_add_frac_dp/n3999 ,
         \fpu_add_frac_dp/n3998 , \fpu_add_frac_dp/n3997 ,
         \fpu_add_frac_dp/n3996 , \fpu_add_frac_dp/n3995 ,
         \fpu_add_frac_dp/n3994 , \fpu_add_frac_dp/n3993 ,
         \fpu_add_frac_dp/n3992 , \fpu_add_frac_dp/n3991 ,
         \fpu_add_frac_dp/n3990 , \fpu_add_frac_dp/n3989 ,
         \fpu_add_frac_dp/n3988 , \fpu_add_frac_dp/n3987 ,
         \fpu_add_frac_dp/n3986 , \fpu_add_frac_dp/n3985 ,
         \fpu_add_frac_dp/n3984 , \fpu_add_frac_dp/n3983 ,
         \fpu_add_frac_dp/n3982 , \fpu_add_frac_dp/n3981 ,
         \fpu_add_frac_dp/n3980 , \fpu_add_frac_dp/n3979 ,
         \fpu_add_frac_dp/n3978 , \fpu_add_frac_dp/n3977 ,
         \fpu_add_frac_dp/n3976 , \fpu_add_frac_dp/n3975 ,
         \fpu_add_frac_dp/n3974 , \fpu_add_frac_dp/n3973 ,
         \fpu_add_frac_dp/n3972 , \fpu_add_frac_dp/n3971 ,
         \fpu_add_frac_dp/n3970 , \fpu_add_frac_dp/n3969 ,
         \fpu_add_frac_dp/n3968 , \fpu_add_frac_dp/n3967 ,
         \fpu_add_frac_dp/n3966 , \fpu_add_frac_dp/n3965 ,
         \fpu_add_frac_dp/n3964 , \fpu_add_frac_dp/n3963 ,
         \fpu_add_frac_dp/n3962 , \fpu_add_frac_dp/n3961 ,
         \fpu_add_frac_dp/n3960 , \fpu_add_frac_dp/n3959 ,
         \fpu_add_frac_dp/n3958 , \fpu_add_frac_dp/n3957 ,
         \fpu_add_frac_dp/n3956 , \fpu_add_frac_dp/n3955 ,
         \fpu_add_frac_dp/n3954 , \fpu_add_frac_dp/n3953 ,
         \fpu_add_frac_dp/n3952 , \fpu_add_frac_dp/n3951 ,
         \fpu_add_frac_dp/n3950 , \fpu_add_frac_dp/n3949 ,
         \fpu_add_frac_dp/n3948 , \fpu_add_frac_dp/n3947 ,
         \fpu_add_frac_dp/n3946 , \fpu_add_frac_dp/n3945 ,
         \fpu_add_frac_dp/n3944 , \fpu_add_frac_dp/n3943 ,
         \fpu_add_frac_dp/n3942 , \fpu_add_frac_dp/n3941 ,
         \fpu_add_frac_dp/n3940 , \fpu_add_frac_dp/n3939 ,
         \fpu_add_frac_dp/n3938 , \fpu_add_frac_dp/n3937 ,
         \fpu_add_frac_dp/n3936 , \fpu_add_frac_dp/n3935 ,
         \fpu_add_frac_dp/n3934 , \fpu_add_frac_dp/n3933 ,
         \fpu_add_frac_dp/n3932 , \fpu_add_frac_dp/n3931 ,
         \fpu_add_frac_dp/n3930 , \fpu_add_frac_dp/n3929 ,
         \fpu_add_frac_dp/n3928 , \fpu_add_frac_dp/n3927 ,
         \fpu_add_frac_dp/n3926 , \fpu_add_frac_dp/n3925 ,
         \fpu_add_frac_dp/n3924 , \fpu_add_frac_dp/n3923 ,
         \fpu_add_frac_dp/n3922 , \fpu_add_frac_dp/n3921 ,
         \fpu_add_frac_dp/n3920 , \fpu_add_frac_dp/n3919 ,
         \fpu_add_frac_dp/n3918 , \fpu_add_frac_dp/n3917 ,
         \fpu_add_frac_dp/n3916 , \fpu_add_frac_dp/n3915 ,
         \fpu_add_frac_dp/n3914 , \fpu_add_frac_dp/n3913 ,
         \fpu_add_frac_dp/n3912 , \fpu_add_frac_dp/n3911 ,
         \fpu_add_frac_dp/n3910 , \fpu_add_frac_dp/n3909 ,
         \fpu_add_frac_dp/n3908 , \fpu_add_frac_dp/n3907 ,
         \fpu_add_frac_dp/n3906 , \fpu_add_frac_dp/n3905 ,
         \fpu_add_frac_dp/n3904 , \fpu_add_frac_dp/n3903 ,
         \fpu_add_frac_dp/n3902 , \fpu_add_frac_dp/n3901 ,
         \fpu_add_frac_dp/n3900 , \fpu_add_frac_dp/n3899 ,
         \fpu_add_frac_dp/n3898 , \fpu_add_frac_dp/n3897 ,
         \fpu_add_frac_dp/n3896 , \fpu_add_frac_dp/n3895 ,
         \fpu_add_frac_dp/n3894 , \fpu_add_frac_dp/n3893 ,
         \fpu_add_frac_dp/n3892 , \fpu_add_frac_dp/n3891 ,
         \fpu_add_frac_dp/n3890 , \fpu_add_frac_dp/n3889 ,
         \fpu_add_frac_dp/n3888 , \fpu_add_frac_dp/n3887 ,
         \fpu_add_frac_dp/n3886 , \fpu_add_frac_dp/n3885 ,
         \fpu_add_frac_dp/n3884 , \fpu_add_frac_dp/n3883 ,
         \fpu_add_frac_dp/n3882 , \fpu_add_frac_dp/n3881 ,
         \fpu_add_frac_dp/n3880 , \fpu_add_frac_dp/n3879 ,
         \fpu_add_frac_dp/n3878 , \fpu_add_frac_dp/n3877 ,
         \fpu_add_frac_dp/n3876 , \fpu_add_frac_dp/n3875 ,
         \fpu_add_frac_dp/n3874 , \fpu_add_frac_dp/n3873 ,
         \fpu_add_frac_dp/n3872 , \fpu_add_frac_dp/n3871 ,
         \fpu_add_frac_dp/n3870 , \fpu_add_frac_dp/n3869 ,
         \fpu_add_frac_dp/n3868 , \fpu_add_frac_dp/n3867 ,
         \fpu_add_frac_dp/n3866 , \fpu_add_frac_dp/n3865 ,
         \fpu_add_frac_dp/n3864 , \fpu_add_frac_dp/n3863 ,
         \fpu_add_frac_dp/n3862 , \fpu_add_frac_dp/n3861 ,
         \fpu_add_frac_dp/n3860 , \fpu_add_frac_dp/n3859 ,
         \fpu_add_frac_dp/n3858 , \fpu_add_frac_dp/n3857 ,
         \fpu_add_frac_dp/n3856 , \fpu_add_frac_dp/n3855 ,
         \fpu_add_frac_dp/n3854 , \fpu_add_frac_dp/n3853 ,
         \fpu_add_frac_dp/n3852 , \fpu_add_frac_dp/n3851 ,
         \fpu_add_frac_dp/n3850 , \fpu_add_frac_dp/n3849 ,
         \fpu_add_frac_dp/n3848 , \fpu_add_frac_dp/n3847 ,
         \fpu_add_frac_dp/n3846 , \fpu_add_frac_dp/n3845 ,
         \fpu_add_frac_dp/n3844 , \fpu_add_frac_dp/n3843 ,
         \fpu_add_frac_dp/n3842 , \fpu_add_frac_dp/n3841 ,
         \fpu_add_frac_dp/n3840 , \fpu_add_frac_dp/n3839 ,
         \fpu_add_frac_dp/n3838 , \fpu_add_frac_dp/n3837 ,
         \fpu_add_frac_dp/n3836 , \fpu_add_frac_dp/n3835 ,
         \fpu_add_frac_dp/n3834 , \fpu_add_frac_dp/n3833 ,
         \fpu_add_frac_dp/n3832 , \fpu_add_frac_dp/n3831 ,
         \fpu_add_frac_dp/n3830 , \fpu_add_frac_dp/n3829 ,
         \fpu_add_frac_dp/n3828 , \fpu_add_frac_dp/n3827 ,
         \fpu_add_frac_dp/n3826 , \fpu_add_frac_dp/n3825 ,
         \fpu_add_frac_dp/n3824 , \fpu_add_frac_dp/n3823 ,
         \fpu_add_frac_dp/n3822 , \fpu_add_frac_dp/n3821 ,
         \fpu_add_frac_dp/n3820 , \fpu_add_frac_dp/n3819 ,
         \fpu_add_frac_dp/n3818 , \fpu_add_frac_dp/n3817 ,
         \fpu_add_frac_dp/n3816 , \fpu_add_frac_dp/n3815 ,
         \fpu_add_frac_dp/n3814 , \fpu_add_frac_dp/n3813 ,
         \fpu_add_frac_dp/n3812 , \fpu_add_frac_dp/n3811 ,
         \fpu_add_frac_dp/n3810 , \fpu_add_frac_dp/n3809 ,
         \fpu_add_frac_dp/n3808 , \fpu_add_frac_dp/n3807 ,
         \fpu_add_frac_dp/n3806 , \fpu_add_frac_dp/n3805 ,
         \fpu_add_frac_dp/n3804 , \fpu_add_frac_dp/n3803 ,
         \fpu_add_frac_dp/n3802 , \fpu_add_frac_dp/n3801 ,
         \fpu_add_frac_dp/n3800 , \fpu_add_frac_dp/n3799 ,
         \fpu_add_frac_dp/n3798 , \fpu_add_frac_dp/n3797 ,
         \fpu_add_frac_dp/n3796 , \fpu_add_frac_dp/n3795 ,
         \fpu_add_frac_dp/n3794 , \fpu_add_frac_dp/n3792 ,
         \fpu_add_frac_dp/n3791 , \fpu_add_frac_dp/n3790 ,
         \fpu_add_frac_dp/n3789 , \fpu_add_frac_dp/n3788 ,
         \fpu_add_frac_dp/n3787 , \fpu_add_frac_dp/n3786 ,
         \fpu_add_frac_dp/n3785 , \fpu_add_frac_dp/n3784 ,
         \fpu_add_frac_dp/n3783 , \fpu_add_frac_dp/n3782 ,
         \fpu_add_frac_dp/n3781 , \fpu_add_frac_dp/n3780 ,
         \fpu_add_frac_dp/n3779 , \fpu_add_frac_dp/n3778 ,
         \fpu_add_frac_dp/n3777 , \fpu_add_frac_dp/n3776 ,
         \fpu_add_frac_dp/n3775 , \fpu_add_frac_dp/n3774 ,
         \fpu_add_frac_dp/n3773 , \fpu_add_frac_dp/n3772 ,
         \fpu_add_frac_dp/n3771 , \fpu_add_frac_dp/n3770 ,
         \fpu_add_frac_dp/n3769 , \fpu_add_frac_dp/n3768 ,
         \fpu_add_frac_dp/n3767 , \fpu_add_frac_dp/n3766 ,
         \fpu_add_frac_dp/n3765 , \fpu_add_frac_dp/n3764 ,
         \fpu_add_frac_dp/n3763 , \fpu_add_frac_dp/n3762 ,
         \fpu_add_frac_dp/n3761 , \fpu_add_frac_dp/n3760 ,
         \fpu_add_frac_dp/n3759 , \fpu_add_frac_dp/n3758 ,
         \fpu_add_frac_dp/n3757 , \fpu_add_frac_dp/n3756 ,
         \fpu_add_frac_dp/n3755 , \fpu_add_frac_dp/n3754 ,
         \fpu_add_frac_dp/n3753 , \fpu_add_frac_dp/n3752 ,
         \fpu_add_frac_dp/n3751 , \fpu_add_frac_dp/n3750 ,
         \fpu_add_frac_dp/n3749 , \fpu_add_frac_dp/n3748 ,
         \fpu_add_frac_dp/n3747 , \fpu_add_frac_dp/n3746 ,
         \fpu_add_frac_dp/n3745 , \fpu_add_frac_dp/n3744 ,
         \fpu_add_frac_dp/n3743 , \fpu_add_frac_dp/n3742 ,
         \fpu_add_frac_dp/n3741 , \fpu_add_frac_dp/n3740 ,
         \fpu_add_frac_dp/n3739 , \fpu_add_frac_dp/n3738 ,
         \fpu_add_frac_dp/n3737 , \fpu_add_frac_dp/n3736 ,
         \fpu_add_frac_dp/n3735 , \fpu_add_frac_dp/n3734 ,
         \fpu_add_frac_dp/n3733 , \fpu_add_frac_dp/n3732 ,
         \fpu_add_frac_dp/n3731 , \fpu_add_frac_dp/n3730 ,
         \fpu_add_frac_dp/n3729 , \fpu_add_frac_dp/n3728 ,
         \fpu_add_frac_dp/n3727 , \fpu_add_frac_dp/n3726 ,
         \fpu_add_frac_dp/n3725 , \fpu_add_frac_dp/n3724 ,
         \fpu_add_frac_dp/n3723 , \fpu_add_frac_dp/n3722 ,
         \fpu_add_frac_dp/n3721 , \fpu_add_frac_dp/n3720 ,
         \fpu_add_frac_dp/n3719 , \fpu_add_frac_dp/n3718 ,
         \fpu_add_frac_dp/n3717 , \fpu_add_frac_dp/n3716 ,
         \fpu_add_frac_dp/n3715 , \fpu_add_frac_dp/n3714 ,
         \fpu_add_frac_dp/n3713 , \fpu_add_frac_dp/n3712 ,
         \fpu_add_frac_dp/n3711 , \fpu_add_frac_dp/n3710 ,
         \fpu_add_frac_dp/n3709 , \fpu_add_frac_dp/n3708 ,
         \fpu_add_frac_dp/n3707 , \fpu_add_frac_dp/n3706 ,
         \fpu_add_frac_dp/n3705 , \fpu_add_frac_dp/n3704 ,
         \fpu_add_frac_dp/n3703 , \fpu_add_frac_dp/n3702 ,
         \fpu_add_frac_dp/n3701 , \fpu_add_frac_dp/n3700 ,
         \fpu_add_frac_dp/n3699 , \fpu_add_frac_dp/n3698 ,
         \fpu_add_frac_dp/n3697 , \fpu_add_frac_dp/n3696 ,
         \fpu_add_frac_dp/n3695 , \fpu_add_frac_dp/n3694 ,
         \fpu_add_frac_dp/n3693 , \fpu_add_frac_dp/n3692 ,
         \fpu_add_frac_dp/n3691 , \fpu_add_frac_dp/n3690 ,
         \fpu_add_frac_dp/n3689 , \fpu_add_frac_dp/n3688 ,
         \fpu_add_frac_dp/n3687 , \fpu_add_frac_dp/n3686 ,
         \fpu_add_frac_dp/n3685 , \fpu_add_frac_dp/n3684 ,
         \fpu_add_frac_dp/n3683 , \fpu_add_frac_dp/n3682 ,
         \fpu_add_frac_dp/n3681 , \fpu_add_frac_dp/n3680 ,
         \fpu_add_frac_dp/n3679 , \fpu_add_frac_dp/n3678 ,
         \fpu_add_frac_dp/n3677 , \fpu_add_frac_dp/n3676 ,
         \fpu_add_frac_dp/n3675 , \fpu_add_frac_dp/n3674 ,
         \fpu_add_frac_dp/n3673 , \fpu_add_frac_dp/n3672 ,
         \fpu_add_frac_dp/n3671 , \fpu_add_frac_dp/n3670 ,
         \fpu_add_frac_dp/n3669 , \fpu_add_frac_dp/n3668 ,
         \fpu_add_frac_dp/n3667 , \fpu_add_frac_dp/n3666 ,
         \fpu_add_frac_dp/n3665 , \fpu_add_frac_dp/n3664 ,
         \fpu_add_frac_dp/n3663 , \fpu_add_frac_dp/n3662 ,
         \fpu_add_frac_dp/n3661 , \fpu_add_frac_dp/n3660 ,
         \fpu_add_frac_dp/n3659 , \fpu_add_frac_dp/n3658 ,
         \fpu_add_frac_dp/n3657 , \fpu_add_frac_dp/n3656 ,
         \fpu_add_frac_dp/n3655 , \fpu_add_frac_dp/n3654 ,
         \fpu_add_frac_dp/n3653 , \fpu_add_frac_dp/n3652 ,
         \fpu_add_frac_dp/n3651 , \fpu_add_frac_dp/n3650 ,
         \fpu_add_frac_dp/n3649 , \fpu_add_frac_dp/n3648 ,
         \fpu_add_frac_dp/n3647 , \fpu_add_frac_dp/n3646 ,
         \fpu_add_frac_dp/n3645 , \fpu_add_frac_dp/n3644 ,
         \fpu_add_frac_dp/n3643 , \fpu_add_frac_dp/n3642 ,
         \fpu_add_frac_dp/n3641 , \fpu_add_frac_dp/n3640 ,
         \fpu_add_frac_dp/n3639 , \fpu_add_frac_dp/n3638 ,
         \fpu_add_frac_dp/n3637 , \fpu_add_frac_dp/n3636 ,
         \fpu_add_frac_dp/n3635 , \fpu_add_frac_dp/n3634 ,
         \fpu_add_frac_dp/n3633 , \fpu_add_frac_dp/n3632 ,
         \fpu_add_frac_dp/n3631 , \fpu_add_frac_dp/n3630 ,
         \fpu_add_frac_dp/n3629 , \fpu_add_frac_dp/n3628 ,
         \fpu_add_frac_dp/n3627 , \fpu_add_frac_dp/n3626 ,
         \fpu_add_frac_dp/n3625 , \fpu_add_frac_dp/n3624 ,
         \fpu_add_frac_dp/n3623 , \fpu_add_frac_dp/n3622 ,
         \fpu_add_frac_dp/n3621 , \fpu_add_frac_dp/n3620 ,
         \fpu_add_frac_dp/n3619 , \fpu_add_frac_dp/n3618 ,
         \fpu_add_frac_dp/n3617 , \fpu_add_frac_dp/n3616 ,
         \fpu_add_frac_dp/n3615 , \fpu_add_frac_dp/n3614 ,
         \fpu_add_frac_dp/n3613 , \fpu_add_frac_dp/n3612 ,
         \fpu_add_frac_dp/n3611 , \fpu_add_frac_dp/n3610 ,
         \fpu_add_frac_dp/n3609 , \fpu_add_frac_dp/n3608 ,
         \fpu_add_frac_dp/n3607 , \fpu_add_frac_dp/n3606 ,
         \fpu_add_frac_dp/n3605 , \fpu_add_frac_dp/n3604 ,
         \fpu_add_frac_dp/n3603 , \fpu_add_frac_dp/n3602 ,
         \fpu_add_frac_dp/n3601 , \fpu_add_frac_dp/n3600 ,
         \fpu_add_frac_dp/n3599 , \fpu_add_frac_dp/n3598 ,
         \fpu_add_frac_dp/n3597 , \fpu_add_frac_dp/n3596 ,
         \fpu_add_frac_dp/n3595 , \fpu_add_frac_dp/n3594 ,
         \fpu_add_frac_dp/n3593 , \fpu_add_frac_dp/n3592 ,
         \fpu_add_frac_dp/n3591 , \fpu_add_frac_dp/n3590 ,
         \fpu_add_frac_dp/n3589 , \fpu_add_frac_dp/n3588 ,
         \fpu_add_frac_dp/n3587 , \fpu_add_frac_dp/n3586 ,
         \fpu_add_frac_dp/n3585 , \fpu_add_frac_dp/n3584 ,
         \fpu_add_frac_dp/n3583 , \fpu_add_frac_dp/n3582 ,
         \fpu_add_frac_dp/n3581 , \fpu_add_frac_dp/n3580 ,
         \fpu_add_frac_dp/n3579 , \fpu_add_frac_dp/n3578 ,
         \fpu_add_frac_dp/n3577 , \fpu_add_frac_dp/n3576 ,
         \fpu_add_frac_dp/n3575 , \fpu_add_frac_dp/n3574 ,
         \fpu_add_frac_dp/n3573 , \fpu_add_frac_dp/n3572 ,
         \fpu_add_frac_dp/n3571 , \fpu_add_frac_dp/n3570 ,
         \fpu_add_frac_dp/n3569 , \fpu_add_frac_dp/n3568 ,
         \fpu_add_frac_dp/n3567 , \fpu_add_frac_dp/n3566 ,
         \fpu_add_frac_dp/n3565 , \fpu_add_frac_dp/n3564 ,
         \fpu_add_frac_dp/n3563 , \fpu_add_frac_dp/n3562 ,
         \fpu_add_frac_dp/n3561 , \fpu_add_frac_dp/n3560 ,
         \fpu_add_frac_dp/n3559 , \fpu_add_frac_dp/n3558 ,
         \fpu_add_frac_dp/n3557 , \fpu_add_frac_dp/n3556 ,
         \fpu_add_frac_dp/n3555 , \fpu_add_frac_dp/n3554 ,
         \fpu_add_frac_dp/n3553 , \fpu_add_frac_dp/n3552 ,
         \fpu_add_frac_dp/n3551 , \fpu_add_frac_dp/n3550 ,
         \fpu_add_frac_dp/n3549 , \fpu_add_frac_dp/n3548 ,
         \fpu_add_frac_dp/n3547 , \fpu_add_frac_dp/n3546 ,
         \fpu_add_frac_dp/n3545 , \fpu_add_frac_dp/n3544 ,
         \fpu_add_frac_dp/n3543 , \fpu_add_frac_dp/n3542 ,
         \fpu_add_frac_dp/n3541 , \fpu_add_frac_dp/n3540 ,
         \fpu_add_frac_dp/n3539 , \fpu_add_frac_dp/n3538 ,
         \fpu_add_frac_dp/n3537 , \fpu_add_frac_dp/n3536 ,
         \fpu_add_frac_dp/n3535 , \fpu_add_frac_dp/n3534 ,
         \fpu_add_frac_dp/n3533 , \fpu_add_frac_dp/n3532 ,
         \fpu_add_frac_dp/n3531 , \fpu_add_frac_dp/n3530 ,
         \fpu_add_frac_dp/n3529 , \fpu_add_frac_dp/n3528 ,
         \fpu_add_frac_dp/n3527 , \fpu_add_frac_dp/n3526 ,
         \fpu_add_frac_dp/n3525 , \fpu_add_frac_dp/n3524 ,
         \fpu_add_frac_dp/n3523 , \fpu_add_frac_dp/n3522 ,
         \fpu_add_frac_dp/n3521 , \fpu_add_frac_dp/n3520 ,
         \fpu_add_frac_dp/n3519 , \fpu_add_frac_dp/n3518 ,
         \fpu_add_frac_dp/n3517 , \fpu_add_frac_dp/n3516 ,
         \fpu_add_frac_dp/n3515 , \fpu_add_frac_dp/n3514 ,
         \fpu_add_frac_dp/n3513 , \fpu_add_frac_dp/n3512 ,
         \fpu_add_frac_dp/n3511 , \fpu_add_frac_dp/n3510 ,
         \fpu_add_frac_dp/n3509 , \fpu_add_frac_dp/n3508 ,
         \fpu_add_frac_dp/n3507 , \fpu_add_frac_dp/n3506 ,
         \fpu_add_frac_dp/n3505 , \fpu_add_frac_dp/n3504 ,
         \fpu_add_frac_dp/n3503 , \fpu_add_frac_dp/n3502 ,
         \fpu_add_frac_dp/n3501 , \fpu_add_frac_dp/n3500 ,
         \fpu_add_frac_dp/n3499 , \fpu_add_frac_dp/n3498 ,
         \fpu_add_frac_dp/n3497 , \fpu_add_frac_dp/n3496 ,
         \fpu_add_frac_dp/n3495 , \fpu_add_frac_dp/n3494 ,
         \fpu_add_frac_dp/n3493 , \fpu_add_frac_dp/n3492 ,
         \fpu_add_frac_dp/n3491 , \fpu_add_frac_dp/n3490 ,
         \fpu_add_frac_dp/n3489 , \fpu_add_frac_dp/n3488 ,
         \fpu_add_frac_dp/n3487 , \fpu_add_frac_dp/n3486 ,
         \fpu_add_frac_dp/n3485 , \fpu_add_frac_dp/n3484 ,
         \fpu_add_frac_dp/n3483 , \fpu_add_frac_dp/n3482 ,
         \fpu_add_frac_dp/n3481 , \fpu_add_frac_dp/n3480 ,
         \fpu_add_frac_dp/n3479 , \fpu_add_frac_dp/n3478 ,
         \fpu_add_frac_dp/n3477 , \fpu_add_frac_dp/n3476 ,
         \fpu_add_frac_dp/n3475 , \fpu_add_frac_dp/n3474 ,
         \fpu_add_frac_dp/n3473 , \fpu_add_frac_dp/n3472 ,
         \fpu_add_frac_dp/n3471 , \fpu_add_frac_dp/n3470 ,
         \fpu_add_frac_dp/n3469 , \fpu_add_frac_dp/n3468 ,
         \fpu_add_frac_dp/n3467 , \fpu_add_frac_dp/n3466 ,
         \fpu_add_frac_dp/n3465 , \fpu_add_frac_dp/n3464 ,
         \fpu_add_frac_dp/n3463 , \fpu_add_frac_dp/n3462 ,
         \fpu_add_frac_dp/n3461 , \fpu_add_frac_dp/n3460 ,
         \fpu_add_frac_dp/n3459 , \fpu_add_frac_dp/n3458 ,
         \fpu_add_frac_dp/n3457 , \fpu_add_frac_dp/n3456 ,
         \fpu_add_frac_dp/n3455 , \fpu_add_frac_dp/n3454 ,
         \fpu_add_frac_dp/n3453 , \fpu_add_frac_dp/n3452 ,
         \fpu_add_frac_dp/n3451 , \fpu_add_frac_dp/n3450 ,
         \fpu_add_frac_dp/n3449 , \fpu_add_frac_dp/n3448 ,
         \fpu_add_frac_dp/n3447 , \fpu_add_frac_dp/n3446 ,
         \fpu_add_frac_dp/n3445 , \fpu_add_frac_dp/n3444 ,
         \fpu_add_frac_dp/n3443 , \fpu_add_frac_dp/n3442 ,
         \fpu_add_frac_dp/n3441 , \fpu_add_frac_dp/n3440 ,
         \fpu_add_frac_dp/n3439 , \fpu_add_frac_dp/n3438 ,
         \fpu_add_frac_dp/n3437 , \fpu_add_frac_dp/n3436 ,
         \fpu_add_frac_dp/n3435 , \fpu_add_frac_dp/n3434 ,
         \fpu_add_frac_dp/n3433 , \fpu_add_frac_dp/n3432 ,
         \fpu_add_frac_dp/n3431 , \fpu_add_frac_dp/n3430 ,
         \fpu_add_frac_dp/n3429 , \fpu_add_frac_dp/n3428 ,
         \fpu_add_frac_dp/n3427 , \fpu_add_frac_dp/n3426 ,
         \fpu_add_frac_dp/n3425 , \fpu_add_frac_dp/n3424 ,
         \fpu_add_frac_dp/n3423 , \fpu_add_frac_dp/n3422 ,
         \fpu_add_frac_dp/n3421 , \fpu_add_frac_dp/n3420 ,
         \fpu_add_frac_dp/n3419 , \fpu_add_frac_dp/n3418 ,
         \fpu_add_frac_dp/n3417 , \fpu_add_frac_dp/n3416 ,
         \fpu_add_frac_dp/n3415 , \fpu_add_frac_dp/n3414 ,
         \fpu_add_frac_dp/n3413 , \fpu_add_frac_dp/n3412 ,
         \fpu_add_frac_dp/n3411 , \fpu_add_frac_dp/n3410 ,
         \fpu_add_frac_dp/n3409 , \fpu_add_frac_dp/n3408 ,
         \fpu_add_frac_dp/n3407 , \fpu_add_frac_dp/n3406 ,
         \fpu_add_frac_dp/n3405 , \fpu_add_frac_dp/n3404 ,
         \fpu_add_frac_dp/n3403 , \fpu_add_frac_dp/n3402 ,
         \fpu_add_frac_dp/n3401 , \fpu_add_frac_dp/n3400 ,
         \fpu_add_frac_dp/n3399 , \fpu_add_frac_dp/n3398 ,
         \fpu_add_frac_dp/n3397 , \fpu_add_frac_dp/n3396 ,
         \fpu_add_frac_dp/n3395 , \fpu_add_frac_dp/n3394 ,
         \fpu_add_frac_dp/n3393 , \fpu_add_frac_dp/n3392 ,
         \fpu_add_frac_dp/n3391 , \fpu_add_frac_dp/n3390 ,
         \fpu_add_frac_dp/n3389 , \fpu_add_frac_dp/n3388 ,
         \fpu_add_frac_dp/n3387 , \fpu_add_frac_dp/n3386 ,
         \fpu_add_frac_dp/n3385 , \fpu_add_frac_dp/n3384 ,
         \fpu_add_frac_dp/n3383 , \fpu_add_frac_dp/n3382 ,
         \fpu_add_frac_dp/n3381 , \fpu_add_frac_dp/n3380 ,
         \fpu_add_frac_dp/n3379 , \fpu_add_frac_dp/n3378 ,
         \fpu_add_frac_dp/n3377 , \fpu_add_frac_dp/n3376 ,
         \fpu_add_frac_dp/n3375 , \fpu_add_frac_dp/n1391 ,
         \fpu_add_frac_dp/n1384 , \fpu_add_frac_dp/n1382 ,
         \fpu_add_frac_dp/n1355 , \fpu_add_frac_dp/n1354 ,
         \fpu_add_frac_dp/n1352 , \fpu_add_frac_dp/n1335 ,
         \fpu_add_frac_dp/n1333 , \fpu_add_frac_dp/n1332 ,
         \fpu_add_frac_dp/n1315 , \fpu_add_frac_dp/n1314 ,
         \fpu_add_frac_dp/n1215 , \fpu_add_frac_dp/n1213 ,
         \fpu_add_frac_dp/n1123 , \fpu_add_frac_dp/n1122 ,
         \fpu_add_frac_dp/n1119 , \fpu_add_frac_dp/n1115 ,
         \fpu_add_frac_dp/n1109 , \fpu_add_frac_dp/n1107 ,
         \fpu_add_frac_dp/n1106 , \fpu_add_frac_dp/n1105 ,
         \fpu_add_frac_dp/n1104 , \fpu_add_frac_dp/n1103 ,
         \fpu_add_frac_dp/n1096 , \fpu_add_frac_dp/n1095 ,
         \fpu_add_frac_dp/n1094 , \fpu_add_frac_dp/n1093 ,
         \fpu_add_frac_dp/n1090 , \fpu_add_frac_dp/n1089 ,
         \fpu_add_frac_dp/n1088 , \fpu_add_frac_dp/n1087 ,
         \fpu_add_frac_dp/n1086 , \fpu_add_frac_dp/n1085 ,
         \fpu_add_frac_dp/n1084 , \fpu_add_frac_dp/n1083 ,
         \fpu_add_frac_dp/n1082 , \fpu_add_frac_dp/n1070 ,
         \fpu_add_frac_dp/n1067 , \fpu_add_frac_dp/n1056 ,
         \fpu_add_frac_dp/n1050 , \fpu_add_frac_dp/n1048 ,
         \fpu_add_frac_dp/n1045 , \fpu_add_frac_dp/n1044 ,
         \fpu_add_frac_dp/n1007 , \fpu_add_frac_dp/n1006 ,
         \fpu_add_frac_dp/n1005 , \fpu_add_frac_dp/n1004 ,
         \fpu_add_frac_dp/n1003 , \fpu_add_frac_dp/n1002 ,
         \fpu_add_frac_dp/n1001 , \fpu_add_frac_dp/n998 ,
         \fpu_add_frac_dp/n965 , \fpu_add_frac_dp/n945 ,
         \fpu_add_frac_dp/n943 , \fpu_add_frac_dp/n942 ,
         \fpu_add_frac_dp/n940 , \fpu_add_frac_dp/n937 ,
         \fpu_add_frac_dp/n935 , \fpu_add_frac_dp/n934 ,
         \fpu_add_frac_dp/n933 , \fpu_add_frac_dp/n932 ,
         \fpu_add_frac_dp/n931 , \fpu_add_frac_dp/n930 ,
         \fpu_add_frac_dp/n929 , \fpu_add_frac_dp/n928 ,
         \fpu_add_frac_dp/n927 , \fpu_add_frac_dp/n922 ,
         \fpu_add_frac_dp/n921 , \fpu_add_frac_dp/n920 ,
         \fpu_add_frac_dp/n919 , \fpu_add_frac_dp/n918 ,
         \fpu_add_frac_dp/n917 , \fpu_add_frac_dp/n913 ,
         \fpu_add_frac_dp/n912 , \fpu_add_frac_dp/n911 ,
         \fpu_add_frac_dp/n908 , \fpu_add_frac_dp/n907 ,
         \fpu_add_frac_dp/n905 , \fpu_add_frac_dp/n904 ,
         \fpu_add_frac_dp/n903 , \fpu_add_frac_dp/n901 ,
         \fpu_add_frac_dp/n900 , \fpu_add_frac_dp/n898 ,
         \fpu_add_frac_dp/n895 , \fpu_add_frac_dp/n851 ,
         \fpu_add_frac_dp/n848 , \fpu_add_frac_dp/n847 ,
         \fpu_add_frac_dp/n846 , \fpu_add_frac_dp/n845 ,
         \fpu_add_frac_dp/n844 , \fpu_add_frac_dp/n843 ,
         \fpu_add_frac_dp/n841 , \fpu_add_frac_dp/n839 ,
         \fpu_add_frac_dp/n834 , \fpu_add_frac_dp/n833 ,
         \fpu_add_frac_dp/n824 , \fpu_add_frac_dp/n823 ,
         \fpu_add_frac_dp/n822 , \fpu_add_frac_dp/n817 ,
         \fpu_add_frac_dp/n816 , \fpu_add_frac_dp/n815 ,
         \fpu_add_frac_dp/n814 , \fpu_add_frac_dp/n781 ,
         \fpu_add_frac_dp/n780 , \fpu_add_frac_dp/n779 ,
         \fpu_add_frac_dp/n778 , \fpu_add_frac_dp/n777 ,
         \fpu_add_frac_dp/n774 , \fpu_add_frac_dp/n773 ,
         \fpu_add_frac_dp/n772 , \fpu_add_frac_dp/n771 ,
         \fpu_add_frac_dp/n770 , \fpu_add_frac_dp/n769 ,
         \fpu_add_frac_dp/n768 , \fpu_add_frac_dp/n767 ,
         \fpu_add_frac_dp/n766 , \fpu_add_frac_dp/n763 ,
         \fpu_add_frac_dp/n762 , \fpu_add_frac_dp/n761 ,
         \fpu_add_frac_dp/n760 , \fpu_add_frac_dp/n759 ,
         \fpu_add_frac_dp/n758 , \fpu_add_frac_dp/n757 ,
         \fpu_add_frac_dp/n756 , \fpu_add_frac_dp/n755 ,
         \fpu_add_frac_dp/n752 , \fpu_add_frac_dp/n751 ,
         \fpu_add_frac_dp/n750 , \fpu_add_frac_dp/n749 ,
         \fpu_add_frac_dp/n747 , \fpu_add_frac_dp/n745 ,
         \fpu_add_frac_dp/n744 , \fpu_add_frac_dp/n743 ,
         \fpu_add_frac_dp/n741 , \fpu_add_frac_dp/n736 ,
         \fpu_add_frac_dp/n735 , \fpu_add_frac_dp/n734 ,
         \fpu_add_frac_dp/n733 , \fpu_add_frac_dp/n732 ,
         \fpu_add_frac_dp/n731 , \fpu_add_frac_dp/n730 ,
         \fpu_add_frac_dp/n729 , \fpu_add_frac_dp/n728 ,
         \fpu_add_frac_dp/n727 , \fpu_add_frac_dp/n726 ,
         \fpu_add_frac_dp/n725 , \fpu_add_frac_dp/n724 ,
         \fpu_add_frac_dp/n723 , \fpu_add_frac_dp/n722 ,
         \fpu_add_frac_dp/n721 , \fpu_add_frac_dp/n720 ,
         \fpu_add_frac_dp/n719 , \fpu_add_frac_dp/n718 ,
         \fpu_add_frac_dp/n717 , \fpu_add_frac_dp/n716 ,
         \fpu_add_frac_dp/n715 , \fpu_add_frac_dp/n714 ,
         \fpu_add_frac_dp/n713 , \fpu_add_frac_dp/n712 ,
         \fpu_add_frac_dp/n711 , \fpu_add_frac_dp/n710 ,
         \fpu_add_frac_dp/n709 , \fpu_add_frac_dp/n708 ,
         \fpu_add_frac_dp/n707 , \fpu_add_frac_dp/n706 ,
         \fpu_add_frac_dp/n705 , \fpu_add_frac_dp/n704 ,
         \fpu_add_frac_dp/n703 , \fpu_add_frac_dp/n702 ,
         \fpu_add_frac_dp/n701 , \fpu_add_frac_dp/n700 ,
         \fpu_add_frac_dp/n699 , \fpu_add_frac_dp/n698 ,
         \fpu_add_frac_dp/n697 , \fpu_add_frac_dp/n696 ,
         \fpu_add_frac_dp/n695 , \fpu_add_frac_dp/n694 ,
         \fpu_add_frac_dp/n693 , \fpu_add_frac_dp/n692 ,
         \fpu_add_frac_dp/n691 , \fpu_add_frac_dp/n690 ,
         \fpu_add_frac_dp/n689 , \fpu_add_frac_dp/n688 ,
         \fpu_add_frac_dp/n687 , \fpu_add_frac_dp/n686 ,
         \fpu_add_frac_dp/n685 , \fpu_add_frac_dp/n684 ,
         \fpu_add_frac_dp/n683 , \fpu_add_frac_dp/n682 ,
         \fpu_add_frac_dp/n681 , \fpu_add_frac_dp/n680 ,
         \fpu_add_frac_dp/n679 , \fpu_add_frac_dp/n678 ,
         \fpu_add_frac_dp/n677 , \fpu_add_frac_dp/n676 ,
         \fpu_add_frac_dp/n675 , \fpu_add_frac_dp/n674 ,
         \fpu_add_frac_dp/n673 , \fpu_add_frac_dp/n670 ,
         \fpu_add_frac_dp/n668 , \fpu_add_frac_dp/n666 ,
         \fpu_add_frac_dp/n664 , \fpu_add_frac_dp/n662 ,
         \fpu_add_frac_dp/n660 , \fpu_add_frac_dp/n659 ,
         \fpu_add_frac_dp/n658 , \fpu_add_frac_dp/n654 ,
         \fpu_add_frac_dp/n652 , \fpu_add_frac_dp/n650 ,
         \fpu_add_frac_dp/n649 , \fpu_add_frac_dp/n648 ,
         \fpu_add_frac_dp/n647 , \fpu_add_frac_dp/n646 ,
         \fpu_add_frac_dp/n645 , \fpu_add_frac_dp/n644 ,
         \fpu_add_frac_dp/n643 , \fpu_add_frac_dp/n642 ,
         \fpu_add_frac_dp/n641 , \fpu_add_frac_dp/n640 ,
         \fpu_add_frac_dp/n639 , \fpu_add_frac_dp/n638 ,
         \fpu_add_frac_dp/n637 , \fpu_add_frac_dp/n636 ,
         \fpu_add_frac_dp/n635 , \fpu_add_frac_dp/n634 ,
         \fpu_add_frac_dp/n633 , \fpu_add_frac_dp/n632 ,
         \fpu_add_frac_dp/n631 , \fpu_add_frac_dp/n630 ,
         \fpu_add_frac_dp/n629 , \fpu_add_frac_dp/n628 ,
         \fpu_add_frac_dp/n627 , \fpu_add_frac_dp/n626 ,
         \fpu_add_frac_dp/n625 , \fpu_add_frac_dp/n624 ,
         \fpu_add_frac_dp/n623 , \fpu_add_frac_dp/n622 ,
         \fpu_add_frac_dp/n621 , \fpu_add_frac_dp/n620 ,
         \fpu_add_frac_dp/n619 , \fpu_add_frac_dp/n618 ,
         \fpu_add_frac_dp/n617 , \fpu_add_frac_dp/n616 ,
         \fpu_add_frac_dp/n615 , \fpu_add_frac_dp/n614 ,
         \fpu_add_frac_dp/n613 , \fpu_add_frac_dp/n612 ,
         \fpu_add_frac_dp/n611 , \fpu_add_frac_dp/n610 ,
         \fpu_add_frac_dp/n609 , \fpu_add_frac_dp/n608 ,
         \fpu_add_frac_dp/n607 , \fpu_add_frac_dp/n606 ,
         \fpu_add_frac_dp/n605 , \fpu_add_frac_dp/n604 ,
         \fpu_add_frac_dp/n603 , \fpu_add_frac_dp/n602 ,
         \fpu_add_frac_dp/n601 , \fpu_add_frac_dp/n600 ,
         \fpu_add_frac_dp/n599 , \fpu_add_frac_dp/n598 ,
         \fpu_add_frac_dp/n596 , \fpu_add_frac_dp/n594 ,
         \fpu_add_frac_dp/n593 , \fpu_add_frac_dp/n592 ,
         \fpu_add_frac_dp/n589 , \fpu_add_frac_dp/n586 ,
         \fpu_add_frac_dp/n584 , \fpu_add_frac_dp/n583 ,
         \fpu_add_frac_dp/n582 , \fpu_add_frac_dp/n580 ,
         \fpu_add_frac_dp/n579 , \fpu_add_frac_dp/n577 ,
         \fpu_add_frac_dp/n576 , \fpu_add_frac_dp/n575 ,
         \fpu_add_frac_dp/n574 , \fpu_add_frac_dp/n573 ,
         \fpu_add_frac_dp/n572 , \fpu_add_frac_dp/n571 ,
         \fpu_add_frac_dp/n570 , \fpu_add_frac_dp/n569 ,
         \fpu_add_frac_dp/n568 , \fpu_add_frac_dp/n567 ,
         \fpu_add_frac_dp/n566 , \fpu_add_frac_dp/n565 ,
         \fpu_add_frac_dp/n564 , \fpu_add_frac_dp/n563 ,
         \fpu_add_frac_dp/n562 , \fpu_add_frac_dp/n561 ,
         \fpu_add_frac_dp/n560 , \fpu_add_frac_dp/n559 ,
         \fpu_add_frac_dp/n558 , \fpu_add_frac_dp/n557 ,
         \fpu_add_frac_dp/n556 , \fpu_add_frac_dp/n555 ,
         \fpu_add_frac_dp/n554 , \fpu_add_frac_dp/n553 ,
         \fpu_add_frac_dp/n552 , \fpu_add_frac_dp/n551 ,
         \fpu_add_frac_dp/n550 , \fpu_add_frac_dp/n549 ,
         \fpu_add_frac_dp/n548 , \fpu_add_frac_dp/n547 ,
         \fpu_add_frac_dp/n546 , \fpu_add_frac_dp/n545 ,
         \fpu_add_frac_dp/n544 , \fpu_add_frac_dp/n543 ,
         \fpu_add_frac_dp/n542 , \fpu_add_frac_dp/n541 ,
         \fpu_add_frac_dp/n540 , \fpu_add_frac_dp/n539 ,
         \fpu_add_frac_dp/n538 , \fpu_add_frac_dp/n537 ,
         \fpu_add_frac_dp/n536 , \fpu_add_frac_dp/n535 ,
         \fpu_add_frac_dp/n534 , \fpu_add_frac_dp/n533 ,
         \fpu_add_frac_dp/n532 , \fpu_add_frac_dp/n531 ,
         \fpu_add_frac_dp/n530 , \fpu_add_frac_dp/n529 ,
         \fpu_add_frac_dp/n528 , \fpu_add_frac_dp/n527 ,
         \fpu_add_frac_dp/n526 , \fpu_add_frac_dp/n525 ,
         \fpu_add_frac_dp/n524 , \fpu_add_frac_dp/n523 ,
         \fpu_add_frac_dp/n522 , \fpu_add_frac_dp/n521 ,
         \fpu_add_frac_dp/n520 , \fpu_add_frac_dp/n519 ,
         \fpu_add_frac_dp/n518 , \fpu_add_frac_dp/n517 ,
         \fpu_add_frac_dp/n516 , \fpu_add_frac_dp/n515 ,
         \fpu_add_frac_dp/n514 , \fpu_add_frac_dp/n513 ,
         \fpu_add_frac_dp/n512 , \fpu_add_frac_dp/n511 ,
         \fpu_add_frac_dp/n510 , \fpu_add_frac_dp/n509 ,
         \fpu_add_frac_dp/n508 , \fpu_add_frac_dp/n507 ,
         \fpu_add_frac_dp/n506 , \fpu_add_frac_dp/n505 ,
         \fpu_add_frac_dp/n504 , \fpu_add_frac_dp/n503 ,
         \fpu_add_frac_dp/n502 , \fpu_add_frac_dp/n501 ,
         \fpu_add_frac_dp/n500 , \fpu_add_frac_dp/n498 ,
         \fpu_add_frac_dp/n496 , \fpu_add_frac_dp/n494 ,
         \fpu_add_frac_dp/n492 , \fpu_add_frac_dp/n490 ,
         \fpu_add_frac_dp/n488 , \fpu_add_frac_dp/n486 ,
         \fpu_add_frac_dp/n484 , \fpu_add_frac_dp/n482 ,
         \fpu_add_frac_dp/n480 , \fpu_add_frac_dp/n478 ,
         \fpu_add_frac_dp/n476 , \fpu_add_frac_dp/n474 ,
         \fpu_add_frac_dp/n472 , \fpu_add_frac_dp/n470 ,
         \fpu_add_frac_dp/n468 , \fpu_add_frac_dp/n466 ,
         \fpu_add_frac_dp/n464 , \fpu_add_frac_dp/n462 ,
         \fpu_add_frac_dp/n460 , \fpu_add_frac_dp/n458 ,
         \fpu_add_frac_dp/n456 , \fpu_add_frac_dp/n454 ,
         \fpu_add_frac_dp/n452 , \fpu_add_frac_dp/n450 ,
         \fpu_add_frac_dp/n448 , \fpu_add_frac_dp/n446 ,
         \fpu_add_frac_dp/n444 , \fpu_add_frac_dp/n442 ,
         \fpu_add_frac_dp/n440 , \fpu_add_frac_dp/n438 ,
         \fpu_add_frac_dp/n436 , \fpu_add_frac_dp/n434 ,
         \fpu_add_frac_dp/n432 , \fpu_add_frac_dp/n430 ,
         \fpu_add_frac_dp/n428 , \fpu_add_frac_dp/n426 ,
         \fpu_add_frac_dp/n424 , \fpu_add_frac_dp/n422 ,
         \fpu_add_frac_dp/n420 , \fpu_add_frac_dp/n418 ,
         \fpu_add_frac_dp/n416 , \fpu_add_frac_dp/n414 ,
         \fpu_add_frac_dp/n412 , \fpu_add_frac_dp/n410 ,
         \fpu_add_frac_dp/n408 , \fpu_add_frac_dp/n406 ,
         \fpu_add_frac_dp/n404 , \fpu_add_frac_dp/n402 ,
         \fpu_add_frac_dp/n400 , \fpu_add_frac_dp/n398 ,
         \fpu_add_frac_dp/n396 , \fpu_add_frac_dp/n394 ,
         \fpu_add_frac_dp/n392 , \fpu_add_frac_dp/n390 ,
         \fpu_add_frac_dp/n388 , \fpu_add_frac_dp/n386 ,
         \fpu_add_frac_dp/n384 , \fpu_add_frac_dp/n382 ,
         \fpu_add_frac_dp/n380 , \fpu_add_frac_dp/n378 ,
         \fpu_add_frac_dp/n377 , \fpu_add_frac_dp/n376 ,
         \fpu_add_frac_dp/n375 , \fpu_add_frac_dp/n374 ,
         \fpu_add_frac_dp/n373 , \fpu_add_frac_dp/n372 ,
         \fpu_add_frac_dp/n371 , \fpu_add_frac_dp/n370 ,
         \fpu_add_frac_dp/n369 , \fpu_add_frac_dp/n368 ,
         \fpu_add_frac_dp/n367 , \fpu_add_frac_dp/n366 ,
         \fpu_add_frac_dp/n365 , \fpu_add_frac_dp/n364 ,
         \fpu_add_frac_dp/n363 , \fpu_add_frac_dp/n362 ,
         \fpu_add_frac_dp/n361 , \fpu_add_frac_dp/n360 ,
         \fpu_add_frac_dp/n359 , \fpu_add_frac_dp/n358 ,
         \fpu_add_frac_dp/n357 , \fpu_add_frac_dp/n356 ,
         \fpu_add_frac_dp/n355 , \fpu_add_frac_dp/n354 ,
         \fpu_add_frac_dp/n353 , \fpu_add_frac_dp/n352 ,
         \fpu_add_frac_dp/n351 , \fpu_add_frac_dp/n350 ,
         \fpu_add_frac_dp/n349 , \fpu_add_frac_dp/n348 ,
         \fpu_add_frac_dp/n347 , \fpu_add_frac_dp/n346 ,
         \fpu_add_frac_dp/n345 , \fpu_add_frac_dp/n344 ,
         \fpu_add_frac_dp/n343 , \fpu_add_frac_dp/n342 ,
         \fpu_add_frac_dp/n341 , \fpu_add_frac_dp/n340 ,
         \fpu_add_frac_dp/n339 , \fpu_add_frac_dp/n338 ,
         \fpu_add_frac_dp/n337 , \fpu_add_frac_dp/n336 ,
         \fpu_add_frac_dp/n335 , \fpu_add_frac_dp/n334 ,
         \fpu_add_frac_dp/n333 , \fpu_add_frac_dp/n332 ,
         \fpu_add_frac_dp/n331 , \fpu_add_frac_dp/n330 ,
         \fpu_add_frac_dp/n329 , \fpu_add_frac_dp/n328 ,
         \fpu_add_frac_dp/n327 , \fpu_add_frac_dp/n326 ,
         \fpu_add_frac_dp/n325 , \fpu_add_frac_dp/n324 ,
         \fpu_add_frac_dp/n323 , \fpu_add_frac_dp/n322 ,
         \fpu_add_frac_dp/n321 , \fpu_add_frac_dp/n320 ,
         \fpu_add_frac_dp/n319 , \fpu_add_frac_dp/n318 ,
         \fpu_add_frac_dp/n317 , \fpu_add_frac_dp/n316 ,
         \fpu_add_frac_dp/n315 , \fpu_add_frac_dp/n313 ,
         \fpu_add_frac_dp/n311 , \fpu_add_frac_dp/n309 ,
         \fpu_add_frac_dp/n307 , \fpu_add_frac_dp/n305 ,
         \fpu_add_frac_dp/n303 , \fpu_add_frac_dp/n301 ,
         \fpu_add_frac_dp/n299 , \fpu_add_frac_dp/n297 ,
         \fpu_add_frac_dp/n295 , \fpu_add_frac_dp/n293 ,
         \fpu_add_frac_dp/n291 , \fpu_add_frac_dp/n289 ,
         \fpu_add_frac_dp/n287 , \fpu_add_frac_dp/n285 ,
         \fpu_add_frac_dp/n283 , \fpu_add_frac_dp/n282 ,
         \fpu_add_frac_dp/n281 , \fpu_add_frac_dp/n280 ,
         \fpu_add_frac_dp/n279 , \fpu_add_frac_dp/n278 ,
         \fpu_add_frac_dp/n277 , \fpu_add_frac_dp/n276 ,
         \fpu_add_frac_dp/n275 , \fpu_add_frac_dp/n274 ,
         \fpu_add_frac_dp/n273 , \fpu_add_frac_dp/n272 ,
         \fpu_add_frac_dp/n271 , \fpu_add_frac_dp/n270 ,
         \fpu_add_frac_dp/n269 , \fpu_add_frac_dp/n268 ,
         \fpu_add_frac_dp/n267 , \fpu_add_frac_dp/n266 ,
         \fpu_add_frac_dp/n265 , \fpu_add_frac_dp/n264 ,
         \fpu_add_frac_dp/n263 , \fpu_add_frac_dp/n262 ,
         \fpu_add_frac_dp/n261 , \fpu_add_frac_dp/n260 ,
         \fpu_add_frac_dp/n259 , \fpu_add_frac_dp/n258 ,
         \fpu_add_frac_dp/n257 , \fpu_add_frac_dp/n256 ,
         \fpu_add_frac_dp/n255 , \fpu_add_frac_dp/n254 ,
         \fpu_add_frac_dp/n253 , \fpu_add_frac_dp/n252 ,
         \fpu_add_frac_dp/n251 , \fpu_add_frac_dp/n250 ,
         \fpu_add_frac_dp/n249 , \fpu_add_frac_dp/n248 ,
         \fpu_add_frac_dp/n247 , \fpu_add_frac_dp/n246 ,
         \fpu_add_frac_dp/n245 , \fpu_add_frac_dp/n244 ,
         \fpu_add_frac_dp/n243 , \fpu_add_frac_dp/n242 ,
         \fpu_add_frac_dp/n241 , \fpu_add_frac_dp/n240 ,
         \fpu_add_frac_dp/n239 , \fpu_add_frac_dp/n238 ,
         \fpu_add_frac_dp/n237 , \fpu_add_frac_dp/n236 ,
         \fpu_add_frac_dp/n235 , \fpu_add_frac_dp/n234 ,
         \fpu_add_frac_dp/n233 , \fpu_add_frac_dp/n232 ,
         \fpu_add_frac_dp/n231 , \fpu_add_frac_dp/n230 ,
         \fpu_add_frac_dp/n229 , \fpu_add_frac_dp/n228 ,
         \fpu_add_frac_dp/n227 , \fpu_add_frac_dp/n226 ,
         \fpu_add_frac_dp/n225 , \fpu_add_frac_dp/n224 ,
         \fpu_add_frac_dp/n223 , \fpu_add_frac_dp/n222 ,
         \fpu_add_frac_dp/n221 , \fpu_add_frac_dp/n220 ,
         \fpu_add_frac_dp/n219 , \fpu_add_frac_dp/n218 ,
         \fpu_add_frac_dp/n217 , \fpu_add_frac_dp/n216 ,
         \fpu_add_frac_dp/n215 , \fpu_add_frac_dp/n214 ,
         \fpu_add_frac_dp/n213 , \fpu_add_frac_dp/n212 ,
         \fpu_add_frac_dp/n211 , \fpu_add_frac_dp/n210 ,
         \fpu_add_frac_dp/n209 , \fpu_add_frac_dp/n208 ,
         \fpu_add_frac_dp/n207 , \fpu_add_frac_dp/n206 ,
         \fpu_add_frac_dp/n205 , \fpu_add_frac_dp/n204 ,
         \fpu_add_frac_dp/n203 , \fpu_add_frac_dp/n202 ,
         \fpu_add_frac_dp/n201 , \fpu_add_frac_dp/n200 ,
         \fpu_add_frac_dp/n199 , \fpu_add_frac_dp/n198 ,
         \fpu_add_frac_dp/n197 , \fpu_add_frac_dp/n196 ,
         \fpu_add_frac_dp/n195 , \fpu_add_frac_dp/n194 ,
         \fpu_add_frac_dp/n193 , \fpu_add_frac_dp/n192 ,
         \fpu_add_frac_dp/n191 , \fpu_add_frac_dp/n190 ,
         \fpu_add_frac_dp/n189 , \fpu_add_frac_dp/n188 ,
         \fpu_add_frac_dp/n187 , \fpu_add_frac_dp/n134 ,
         \fpu_add_frac_dp/n132 , \fpu_add_frac_dp/n129 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N3 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N8 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N9 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N13 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N14 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N15 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N16 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N17 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N18 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N19 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N20 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N21 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N22 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N23 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N24 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N25 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N26 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N27 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N28 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N29 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N30 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N31 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N32 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N33 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N34 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N35 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N36 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N37 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N38 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N39 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N40 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N41 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N42 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N43 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N44 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N45 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N46 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N47 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N48 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N49 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N50 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N51 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N52 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N53 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N54 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N55 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N56 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N57 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N58 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N59 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N60 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N61 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N62 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N63 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N64 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N65 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N66 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N4 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N5 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N6 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N7 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N8 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N9 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N10 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N11 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N12 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N13 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N14 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N15 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N16 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N17 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N18 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N19 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N20 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N21 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N22 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N23 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N24 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N25 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N26 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N27 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N28 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N29 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N30 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N31 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N32 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N33 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N34 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N35 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N36 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N37 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N38 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N39 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N40 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N41 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N42 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N43 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N44 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N45 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N46 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N47 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N48 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N49 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N50 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N51 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N52 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N53 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N54 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N55 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N56 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N57 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N58 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N59 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N60 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N61 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N62 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N63 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N64 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N65 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N66 ,
         \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N3 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N4 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N5 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N6 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N7 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N8 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N9 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N10 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N11 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N12 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N13 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N14 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N15 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N16 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N17 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N18 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N19 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N20 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N21 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N22 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N23 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N24 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N25 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N26 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N27 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N28 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N29 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N30 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N31 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N32 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N33 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N34 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N35 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N36 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N37 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N38 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N39 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N40 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N41 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N42 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N43 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N44 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N45 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N46 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N47 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N48 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N49 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N50 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N51 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N52 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N53 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N54 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N55 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N56 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N57 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N58 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N59 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N60 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N61 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N62 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N63 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N64 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N65 ,
         \fpu_add_frac_dp/i_a3stg_frac2/N66 ,
         \fpu_add_frac_dp/ckbuf_add_frac_dp/N1 ,
         \fpu_add_frac_dp/ckbuf_add_frac_dp/clken ,
         \fpu_add_frac_dp/a5stg_in_of ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[63] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[62] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[61] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[60] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[59] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[58] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[57] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[56] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[55] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[54] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[53] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[52] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[51] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[50] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[49] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[48] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[47] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[46] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[45] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[44] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[43] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[42] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[41] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[40] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[39] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[38] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[37] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[36] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[35] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[34] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[33] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[32] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[31] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[30] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[29] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[28] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[27] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[26] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[25] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[24] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[23] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[22] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[21] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[20] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[19] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[18] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[17] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[16] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[15] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[14] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[13] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[12] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[11] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[10] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[9] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[8] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[7] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[6] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[5] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[4] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[3] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[2] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre2[1] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[63] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[62] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[61] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[60] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[59] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[58] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[57] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[56] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[55] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[54] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[53] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[52] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[51] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[50] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[49] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[48] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[47] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[46] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[45] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[44] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[43] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[42] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[41] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[40] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[39] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[38] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[37] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[36] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[35] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[34] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[33] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[32] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[31] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[30] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[29] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[28] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[27] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[26] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[25] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[24] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[23] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[22] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[21] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[20] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[19] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[18] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[17] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[16] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[15] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[14] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[13] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[12] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[11] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[10] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[9] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[8] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[7] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[6] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[5] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[4] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[3] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[2] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre3[1] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[63] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[62] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[61] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[60] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[59] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[58] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[57] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[56] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[55] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[54] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[53] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[52] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[51] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[50] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[49] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[48] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[47] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[46] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[45] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[44] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[43] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[42] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[41] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[40] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[39] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[38] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[37] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[36] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[35] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[34] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[33] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[32] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[31] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[30] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[29] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[28] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[27] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[26] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[25] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[24] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[23] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[22] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[21] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[20] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[19] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[18] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[17] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[16] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[15] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[14] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[13] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[12] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[11] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[10] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[9] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[8] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[7] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[6] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[5] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[4] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[3] ,
         \fpu_add_frac_dp/a4stg_rnd_frac_pre1[2] ,
         \fpu_add_frac_dp/a4stg_shl_cnt_dec54_1[1] ,
         \fpu_add_frac_dp/a3stg_fracadd[0] , \fpu_add_frac_dp/a3stg_frac2[63] ,
         \fpu_add_frac_dp/a2stg_shr_cnt[5] ,
         \fpu_add_frac_dp/a2stg_shr_cnt_4[3] ,
         \fpu_add_frac_dp/a2stg_frac2a[58] , \fpu_add_frac_dp/a1stg_in2[3] ,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888;
  assign so = 1'b0;
  assign add_exc_out[1] = 1'b0;

  DFFX1 \fpu_add_ctl/i_a2stg_fracadd_frac2/q_reg[0]  ( .D(\fpu_add_ctl/n540 ), 
        .CLK(rclk), .Q(n155), .QN(\fpu_add_ctl/n1 ) );
  DFFX1 \fpu_add_ctl/i_add_nx_out/q_reg[0]  ( .D(\fpu_add_ctl/n541 ), .CLK(
        rclk), .Q(\fpu_add_ctl/add_nx_out ), .QN(\fpu_add_ctl/n2 ) );
  DFFX1 \fpu_add_ctl/i_add_uf_out/q_reg[0]  ( .D(\fpu_add_ctl/n542 ), .CLK(
        rclk), .Q(add_exc_out[2]), .QN(\fpu_add_ctl/n3 ) );
  DFFX1 \fpu_add_ctl/i_add_of_out_tmp2/q_reg[0]  ( .D(\fpu_add_ctl/n543 ), 
        .CLK(rclk), .Q(\fpu_add_ctl/add_of_out_tmp2 ), .QN(\fpu_add_ctl/n4 )
         );
  DFFX1 \fpu_add_ctl/i_add_of_out_tmp1/q_reg[0]  ( .D(\fpu_add_ctl/n544 ), 
        .CLK(rclk), .Q(n1234), .QN(\fpu_add_ctl/n5 ) );
  DFFX1 \fpu_add_ctl/i_add_nv_out/q_reg[0]  ( .D(\fpu_add_ctl/n545 ), .CLK(
        rclk), .Q(add_exc_out[4]) );
  DFFX1 \fpu_add_ctl/i_a4stg_nx/q_reg[0]  ( .D(\fpu_add_ctl/n546 ), .CLK(rclk), 
        .Q(n1245), .QN(\fpu_add_ctl/n7 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_nx2/q_reg[0]  ( .D(\fpu_add_ctl/n547 ), .CLK(rclk), .Q(n513) );
  DFFX1 \fpu_add_ctl/i_a4stg_of_mask/q_reg[0]  ( .D(\fpu_add_ctl/n548 ), .CLK(
        rclk), .Q(n452), .QN(\fpu_add_ctl/n9 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_of_mask2/q_reg[0]  ( .D(\fpu_add_ctl/n549 ), 
        .CLK(rclk), .Q(n905) );
  DFFX1 \fpu_add_ctl/i_a4stg_nv/q_reg[0]  ( .D(\fpu_add_ctl/n550 ), .CLK(rclk), 
        .Q(n1074) );
  DFFX1 \fpu_add_ctl/i_a4stg_nv2/q_reg[0]  ( .D(\fpu_add_ctl/n551 ), .CLK(rclk), .Q(n512) );
  DFFX1 \fpu_add_ctl/i_a3stg_nx_tmp3/q_reg[0]  ( .D(\fpu_add_ctl/n552 ), .CLK(
        rclk), .Q(n1265), .QN(\fpu_add_ctl/n13 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_nx_tmp2/q_reg[0]  ( .D(\fpu_add_ctl/n553 ), .CLK(
        rclk), .Q(n1272), .QN(\fpu_add_ctl/n14 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_nx_tmp1/q_reg[0]  ( .D(\fpu_add_ctl/n554 ), .CLK(
        rclk), .Q(n1249), .QN(\fpu_add_ctl/n15 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_a2_expadd_11/q_reg[0]  ( .D(\fpu_add_ctl/n555 ), 
        .CLK(rclk), .Q(\fpu_add_ctl/a3stg_a2_expadd_11 ), .QN(
        \fpu_add_ctl/n16 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_of_mask/q_reg[0]  ( .D(\fpu_add_ctl/n556 ), .CLK(
        rclk), .Q(n137) );
  DFFX1 \fpu_add_ctl/i_a3stg_nv/q_reg[0]  ( .D(\fpu_add_ctl/n557 ), .CLK(rclk), 
        .Q(n140) );
  DFFX1 \fpu_add_ctl/i_a2stg_of_mask/q_reg[0]  ( .D(\fpu_add_ctl/n558 ), .CLK(
        rclk), .Q(n1077) );
  DFFX1 \fpu_add_ctl/i_a2stg_nv/q_reg[0]  ( .D(\fpu_add_ctl/n559 ), .CLK(rclk), 
        .Q(n903) );
  DFFX1 \fpu_add_ctl/i_add_cc_out/q_reg[1]  ( .D(\fpu_add_ctl/n560 ), .CLK(
        rclk), .Q(add_cc_out[1]) );
  DFFX1 \fpu_add_ctl/i_add_cc_out/q_reg[0]  ( .D(\fpu_add_ctl/n561 ), .CLK(
        rclk), .Q(add_cc_out[0]) );
  DFFX1 \fpu_add_ctl/i_add_sign_out/q_reg[0]  ( .D(\fpu_add_ctl/n562 ), .CLK(
        rclk), .Q(add_sign_out) );
  DFFX1 \fpu_add_ctl/i_a4stg_cc/q_reg[1]  ( .D(\fpu_add_ctl/n563 ), .CLK(rclk), 
        .Q(n557) );
  DFFX1 \fpu_add_ctl/i_a4stg_cc/q_reg[0]  ( .D(\fpu_add_ctl/n564 ), .CLK(rclk), 
        .Q(n556) );
  DFFX1 \fpu_add_ctl/i_a4stg_sign/q_reg[0]  ( .D(\fpu_add_ctl/n565 ), .CLK(
        rclk), .Q(n444), .QN(\fpu_add_ctl/n337 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_sign2/q_reg[0]  ( .D(\fpu_add_ctl/n566 ), .CLK(
        rclk), .Q(n884) );
  DFFX1 \fpu_add_ctl/i_a3stg_cc/q_reg[1]  ( .D(\fpu_add_ctl/n567 ), .CLK(rclk), 
        .Q(n1083) );
  DFFX1 \fpu_add_ctl/i_a3stg_cc/q_reg[0]  ( .D(\fpu_add_ctl/n568 ), .CLK(rclk), 
        .Q(n1082) );
  DFFX1 \fpu_add_ctl/i_a3stg_sign/q_reg[0]  ( .D(\fpu_add_ctl/n569 ), .CLK(
        rclk), .Q(n149) );
  DFFX1 \fpu_add_ctl/i_a2stg_2inf_in/q_reg[0]  ( .D(\fpu_add_ctl/n570 ), .CLK(
        rclk), .Q(n957), .QN(\fpu_add_ctl/n31 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_2zero_in/q_reg[0]  ( .D(\fpu_add_ctl/n571 ), 
        .CLK(rclk), .Q(n1217), .QN(\fpu_add_ctl/n32 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_qnan_in1/q_reg[0]  ( .D(\fpu_add_ctl/n572 ), 
        .CLK(rclk), .Q(n1068) );
  DFFX1 \fpu_add_ctl/i_a2stg_snan_in1/q_reg[0]  ( .D(\fpu_add_ctl/n573 ), 
        .CLK(rclk), .Q(n422), .QN(\fpu_add_ctl/n311 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_qnan_in2/q_reg[0]  ( .D(\fpu_add_ctl/n574 ), 
        .CLK(rclk), .Q(n1213), .QN(\fpu_add_ctl/n34 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_snan_in2/q_reg[0]  ( .D(\fpu_add_ctl/n575 ), 
        .CLK(rclk), .Q(n1173), .QN(\fpu_add_ctl/n310 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_nan_in2/q_reg[0]  ( .D(\fpu_add_ctl/n576 ), .CLK(
        rclk), .Q(\fpu_add_ctl/a2stg_nan_in2 ), .QN(\fpu_add_ctl/n338 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_nan_in/q_reg[0]  ( .D(\fpu_add_ctl/n577 ), .CLK(
        rclk), .Q(n851), .QN(\fpu_add_ctl/n37 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_in2_gt_in1_exp/q_reg[0]  ( .D(\fpu_add_ctl/n578 ), 
        .CLK(rclk), .Q(\fpu_add_ctl/a2stg_in2_gt_in1_exp ), .QN(
        \fpu_add_ctl/n38 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_in2_eq_in1_exp/q_reg[0]  ( .D(\fpu_add_ctl/n579 ), 
        .CLK(rclk), .Q(n1004), .QN(\fpu_add_ctl/n335 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_in2_gt_in1_frac/q_reg[0]  ( .D(\fpu_add_ctl/n580 ), .CLK(rclk), .Q(n1212), .QN(\fpu_add_ctl/n39 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_in2_neq_in1_frac/q_reg[0]  ( .D(
        \fpu_add_ctl/n581 ), .CLK(rclk), .Q(n1210), .QN(\fpu_add_ctl/n40 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_sub/q_reg[0]  ( .D(\fpu_add_ctl/n582 ), .CLK(rclk), .Q(\fpu_add_ctl/n313 ), .QN(n754) );
  DFFX1 \fpu_add_ctl/i_a2stg_sign2/q_reg[0]  ( .D(\fpu_add_ctl/n583 ), .CLK(
        rclk), .Q(n270), .QN(\fpu_add_ctl/n316 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_sign1/q_reg[0]  ( .D(\fpu_add_ctl/n584 ), .CLK(
        rclk), .Q(n433), .QN(\fpu_add_ctl/n41 ) );
  DFFX1 \fpu_add_ctl/i_add_pipe_active/q_reg[0]  ( .D(
        \fpu_add_ctl/i_add_pipe_active/N7 ), .CLK(rclk), .Q(add_pipe_active)
         );
  DFFX1 \fpu_add_ctl/i_add_fcc_out/q_reg[1]  ( .D(\fpu_add_ctl/n585 ), .CLK(
        rclk), .Q(add_fcc_out[1]) );
  DFFX1 \fpu_add_ctl/i_add_fcc_out/q_reg[0]  ( .D(\fpu_add_ctl/n586 ), .CLK(
        rclk), .Q(add_fcc_out[0]) );
  DFFSSRX1 \fpu_add_ctl/i_add_id_out/q_reg[9]  ( .D(\fpu_add_ctl/n470 ), 
        .RSTB(add_id_out_in[9]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_add_ctl/add_id_out[9] ) );
  DFFSSRX1 \fpu_add_ctl/i_add_id_out/q_reg[8]  ( .D(\fpu_add_ctl/n470 ), 
        .RSTB(add_id_out_in[8]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_add_ctl/add_id_out[8] ) );
  DFFSSRX1 \fpu_add_ctl/i_add_id_out/q_reg[7]  ( .D(\fpu_add_ctl/n470 ), 
        .RSTB(add_id_out_in[7]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_add_ctl/add_id_out[7] ) );
  DFFSSRX1 \fpu_add_ctl/i_add_id_out/q_reg[6]  ( .D(\fpu_add_ctl/n470 ), 
        .RSTB(add_id_out_in[6]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_add_ctl/add_id_out[6] ) );
  DFFSSRX1 \fpu_add_ctl/i_add_id_out/q_reg[5]  ( .D(\fpu_add_ctl/n470 ), 
        .RSTB(add_id_out_in[5]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_add_ctl/add_id_out[5] ) );
  DFFSSRX1 \fpu_add_ctl/i_add_id_out/q_reg[4]  ( .D(\fpu_add_ctl/n470 ), 
        .RSTB(add_id_out_in[4]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_add_ctl/add_id_out[4] ) );
  DFFSSRX1 \fpu_add_ctl/i_add_id_out/q_reg[3]  ( .D(\fpu_add_ctl/n470 ), 
        .RSTB(add_id_out_in[3]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_add_ctl/add_id_out[3] ) );
  DFFSSRX1 \fpu_add_ctl/i_add_id_out/q_reg[2]  ( .D(\fpu_add_ctl/n470 ), 
        .RSTB(add_id_out_in[2]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_add_ctl/add_id_out[2] ) );
  DFFSSRX1 \fpu_add_ctl/i_add_id_out/q_reg[1]  ( .D(\fpu_add_ctl/n470 ), 
        .RSTB(add_id_out_in[1]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_add_ctl/add_id_out[1] ) );
  DFFSSRX1 \fpu_add_ctl/i_add_id_out/q_reg[0]  ( .D(\fpu_add_ctl/n470 ), 
        .RSTB(add_id_out_in[0]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_add_ctl/add_id_out[0] ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[17]  ( .D(\fpu_add_ctl/n606 ), .CLK(
        rclk), .Q(n1242), .QN(\fpu_add_ctl/n65 ) );
  DFFX1 \fpu_add_ctl/i_a5stg_opdec/q_reg[8]  ( .D(\fpu_add_ctl/n612 ), .CLK(
        rclk), .Q(n1157), .QN(\fpu_add_ctl/n66 ) );
  DFFX1 \fpu_add_ctl/i_a6stg_opdec/q_reg[4]  ( .D(\fpu_add_ctl/n607 ), .CLK(
        rclk), .Q(a6stg_dbl_dst) );
  DFFX1 \fpu_add_ctl/i_a5stg_opdec/q_reg[7]  ( .D(\fpu_add_ctl/n613 ), .CLK(
        rclk), .Q(n1073) );
  DFFX1 \fpu_add_ctl/i_a6stg_opdec/q_reg[3]  ( .D(\fpu_add_ctl/n608 ), .CLK(
        rclk), .Q(a6stg_sng_dst) );
  DFFX1 \fpu_add_ctl/i_a5stg_opdec/q_reg[6]  ( .D(\fpu_add_ctl/n614 ), .CLK(
        rclk), .Q(n1072) );
  DFFX1 \fpu_add_ctl/i_a6stg_opdec/q_reg[2]  ( .D(\fpu_add_ctl/n609 ), .CLK(
        rclk), .Q(a6stg_long_dst) );
  DFFX1 \fpu_add_ctl/i_a5stg_opdec/q_reg[5]  ( .D(\fpu_add_ctl/n615 ), .CLK(
        rclk), .Q(n1071) );
  DFFX1 \fpu_add_ctl/i_a6stg_opdec/q_reg[1]  ( .D(\fpu_add_ctl/n610 ), .CLK(
        rclk), .Q(a6stg_int_dst) );
  DFFX1 \fpu_add_ctl/i_a5stg_opdec/q_reg[4]  ( .D(\fpu_add_ctl/n616 ), .CLK(
        rclk), .Q(n1070) );
  DFFX1 \fpu_add_ctl/i_a6stg_opdec/q_reg[0]  ( .D(\fpu_add_ctl/n611 ), .CLK(
        rclk), .Q(a6stg_fcmpop) );
  DFFX1 \fpu_add_ctl/i_a5stg_opdec/q_reg[3]  ( .D(\fpu_add_ctl/n617 ), .CLK(
        rclk), .Q(n1069) );
  DFFX1 \fpu_add_ctl/i_a5stg_opdec/q_reg[2]  ( .D(\fpu_add_ctl/n618 ), .CLK(
        rclk), .Q(n622), .QN(\fpu_add_ctl/n315 ) );
  DFFX1 \fpu_add_ctl/i_a5stg_opdec/q_reg[1]  ( .D(\fpu_add_ctl/n619 ), .CLK(
        rclk), .Q(n552), .QN(\fpu_add_ctl/n77 ) );
  DFFX1 \fpu_add_ctl/i_a5stg_opdec/q_reg[0]  ( .D(\fpu_add_ctl/n620 ), .CLK(
        rclk), .Q(n108), .QN(\fpu_add_ctl/n78 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[16]  ( .D(\fpu_add_ctl/n621 ), .CLK(
        rclk), .Q(n339), .QN(\fpu_add_ctl/n79 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[15]  ( .D(\fpu_add_ctl/n622 ), .CLK(
        rclk), .Q(n136) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[14]  ( .D(\fpu_add_ctl/n623 ), .CLK(
        rclk), .Q(n135) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[13]  ( .D(\fpu_add_ctl/n624 ), .CLK(
        rclk), .Q(n333) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[12]  ( .D(\fpu_add_ctl/n625 ), .CLK(
        rclk), .Q(n134) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[11]  ( .D(\fpu_add_ctl/n626 ), .CLK(
        rclk), .Q(n927), .QN(\fpu_add_ctl/n939 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[10]  ( .D(\fpu_add_ctl/n627 ), .CLK(
        rclk), .Q(n490), .QN(\fpu_add_ctl/n334 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[9]  ( .D(\fpu_add_ctl/n628 ), .CLK(
        rclk), .Q(n1246), .QN(\fpu_add_ctl/n85 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[8]  ( .D(\fpu_add_ctl/n629 ), .CLK(
        rclk), .Q(n324), .QN(\fpu_add_ctl/n86 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[7]  ( .D(\fpu_add_ctl/n630 ), .CLK(
        rclk), .Q(\fpu_add_ctl/n319 ), .QN(n642) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[6]  ( .D(\fpu_add_ctl/n631 ), .CLK(
        rclk), .Q(n420), .QN(\fpu_add_ctl/n941 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[5]  ( .D(\fpu_add_ctl/n632 ), .CLK(
        rclk), .Q(n148), .QN(\fpu_add_ctl/n323 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[4]  ( .D(\fpu_add_ctl/n633 ), .CLK(
        rclk), .Q(n21), .QN(\fpu_add_ctl/n322 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[3]  ( .D(\fpu_add_ctl/n634 ), .CLK(
        rclk), .Q(n55), .QN(\fpu_add_ctl/n89 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[2]  ( .D(\fpu_add_ctl/n635 ), .CLK(
        rclk), .Q(n492), .QN(\fpu_add_ctl/n90 ) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[1]  ( .D(\fpu_add_ctl/n636 ), .CLK(
        rclk), .Q(n1032) );
  DFFX1 \fpu_add_ctl/i_a4stg_opdec/q_reg[0]  ( .D(\fpu_add_ctl/n637 ), .CLK(
        rclk), .Q(n1031) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[18]  ( .D(\fpu_add_ctl/n638 ), .CLK(
        rclk), .Q(n576) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[17]  ( .D(\fpu_add_ctl/n639 ), .CLK(
        rclk), .Q(\fpu_add_ctl/n325 ), .QN(\fpu_add_ctl/n255 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[16]  ( .D(\fpu_add_ctl/n640 ), .CLK(
        rclk), .Q(n575) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[15]  ( .D(\fpu_add_ctl/n641 ), .CLK(
        rclk), .Q(n574) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[14]  ( .D(\fpu_add_ctl/n642 ), .CLK(
        rclk), .Q(n1030) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[13]  ( .D(\fpu_add_ctl/n643 ), .CLK(
        rclk), .Q(n549), .QN(\fpu_add_ctl/n97 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[11]  ( .D(\fpu_add_ctl/n645 ), .CLK(
        rclk), .Q(n1029) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[10]  ( .D(\fpu_add_ctl/n646 ), .CLK(
        rclk), .Q(n336) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[9]  ( .D(\fpu_add_ctl/n647 ), .CLK(
        rclk), .Q(n1028) );
  DFFX1 \fpu_add_ctl/i_a4stg_rnd_mode/q_reg[0]  ( .D(\fpu_add_ctl/n649 ), 
        .CLK(rclk), .Q(\fpu_add_ctl/n307 ), .QN(n1084) );
  DFFX1 \fpu_add_ctl/i_a4stg_rnd_mode/q_reg[1]  ( .D(\fpu_add_ctl/n648 ), 
        .CLK(rclk), .Q(n291), .QN(\fpu_add_ctl/n937 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[8]  ( .D(\fpu_add_ctl/n650 ), .CLK(
        rclk), .Q(n455), .QN(\fpu_add_ctl/n101 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[7]  ( .D(\fpu_add_ctl/n651 ), .CLK(
        rclk), .Q(n895), .QN(\fpu_add_ctl/n102 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[6]  ( .D(\fpu_add_ctl/n652 ), .CLK(
        rclk), .Q(n1027) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[5]  ( .D(\fpu_add_ctl/n653 ), .CLK(
        rclk), .Q(n1026) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[4]  ( .D(\fpu_add_ctl/n654 ), .CLK(
        rclk), .Q(n1025) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[3]  ( .D(\fpu_add_ctl/n655 ), .CLK(
        rclk), .Q(\fpu_add_ctl/a3stg_opdec_9_0[3] ), .QN(a3stg_fdtos_inv) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[2]  ( .D(\fpu_add_ctl/n656 ), .CLK(
        rclk), .Q(n1024) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[1]  ( .D(\fpu_add_ctl/n657 ), .CLK(
        rclk), .Q(n573) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[0]  ( .D(\fpu_add_ctl/n658 ), .CLK(
        rclk), .Q(n572) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[20]  ( .D(\fpu_add_ctl/n671 ), .CLK(
        rclk), .Q(n547), .QN(\fpu_add_ctl/n109 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[21]  ( .D(\fpu_add_ctl/n670 ), .CLK(
        rclk), .Q(n1008), .QN(\fpu_add_ctl/n110 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[8]  ( .D(\fpu_add_ctl/n682 ), .CLK(
        rclk), .Q(n858) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[22]  ( .D(\fpu_add_ctl/n669 ), .CLK(
        rclk), .Q(n356) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[28]  ( .D(\fpu_add_ctl/n661 ), .CLK(
        rclk), .Q(n1201), .QN(\fpu_add_ctl/n113 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[30]  ( .D(\fpu_add_ctl/n659 ), .CLK(
        rclk), .Q(n1023) );
  DFFX1 \fpu_add_ctl/i_a1stg_dblop/q_reg[0]  ( .D(\fpu_add_ctl/n689 ), .CLK(
        rclk), .Q(n295) );
  DFFX1 \fpu_add_ctl/i_a1stg_sngop/q_reg[0]  ( .D(\fpu_add_ctl/n601 ), .CLK(
        rclk), .Q(n662), .QN(\fpu_add_ctl/n116 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in2_exp_neq_ffs/q_reg[0]  ( .D(\fpu_add_ctl/n600 ), .CLK(rclk), .Q(\fpu_add_ctl/n317 ), .QN(n338) );
  DFFX1 \fpu_add_ctl/i_a1stg_in2_exp_eq_0/q_reg[0]  ( .D(\fpu_add_ctl/n599 ), 
        .CLK(rclk), .Q(n1086), .QN(\fpu_add_ctl/n117 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in2_53_32_neq_0/q_reg[0]  ( .D(\fpu_add_ctl/n598 ), .CLK(rclk), .Q(n730), .QN(\fpu_add_ctl/n118 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in2_50_0_neq_0/q_reg[0]  ( .D(\fpu_add_ctl/n597 ), 
        .CLK(rclk), .Q(n731), .QN(\fpu_add_ctl/n119 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in2_63/q_reg[0]  ( .D(\fpu_add_ctl/n596 ), .CLK(
        rclk), .Q(n649), .QN(\fpu_add_ctl/n940 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in2_54/q_reg[0]  ( .D(\fpu_add_ctl/n595 ), .CLK(
        rclk), .Q(n847), .QN(\fpu_add_ctl/n333 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in2_51/q_reg[0]  ( .D(\fpu_add_ctl/n594 ), .CLK(
        rclk), .Q(n460), .QN(\fpu_add_ctl/n121 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in1_exp_neq_ffs/q_reg[0]  ( .D(\fpu_add_ctl/n593 ), .CLK(rclk), .Q(n598), .QN(\fpu_add_ctl/n324 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in1_exp_eq_0/q_reg[0]  ( .D(\fpu_add_ctl/n592 ), 
        .CLK(rclk), .Q(n1085), .QN(\fpu_add_ctl/n122 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in1_53_32_neq_0/q_reg[0]  ( .D(\fpu_add_ctl/n591 ), .CLK(rclk), .Q(n743), .QN(\fpu_add_ctl/n123 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in1_50_0_neq_0/q_reg[0]  ( .D(\fpu_add_ctl/n590 ), 
        .CLK(rclk), .Q(n744), .QN(\fpu_add_ctl/n124 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in1_63/q_reg[0]  ( .D(\fpu_add_ctl/n589 ), .CLK(
        rclk), .Q(n897), .QN(\fpu_add_ctl/n125 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in1_54/q_reg[0]  ( .D(\fpu_add_ctl/n588 ), .CLK(
        rclk), .Q(n1120), .QN(\fpu_add_ctl/n332 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_in1_51/q_reg[0]  ( .D(\fpu_add_ctl/n587 ), .CLK(
        rclk), .Q(n1119), .QN(\fpu_add_ctl/n127 ) );
  DFFSSRX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[3]  ( .D(a1stg_fdtos), .RSTB(
        \fpu_add_ctl/n47 ), .SETB(\fpu_add_ctl/n426 ), .CLK(rclk), .Q(n91), 
        .QN(\fpu_add_ctl/n336 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[6]  ( .D(\fpu_add_ctl/n684 ), .CLK(
        rclk), .Q(n571) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[13]  ( .D(\fpu_add_ctl/n677 ), .CLK(
        rclk), .Q(n128), .QN(\fpu_add_ctl/n129 ) );
  DFFSSRX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[19]  ( .D(a1stg_fsdtoix), .RSTB(
        \fpu_add_ctl/n47 ), .SETB(\fpu_add_ctl/n416 ), .CLK(rclk), .Q(
        \fpu_add_ctl/n329 ), .QN(\fpu_add_ctl/n252 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[26]  ( .D(\fpu_add_ctl/n663 ), .CLK(
        rclk), .Q(n506), .QN(\fpu_add_ctl/n130 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[29]  ( .D(\fpu_add_ctl/n660 ), .CLK(
        rclk), .Q(n651) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[14]  ( .D(\fpu_add_ctl/n676 ), .CLK(
        rclk), .Q(n1076) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[15]  ( .D(\fpu_add_ctl/n675 ), .CLK(
        rclk), .Q(n553), .QN(\fpu_add_ctl/n133 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[16]  ( .D(\fpu_add_ctl/n674 ), .CLK(
        rclk), .Q(n569) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[17]  ( .D(\fpu_add_ctl/n673 ), .CLK(
        rclk), .Q(n1022) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[4]  ( .D(\fpu_add_ctl/n685 ), .CLK(
        rclk), .Q(n570) );
  DFFSSRX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[5]  ( .D(\fpu_add_ctl/n47 ), 
        .RSTB(a1stg_faddsubs), .SETB(\fpu_add_ctl/n425 ), .CLK(rclk), .Q(n562)
         );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[27]  ( .D(\fpu_add_ctl/n662 ), .CLK(
        rclk), .Q(n1200), .QN(\fpu_add_ctl/n138 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[23]  ( .D(\fpu_add_ctl/n668 ), .CLK(
        rclk), .Q(n1187), .QN(\fpu_add_ctl/n139 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_faddsubopa/q_reg[0]  ( .D(\fpu_add_ctl/n666 ), 
        .CLK(rclk), .Q(n1233), .QN(\fpu_add_ctl/n140 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_faddsubopa/q_reg[1]  ( .D(\fpu_add_ctl/n665 ), 
        .CLK(rclk), .Q(n1218), .QN(\fpu_add_ctl/n141 ) );
  DFFX1 \fpu_add_ctl/i_a3stg_opdec/q_reg[12]  ( .D(\fpu_add_ctl/n644 ), .CLK(
        rclk), .Q(n133), .QN(\fpu_add_ctl/n142 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[24]  ( .D(\fpu_add_ctl/n667 ), .CLK(
        rclk), .Q(n640), .QN(\fpu_add_ctl/n938 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[9]  ( .D(\fpu_add_ctl/n681 ), .CLK(
        rclk), .Q(n511), .QN(\fpu_add_ctl/n143 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[25]  ( .D(\fpu_add_ctl/n664 ), .CLK(
        rclk), .Q(n1214), .QN(\fpu_add_ctl/n144 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[1]  ( .D(\fpu_add_ctl/n687 ), .CLK(
        rclk), .Q(n1001) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[10]  ( .D(\fpu_add_ctl/n680 ), .CLK(
        rclk), .Q(n757) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[12]  ( .D(\fpu_add_ctl/n678 ), .CLK(
        rclk), .Q(n421), .QN(\fpu_add_ctl/n147 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[18]  ( .D(\fpu_add_ctl/n672 ), .CLK(
        rclk), .Q(n258) );
  DFFX1 \fpu_add_ctl/i_a1stg_op/q_reg[7]  ( .D(\fpu_add_ctl/n752 ), .CLK(rclk), 
        .Q(\fpu_add_ctl/n314 ), .QN(n172) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[2]  ( .D(\fpu_add_ctl/n686 ), .CLK(
        rclk), .Q(n560) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[11]  ( .D(\fpu_add_ctl/n679 ), .CLK(
        rclk), .Q(n718), .QN(\fpu_add_ctl/n150 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_op/q_reg[6]  ( .D(\fpu_add_ctl/n751 ), .CLK(rclk), 
        .Q(\fpu_add_ctl/n312 ), .QN(n254) );
  DFFX1 \fpu_add_ctl/i_a1stg_op/q_reg[5]  ( .D(\fpu_add_ctl/n750 ), .CLK(rclk), 
        .Q(n84) );
  DFFX1 \fpu_add_ctl/i_a1stg_op/q_reg[4]  ( .D(\fpu_add_ctl/n749 ), .CLK(rclk), 
        .Q(n585), .QN(\fpu_add_ctl/n303 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_op/q_reg[3]  ( .D(\fpu_add_ctl/n748 ), .CLK(rclk), 
        .Q(n595), .QN(\fpu_add_ctl/n321 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_op/q_reg[2]  ( .D(\fpu_add_ctl/n747 ), .CLK(rclk), 
        .Q(n18), .QN(\fpu_add_ctl/n318 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_op/q_reg[1]  ( .D(\fpu_add_ctl/n746 ), .CLK(rclk), 
        .Q(n829), .QN(\fpu_add_ctl/n936 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_op/q_reg[0]  ( .D(\fpu_add_ctl/n745 ), .CLK(rclk), 
        .Q(\fpu_add_ctl/n320 ), .QN(n158) );
  DFFX1 \fpu_add_ctl/i_a4stg_fcc/q_reg[1]  ( .D(\fpu_add_ctl/n737 ), .CLK(rclk), .Q(n555) );
  DFFX1 \fpu_add_ctl/i_a3stg_fcc/q_reg[1]  ( .D(\fpu_add_ctl/n739 ), .CLK(rclk), .Q(n1013) );
  DFFX1 \fpu_add_ctl/i_a2stg_fcc/q_reg[1]  ( .D(\fpu_add_ctl/n741 ), .CLK(rclk), .Q(n564) );
  DFFX1 \fpu_add_ctl/i_a1stg_fcc/q_reg[1]  ( .D(\fpu_add_ctl/n744 ), .CLK(rclk), .Q(n1011) );
  DFFX1 \fpu_add_ctl/i_a4stg_fcc/q_reg[0]  ( .D(\fpu_add_ctl/n738 ), .CLK(rclk), .Q(n554) );
  DFFX1 \fpu_add_ctl/i_a3stg_fcc/q_reg[0]  ( .D(\fpu_add_ctl/n740 ), .CLK(rclk), .Q(n1012) );
  DFFX1 \fpu_add_ctl/i_a2stg_fcc/q_reg[0]  ( .D(\fpu_add_ctl/n742 ), .CLK(rclk), .Q(n563) );
  DFFX1 \fpu_add_ctl/i_a1stg_fcc/q_reg[0]  ( .D(\fpu_add_ctl/n743 ), .CLK(rclk), .Q(n1010) );
  DFFX1 \fpu_add_ctl/i_a5stg_id/q_reg[6]  ( .D(\fpu_add_ctl/n705 ), .CLK(rclk), 
        .Q(n888) );
  DFFX1 \fpu_add_ctl/i_a4stg_id/q_reg[6]  ( .D(\fpu_add_ctl/n715 ), .CLK(rclk), 
        .Q(n350) );
  DFFX1 \fpu_add_ctl/i_a5stg_id/q_reg[7]  ( .D(\fpu_add_ctl/n704 ), .CLK(rclk), 
        .Q(n887) );
  DFFX1 \fpu_add_ctl/i_a4stg_id/q_reg[7]  ( .D(\fpu_add_ctl/n714 ), .CLK(rclk), 
        .Q(n349) );
  DFFX1 \fpu_add_ctl/i_a5stg_id/q_reg[8]  ( .D(\fpu_add_ctl/n703 ), .CLK(rclk), 
        .Q(n886) );
  DFFX1 \fpu_add_ctl/i_a4stg_id/q_reg[8]  ( .D(\fpu_add_ctl/n713 ), .CLK(rclk), 
        .Q(n348) );
  DFFX1 \fpu_add_ctl/i_a5stg_id/q_reg[9]  ( .D(\fpu_add_ctl/n702 ), .CLK(rclk), 
        .Q(n885) );
  DFFX1 \fpu_add_ctl/i_a4stg_id/q_reg[9]  ( .D(\fpu_add_ctl/n712 ), .CLK(rclk), 
        .Q(n347) );
  DFFX1 \fpu_add_ctl/i_a5stg_id/q_reg[2]  ( .D(\fpu_add_ctl/n709 ), .CLK(rclk), 
        .Q(n892) );
  DFFX1 \fpu_add_ctl/i_a4stg_id/q_reg[2]  ( .D(\fpu_add_ctl/n719 ), .CLK(rclk), 
        .Q(n354) );
  DFFX1 \fpu_add_ctl/i_a5stg_id/q_reg[3]  ( .D(\fpu_add_ctl/n708 ), .CLK(rclk), 
        .Q(n891) );
  DFFX1 \fpu_add_ctl/i_a4stg_id/q_reg[3]  ( .D(\fpu_add_ctl/n718 ), .CLK(rclk), 
        .Q(n353) );
  DFFX1 \fpu_add_ctl/i_a5stg_id/q_reg[4]  ( .D(\fpu_add_ctl/n707 ), .CLK(rclk), 
        .Q(n890) );
  DFFX1 \fpu_add_ctl/i_a4stg_id/q_reg[4]  ( .D(\fpu_add_ctl/n717 ), .CLK(rclk), 
        .Q(n352) );
  DFFX1 \fpu_add_ctl/i_a5stg_id/q_reg[5]  ( .D(\fpu_add_ctl/n706 ), .CLK(rclk), 
        .Q(n889) );
  DFFX1 \fpu_add_ctl/i_a4stg_id/q_reg[5]  ( .D(\fpu_add_ctl/n716 ), .CLK(rclk), 
        .Q(n351) );
  DFFX1 \fpu_add_ctl/i_a3stg_id/q_reg[4]  ( .D(\fpu_add_ctl/n722 ), .CLK(rclk), 
        .Q(n89), .QN(\fpu_add_ctl/n177 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_id/q_reg[4]  ( .D(\fpu_add_ctl/n727 ), .CLK(rclk), 
        .Q(n1017) );
  DFFX1 \fpu_add_ctl/i_a1stg_id/q_reg[4]  ( .D(\fpu_add_ctl/n736 ), .CLK(rclk), 
        .Q(n566) );
  DFFX1 \fpu_add_ctl/i_a3stg_id/q_reg[3]  ( .D(\fpu_add_ctl/n723 ), .CLK(rclk), 
        .Q(n269), .QN(\fpu_add_ctl/n308 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_id/q_reg[3]  ( .D(\fpu_add_ctl/n728 ), .CLK(rclk), 
        .Q(n1016) );
  DFFX1 \fpu_add_ctl/i_a1stg_id/q_reg[3]  ( .D(\fpu_add_ctl/n735 ), .CLK(rclk), 
        .Q(n565) );
  DFFX1 \fpu_add_ctl/i_a3stg_id/q_reg[2]  ( .D(\fpu_add_ctl/n724 ), .CLK(rclk), 
        .Q(\fpu_add_ctl/a3stg_id[2] ), .QN(\fpu_add_ctl/n326 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_id/q_reg[2]  ( .D(\fpu_add_ctl/n729 ), .CLK(rclk), 
        .Q(\fpu_add_ctl/a2stg_id[2] ), .QN(\fpu_add_ctl/n182 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_id/q_reg[2]  ( .D(\fpu_add_ctl/n734 ), .CLK(rclk), 
        .Q(n1216), .QN(\fpu_add_ctl/n183 ) );
  DFFX1 \fpu_add_ctl/i_a5stg_id/q_reg[1]  ( .D(\fpu_add_ctl/n710 ), .CLK(rclk), 
        .Q(n893) );
  DFFX1 \fpu_add_ctl/i_a4stg_id/q_reg[1]  ( .D(\fpu_add_ctl/n720 ), .CLK(rclk), 
        .Q(n341) );
  DFFX1 \fpu_add_ctl/i_a3stg_id/q_reg[1]  ( .D(\fpu_add_ctl/n725 ), .CLK(rclk), 
        .Q(n1019) );
  DFFX1 \fpu_add_ctl/i_a2stg_id/q_reg[1]  ( .D(\fpu_add_ctl/n730 ), .CLK(rclk), 
        .Q(n568) );
  DFFX1 \fpu_add_ctl/i_a1stg_id/q_reg[1]  ( .D(\fpu_add_ctl/n733 ), .CLK(rclk), 
        .Q(n1015) );
  DFFX1 \fpu_add_ctl/i_a5stg_id/q_reg[0]  ( .D(\fpu_add_ctl/n711 ), .CLK(rclk), 
        .Q(n894) );
  DFFX1 \fpu_add_ctl/i_a4stg_id/q_reg[0]  ( .D(\fpu_add_ctl/n721 ), .CLK(rclk), 
        .Q(n342) );
  DFFX1 \fpu_add_ctl/i_a3stg_id/q_reg[0]  ( .D(\fpu_add_ctl/n726 ), .CLK(rclk), 
        .Q(n1018) );
  DFFX1 \fpu_add_ctl/i_a2stg_id/q_reg[0]  ( .D(\fpu_add_ctl/n731 ), .CLK(rclk), 
        .Q(n567) );
  DFFX1 \fpu_add_ctl/i_a1stg_id/q_reg[0]  ( .D(\fpu_add_ctl/n732 ), .CLK(rclk), 
        .Q(n1014) );
  DFFX1 \fpu_add_ctl/i_a4stg_rnd_mode2/q_reg[1]  ( .D(\fpu_add_ctl/n694 ), 
        .CLK(rclk), .Q(n883) );
  DFFX1 \fpu_add_ctl/i_a3stg_rnd_mode/q_reg[1]  ( .D(\fpu_add_ctl/n696 ), 
        .CLK(rclk), .Q(n147) );
  DFFX1 \fpu_add_ctl/i_a2stg_rnd_mode/q_reg[1]  ( .D(\fpu_add_ctl/n698 ), 
        .CLK(rclk), .Q(n504), .QN(\fpu_add_ctl/n196 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_rnd_mode/q_reg[1]  ( .D(\fpu_add_ctl/n701 ), 
        .CLK(rclk), .Q(n1021) );
  DFFX1 \fpu_add_ctl/i_a4stg_rnd_mode2/q_reg[0]  ( .D(\fpu_add_ctl/n695 ), 
        .CLK(rclk), .Q(n882) );
  DFFX1 \fpu_add_ctl/i_a3stg_rnd_mode/q_reg[0]  ( .D(\fpu_add_ctl/n697 ), 
        .CLK(rclk), .Q(n146) );
  DFFX1 \fpu_add_ctl/i_a2stg_rnd_mode/q_reg[0]  ( .D(\fpu_add_ctl/n699 ), 
        .CLK(rclk), .Q(n505), .QN(\fpu_add_ctl/n200 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_rnd_mode/q_reg[0]  ( .D(\fpu_add_ctl/n700 ), 
        .CLK(rclk), .Q(n1020) );
  DFFX1 \fpu_add_ctl/i_a1stg_dblopa/q_reg[3]  ( .D(\fpu_add_ctl/n693 ), .CLK(
        rclk), .Q(n915), .QN(\fpu_add_ctl/n202 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_dblopa/q_reg[2]  ( .D(\fpu_add_ctl/n692 ), .CLK(
        rclk), .Q(n325), .QN(\fpu_add_ctl/n309 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_dblopa/q_reg[1]  ( .D(\fpu_add_ctl/n691 ), .CLK(
        rclk), .Q(n44), .QN(\fpu_add_ctl/n203 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_dblopa/q_reg[0]  ( .D(\fpu_add_ctl/n690 ), .CLK(
        rclk), .Q(n700), .QN(\fpu_add_ctl/n327 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_sngopa/q_reg[3]  ( .D(\fpu_add_ctl/n605 ), .CLK(
        rclk), .Q(n129) );
  DFFX1 \fpu_add_ctl/i_a1stg_sngopa/q_reg[2]  ( .D(\fpu_add_ctl/n604 ), .CLK(
        rclk), .Q(n692), .QN(\fpu_add_ctl/n330 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_sngopa/q_reg[1]  ( .D(\fpu_add_ctl/n603 ), .CLK(
        rclk), .Q(n102), .QN(\fpu_add_ctl/n205 ) );
  DFFX1 \fpu_add_ctl/i_a1stg_sngopa/q_reg[0]  ( .D(\fpu_add_ctl/n602 ), .CLK(
        rclk), .Q(n701), .QN(\fpu_add_ctl/n328 ) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[7]  ( .D(\fpu_add_ctl/n683 ), .CLK(
        rclk), .Q(n355) );
  DFFX1 \fpu_add_ctl/i_a2stg_opdec/q_reg[0]  ( .D(\fpu_add_ctl/n688 ), .CLK(
        rclk), .Q(n849), .QN(\fpu_add_ctl/n207 ) );
  DFFSSRX1 \fpu_add_ctl/i_a6stg_opdec/q_reg[5]  ( .D(\fpu_add_ctl/n49 ), 
        .RSTB(\fpu_add_ctl/n441 ), .SETB(n586), .CLK(rclk), .QN(
        \fpu_add_ctl/n269 ) );
  DFFARX1 \fpu_add_ctl/dffrl_add_ctl/q_reg[0]  ( .D(
        \fpu_add_ctl/dffrl_add_ctl/N4 ), .CLK(rclk), .RSTB(arst_l), .Q(
        \fpu_add_ctl/add_ctl_rst_l ), .QN(\fpu_add_ctl/n210 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[10]  ( .D(\fpu_add_exp_dp/n507 ), 
        .CLK(n1566), .Q(n1238), .QN(\fpu_add_exp_dp/n1 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[9]  ( .D(\fpu_add_exp_dp/n508 ), 
        .CLK(n1566), .Q(n1232), .QN(\fpu_add_exp_dp/n2 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[8]  ( .D(\fpu_add_exp_dp/n509 ), 
        .CLK(n1566), .Q(n1231), .QN(\fpu_add_exp_dp/n3 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[7]  ( .D(\fpu_add_exp_dp/n510 ), 
        .CLK(n1566), .Q(n1230), .QN(\fpu_add_exp_dp/n4 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[6]  ( .D(\fpu_add_exp_dp/n511 ), 
        .CLK(n1566), .Q(n1229), .QN(\fpu_add_exp_dp/n5 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[5]  ( .D(\fpu_add_exp_dp/n512 ), 
        .CLK(n1566), .Q(n1228), .QN(\fpu_add_exp_dp/n6 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[4]  ( .D(\fpu_add_exp_dp/n513 ), 
        .CLK(n1566), .Q(n1227), .QN(\fpu_add_exp_dp/n7 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[3]  ( .D(\fpu_add_exp_dp/n514 ), 
        .CLK(n1566), .Q(n1226), .QN(\fpu_add_exp_dp/n8 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[2]  ( .D(\fpu_add_exp_dp/n515 ), 
        .CLK(n1566), .Q(n1225), .QN(\fpu_add_exp_dp/n9 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[1]  ( .D(\fpu_add_exp_dp/n516 ), 
        .CLK(n1566), .Q(n1237), .QN(\fpu_add_exp_dp/n10 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out4/q_reg[0]  ( .D(\fpu_add_exp_dp/n517 ), 
        .CLK(n1565), .Q(n1236), .QN(\fpu_add_exp_dp/n11 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[10]  ( .D(\fpu_add_exp_dp/n518 ), 
        .CLK(\fpu_add_exp_dp/n448 ), .Q(\fpu_add_exp_dp/add_exp_out3[10] ), 
        .QN(\fpu_add_exp_dp/n12 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[9]  ( .D(\fpu_add_exp_dp/n519 ), 
        .CLK(\fpu_add_exp_dp/n448 ), .Q(\fpu_add_exp_dp/add_exp_out3[9] ), 
        .QN(\fpu_add_exp_dp/n13 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[8]  ( .D(\fpu_add_exp_dp/n520 ), 
        .CLK(\fpu_add_exp_dp/n448 ), .Q(\fpu_add_exp_dp/add_exp_out3[8] ), 
        .QN(\fpu_add_exp_dp/n14 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[7]  ( .D(\fpu_add_exp_dp/n521 ), 
        .CLK(n1585), .Q(\fpu_add_exp_dp/add_exp_out3[7] ), .QN(
        \fpu_add_exp_dp/n15 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[6]  ( .D(\fpu_add_exp_dp/n522 ), 
        .CLK(\fpu_add_exp_dp/n448 ), .Q(\fpu_add_exp_dp/add_exp_out3[6] ), 
        .QN(\fpu_add_exp_dp/n16 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[5]  ( .D(\fpu_add_exp_dp/n523 ), 
        .CLK(n1585), .Q(\fpu_add_exp_dp/add_exp_out3[5] ), .QN(
        \fpu_add_exp_dp/n17 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[4]  ( .D(\fpu_add_exp_dp/n524 ), 
        .CLK(\fpu_add_exp_dp/n448 ), .Q(\fpu_add_exp_dp/add_exp_out3[4] ), 
        .QN(\fpu_add_exp_dp/n18 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[3]  ( .D(\fpu_add_exp_dp/n525 ), 
        .CLK(n1567), .Q(\fpu_add_exp_dp/add_exp_out3[3] ), .QN(
        \fpu_add_exp_dp/n19 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[2]  ( .D(\fpu_add_exp_dp/n526 ), 
        .CLK(n1585), .Q(\fpu_add_exp_dp/add_exp_out3[2] ), .QN(
        \fpu_add_exp_dp/n20 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[1]  ( .D(\fpu_add_exp_dp/n527 ), 
        .CLK(n1567), .Q(\fpu_add_exp_dp/add_exp_out3[1] ), .QN(
        \fpu_add_exp_dp/n21 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out3/q_reg[0]  ( .D(\fpu_add_exp_dp/n528 ), 
        .CLK(n1567), .Q(\fpu_add_exp_dp/add_exp_out3[0] ), .QN(
        \fpu_add_exp_dp/n22 ) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[10]  ( .D(\fpu_add_exp_dp/n529 ), 
        .CLK(n1565), .Q(n443) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[9]  ( .D(\fpu_add_exp_dp/n530 ), 
        .CLK(n1565), .Q(n441) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[8]  ( .D(\fpu_add_exp_dp/n531 ), 
        .CLK(n1565), .Q(n442) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[7]  ( .D(\fpu_add_exp_dp/n532 ), 
        .CLK(n1565), .Q(n732) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[6]  ( .D(\fpu_add_exp_dp/n533 ), 
        .CLK(n1565), .Q(n733) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[5]  ( .D(\fpu_add_exp_dp/n534 ), 
        .CLK(n1565), .Q(n734) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[4]  ( .D(\fpu_add_exp_dp/n535 ), 
        .CLK(n1565), .Q(n735) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[3]  ( .D(\fpu_add_exp_dp/n536 ), 
        .CLK(n1565), .Q(n736) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[2]  ( .D(\fpu_add_exp_dp/n537 ), 
        .CLK(n1565), .Q(n737) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[1]  ( .D(\fpu_add_exp_dp/n538 ), 
        .CLK(n1565), .Q(n738) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out2/q_reg[0]  ( .D(\fpu_add_exp_dp/n539 ), 
        .CLK(n1565), .Q(n764) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[10]  ( .D(\fpu_add_exp_dp/n540 ), 
        .CLK(n1567), .Q(n760) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[9]  ( .D(\fpu_add_exp_dp/n541 ), 
        .CLK(n1567), .Q(n758) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[8]  ( .D(\fpu_add_exp_dp/n542 ), 
        .CLK(n1567), .Q(n759) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[7]  ( .D(\fpu_add_exp_dp/n543 ), 
        .CLK(n1567), .Q(n434) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[6]  ( .D(\fpu_add_exp_dp/n544 ), 
        .CLK(n1567), .Q(n435) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[5]  ( .D(\fpu_add_exp_dp/n545 ), 
        .CLK(n1567), .Q(n436) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[4]  ( .D(\fpu_add_exp_dp/n546 ), 
        .CLK(n1567), .Q(n437) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[3]  ( .D(\fpu_add_exp_dp/n547 ), 
        .CLK(n1567), .Q(n438) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[2]  ( .D(\fpu_add_exp_dp/n548 ), 
        .CLK(n1567), .Q(n439) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[1]  ( .D(\fpu_add_exp_dp/n549 ), 
        .CLK(n1566), .Q(n440) );
  DFFX1 \fpu_add_exp_dp/i_add_exp_out1/q_reg[0]  ( .D(\fpu_add_exp_dp/n550 ), 
        .CLK(n1566), .Q(n454) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[11]  ( .D(\fpu_add_exp_dp/n552 ), 
        .CLK(n1572), .Q(\fpu_add_exp_dp/a4stg_exp2[11] ), .QN(
        \fpu_add_exp_dp/n46 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[10]  ( .D(\fpu_add_exp_dp/n553 ), 
        .CLK(n1573), .Q(n663), .QN(\fpu_add_exp_dp/n451 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[9]  ( .D(\fpu_add_exp_dp/n554 ), 
        .CLK(n1572), .Q(\fpu_add_exp_dp/a4stg_exp2[9] ), .QN(
        \fpu_add_exp_dp/n48 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[8]  ( .D(\fpu_add_exp_dp/n555 ), 
        .CLK(n1572), .Q(\fpu_add_exp_dp/a4stg_exp2[8] ), .QN(
        \fpu_add_exp_dp/n450 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[7]  ( .D(\fpu_add_exp_dp/n556 ), 
        .CLK(n1572), .Q(\fpu_add_exp_dp/a4stg_exp2[7] ), .QN(
        \fpu_add_exp_dp/n50 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[6]  ( .D(\fpu_add_exp_dp/n557 ), 
        .CLK(n1573), .Q(n666), .QN(\fpu_add_exp_dp/n452 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[5]  ( .D(\fpu_add_exp_dp/n558 ), 
        .CLK(n1572), .Q(n761), .QN(\fpu_add_exp_dp/n441 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[4]  ( .D(\fpu_add_exp_dp/n559 ), 
        .CLK(n1571), .Q(\fpu_add_exp_dp/a4stg_exp2[4] ), .QN(
        \fpu_add_exp_dp/n440 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[3]  ( .D(\fpu_add_exp_dp/n560 ), 
        .CLK(n1571), .Q(\fpu_add_exp_dp/a4stg_exp2[3] ), .QN(
        \fpu_add_exp_dp/n439 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[2]  ( .D(\fpu_add_exp_dp/n561 ), 
        .CLK(n1571), .Q(\fpu_add_exp_dp/a4stg_exp2[2] ), .QN(
        \fpu_add_exp_dp/n438 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[1]  ( .D(\fpu_add_exp_dp/n562 ), 
        .CLK(n1572), .Q(n643), .QN(\fpu_add_exp_dp/n437 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp2/q_reg[0]  ( .D(\fpu_add_exp_dp/n563 ), 
        .CLK(n1571), .Q(\fpu_add_exp_dp/a4stg_exp2[0] ), .QN(
        \fpu_add_exp_dp/n57 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[11]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N14 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre2[11] ), .QN(\fpu_add_exp_dp/n60 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[11]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N14 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[11] ), .QN(\fpu_add_exp_dp/n61 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[10]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N13 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre2[10] ), .QN(\fpu_add_exp_dp/n62 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[10]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N13 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[10] ), .QN(\fpu_add_exp_dp/n63 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[9]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N12 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre2[9] ), .QN(\fpu_add_exp_dp/n64 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[9]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N12 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[9] ), .QN(\fpu_add_exp_dp/n65 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[8]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N11 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre2[8] ), .QN(\fpu_add_exp_dp/n66 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[8]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N11 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[8] ), .QN(\fpu_add_exp_dp/n67 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[7]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N10 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre2[7] ), .QN(\fpu_add_exp_dp/n68 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[7]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N10 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[7] ), .QN(\fpu_add_exp_dp/n69 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[6]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N9 ), .CLK(\fpu_add_exp_dp/n448 ), 
        .Q(\fpu_add_exp_dp/a4stg_exp_pre2[6] ), .QN(\fpu_add_exp_dp/n70 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[6]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N9 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[6] ), .QN(\fpu_add_exp_dp/n71 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[5]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N8 ), .CLK(\fpu_add_exp_dp/n448 ), 
        .Q(\fpu_add_exp_dp/a4stg_exp_pre2[5] ), .QN(\fpu_add_exp_dp/n72 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[5]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N8 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[5] ), .QN(\fpu_add_exp_dp/n73 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[4]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N7 ), .CLK(\fpu_add_exp_dp/n448 ), 
        .Q(\fpu_add_exp_dp/a4stg_exp_pre2[4] ), .QN(\fpu_add_exp_dp/n74 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[4]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N7 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[4] ), .QN(\fpu_add_exp_dp/n75 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[3]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N6 ), .CLK(\fpu_add_exp_dp/n448 ), 
        .Q(\fpu_add_exp_dp/a4stg_exp_pre2[3] ), .QN(\fpu_add_exp_dp/n76 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[3]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N6 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[3] ), .QN(\fpu_add_exp_dp/n77 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[2]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N5 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre2[2] ), .QN(\fpu_add_exp_dp/n78 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[2]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N5 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[2] ), .QN(\fpu_add_exp_dp/n79 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[1]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N4 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre2[1] ), .QN(\fpu_add_exp_dp/n80 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[1]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N4 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[1] ), .QN(\fpu_add_exp_dp/n81 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre2/q_reg[0]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre2/N3 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre2[0] ), .QN(\fpu_add_exp_dp/n82 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre4/q_reg[0]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N3 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre4[0] ), .QN(\fpu_add_exp_dp/n83 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[11]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N14 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[11] ), .QN(\fpu_add_exp_dp/n85 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[10]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N13 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[10] ), .QN(\fpu_add_exp_dp/n86 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[9]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N12 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[9] ), .QN(\fpu_add_exp_dp/n87 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[8]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N11 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[8] ), .QN(\fpu_add_exp_dp/n88 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[7]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N10 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[7] ), .QN(\fpu_add_exp_dp/n89 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[6]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N9 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[6] ), .QN(\fpu_add_exp_dp/n90 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[5]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N8 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[5] ), .QN(\fpu_add_exp_dp/n91 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[4]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N7 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[4] ), .QN(\fpu_add_exp_dp/n92 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[3]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N6 ), .CLK(n1568), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[3] ), .QN(\fpu_add_exp_dp/n93 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[2]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N5 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[2] ), .QN(\fpu_add_exp_dp/n94 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[1]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N4 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[1] ), .QN(\fpu_add_exp_dp/n95 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre3/q_reg[0]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N3 ), .CLK(n1569), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre3[0] ), .QN(\fpu_add_exp_dp/n96 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[11]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N14 ), .CLK(n1571), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[11] ), .QN(\fpu_add_exp_dp/n98 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[10]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N13 ), .CLK(n1571), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[10] ), .QN(\fpu_add_exp_dp/n99 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[9]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N12 ), .CLK(n1571), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[9] ), .QN(\fpu_add_exp_dp/n100 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[8]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N11 ), .CLK(n1571), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[8] ), .QN(\fpu_add_exp_dp/n101 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[7]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N10 ), .CLK(n1571), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[7] ), .QN(\fpu_add_exp_dp/n102 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[6]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N9 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[6] ), .QN(\fpu_add_exp_dp/n103 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[5]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N8 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[5] ), .QN(\fpu_add_exp_dp/n104 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[4]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N7 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[4] ), .QN(\fpu_add_exp_dp/n105 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[3]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N6 ), .CLK(n1570), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[3] ), .QN(\fpu_add_exp_dp/n106 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[2]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N5 ), .CLK(n1571), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[2] ), .QN(\fpu_add_exp_dp/n107 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[1]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N4 ), .CLK(n1571), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[1] ), .QN(\fpu_add_exp_dp/n108 ) );
  DFFX1 \fpu_add_exp_dp/i_a4stg_exp_pre1/q_reg[0]  ( .D(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N3 ), .CLK(n1571), .Q(
        \fpu_add_exp_dp/a4stg_exp_pre1[0] ), .QN(\fpu_add_exp_dp/n109 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[11]  ( .D(\fpu_add_exp_dp/n565 ), 
        .CLK(n1575), .Q(n728), .QN(\fpu_add_exp_dp/n447 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[10]  ( .D(\fpu_add_exp_dp/n566 ), 
        .CLK(n1573), .Q(n181), .QN(\fpu_add_exp_dp/n446 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[9]  ( .D(\fpu_add_exp_dp/n567 ), 
        .CLK(n1573), .Q(n17), .QN(\fpu_add_exp_dp/n443 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[8]  ( .D(\fpu_add_exp_dp/n568 ), 
        .CLK(n1573), .Q(n71), .QN(\fpu_add_exp_dp/n445 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[7]  ( .D(\fpu_add_exp_dp/n569 ), 
        .CLK(n1572), .Q(n256), .QN(\fpu_add_exp_dp/n442 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[6]  ( .D(\fpu_add_exp_dp/n570 ), 
        .CLK(n1573), .Q(n160), .QN(\fpu_add_exp_dp/n435 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[5]  ( .D(\fpu_add_exp_dp/n571 ), 
        .CLK(n1572), .Q(n69), .QN(\fpu_add_exp_dp/n433 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[4]  ( .D(\fpu_add_exp_dp/n572 ), 
        .CLK(n1572), .Q(n67), .QN(\fpu_add_exp_dp/n432 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[3]  ( .D(\fpu_add_exp_dp/n573 ), 
        .CLK(n1572), .Q(n178), .QN(\fpu_add_exp_dp/n434 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[2]  ( .D(\fpu_add_exp_dp/n574 ), 
        .CLK(n1572), .Q(n159), .QN(\fpu_add_exp_dp/n431 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[1]  ( .D(\fpu_add_exp_dp/n575 ), 
        .CLK(n1572), .Q(n72), .QN(\fpu_add_exp_dp/n436 ) );
  DFFX1 \fpu_add_exp_dp/i_a3stg_exp/q_reg[0]  ( .D(\fpu_add_exp_dp/n576 ), 
        .CLK(n1573), .Q(n583), .QN(\fpu_add_exp_dp/n444 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[12]  ( .D(
        \fpu_add_exp_dp/n577 ), .CLK(n1576), .Q(n694) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[11]  ( .D(
        \fpu_add_exp_dp/n578 ), .CLK(n1576), .Q(n629), .QN(
        \fpu_add_exp_dp/n111 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[10]  ( .D(
        \fpu_add_exp_dp/n579 ), .CLK(n1576), .Q(n298), .QN(
        \fpu_add_exp_dp/n112 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[9]  ( .D(
        \fpu_add_exp_dp/n580 ), .CLK(n1576), .Q(n300), .QN(
        \fpu_add_exp_dp/n113 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[8]  ( .D(
        \fpu_add_exp_dp/n581 ), .CLK(n1576), .Q(n301), .QN(
        \fpu_add_exp_dp/n114 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[7]  ( .D(
        \fpu_add_exp_dp/n582 ), .CLK(n1576), .Q(n308), .QN(
        \fpu_add_exp_dp/n115 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[6]  ( .D(
        \fpu_add_exp_dp/n583 ), .CLK(n1576), .Q(n302), .QN(
        \fpu_add_exp_dp/n116 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[5]  ( .D(
        \fpu_add_exp_dp/n584 ), .CLK(n1576), .Q(n299), .QN(
        \fpu_add_exp_dp/n117 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[4]  ( .D(
        \fpu_add_exp_dp/n585 ), .CLK(n1576), .Q(n303), .QN(
        \fpu_add_exp_dp/n118 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[3]  ( .D(
        \fpu_add_exp_dp/n586 ), .CLK(n1575), .Q(n304), .QN(
        \fpu_add_exp_dp/n119 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[2]  ( .D(
        \fpu_add_exp_dp/n587 ), .CLK(n1575), .Q(n305), .QN(
        \fpu_add_exp_dp/n120 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[1]  ( .D(
        \fpu_add_exp_dp/n588 ), .CLK(n1575), .Q(n297), .QN(
        \fpu_add_exp_dp/n121 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expadd2_in2/q_reg[0]  ( .D(
        \fpu_add_exp_dp/n589 ), .CLK(n1575), .Q(n830), .QN(
        \fpu_add_exp_dp/n122 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[11]  ( .D(\fpu_add_exp_dp/n591 ), 
        .CLK(n1575), .Q(n316), .QN(\fpu_add_exp_dp/n124 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[10]  ( .D(\fpu_add_exp_dp/n592 ), 
        .CLK(n1575), .Q(n680), .QN(\fpu_add_exp_dp/n125 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[9]  ( .D(\fpu_add_exp_dp/n593 ), 
        .CLK(n1575), .Q(n681), .QN(\fpu_add_exp_dp/n126 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[8]  ( .D(\fpu_add_exp_dp/n594 ), 
        .CLK(n1575), .Q(n682), .QN(\fpu_add_exp_dp/n127 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[7]  ( .D(\fpu_add_exp_dp/n595 ), 
        .CLK(n1575), .Q(n683), .QN(\fpu_add_exp_dp/n128 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[6]  ( .D(\fpu_add_exp_dp/n596 ), 
        .CLK(n1575), .Q(n661), .QN(\fpu_add_exp_dp/n129 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[5]  ( .D(\fpu_add_exp_dp/n597 ), 
        .CLK(n1575), .Q(n684), .QN(\fpu_add_exp_dp/n130 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[4]  ( .D(\fpu_add_exp_dp/n598 ), 
        .CLK(n1574), .Q(n685), .QN(\fpu_add_exp_dp/n131 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[3]  ( .D(\fpu_add_exp_dp/n599 ), 
        .CLK(n1574), .Q(n686), .QN(\fpu_add_exp_dp/n132 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[2]  ( .D(\fpu_add_exp_dp/n600 ), 
        .CLK(n1574), .Q(n687), .QN(\fpu_add_exp_dp/n133 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[1]  ( .D(\fpu_add_exp_dp/n601 ), 
        .CLK(n1574), .Q(n676), .QN(\fpu_add_exp_dp/n134 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_expa/q_reg[0]  ( .D(\fpu_add_exp_dp/n602 ), 
        .CLK(n1574), .Q(n315), .QN(\fpu_add_exp_dp/n135 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[11]  ( .D(\fpu_add_exp_dp/n603 ), 
        .CLK(n1574), .Q(n725), .QN(\fpu_add_exp_dp/n136 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[10]  ( .D(\fpu_add_exp_dp/n604 ), 
        .CLK(n1574), .Q(n289), .QN(\fpu_add_exp_dp/n137 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[9]  ( .D(\fpu_add_exp_dp/n605 ), 
        .CLK(n1574), .Q(n88) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[8]  ( .D(\fpu_add_exp_dp/n606 ), 
        .CLK(n1574), .Q(n35) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[7]  ( .D(\fpu_add_exp_dp/n607 ), 
        .CLK(n1574), .Q(n221) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[6]  ( .D(\fpu_add_exp_dp/n608 ), 
        .CLK(n1574), .Q(n711), .QN(\fpu_add_exp_dp/n141 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[5]  ( .D(\fpu_add_exp_dp/n609 ), 
        .CLK(n1574), .Q(n646), .QN(\fpu_add_exp_dp/n142 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[4]  ( .D(\fpu_add_exp_dp/n610 ), 
        .CLK(n1573), .Q(n648), .QN(\fpu_add_exp_dp/n143 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[3]  ( .D(\fpu_add_exp_dp/n611 ), 
        .CLK(n1573), .Q(n290), .QN(\fpu_add_exp_dp/n144 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[2]  ( .D(\fpu_add_exp_dp/n612 ), 
        .CLK(n1573), .Q(n287), .QN(\fpu_add_exp_dp/n145 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[1]  ( .D(\fpu_add_exp_dp/n613 ), 
        .CLK(n1573), .Q(n73), .QN(\fpu_add_exp_dp/n146 ) );
  DFFX1 \fpu_add_exp_dp/i_a2stg_exp/q_reg[0]  ( .D(\fpu_add_exp_dp/n614 ), 
        .CLK(n1573), .Q(n645), .QN(\fpu_add_exp_dp/n147 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[10]  ( .D(
        \fpu_add_exp_dp/n615 ), .CLK(n1577), .Q(
        \fpu_add_exp_dp/a1stg_expadd3_in2[10] ), .QN(\fpu_add_exp_dp/n47 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[9]  ( .D(
        \fpu_add_exp_dp/n616 ), .CLK(n1577), .Q(n445), .QN(
        \fpu_add_exp_dp/n149 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[8]  ( .D(
        \fpu_add_exp_dp/n617 ), .CLK(n1577), .Q(n446), .QN(
        \fpu_add_exp_dp/n150 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[7]  ( .D(
        \fpu_add_exp_dp/n618 ), .CLK(n1585), .Q(n323) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[6]  ( .D(
        \fpu_add_exp_dp/n619 ), .CLK(n1585), .Q(n322) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[5]  ( .D(
        \fpu_add_exp_dp/n620 ), .CLK(n1585), .Q(n321) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[4]  ( .D(
        \fpu_add_exp_dp/n621 ), .CLK(n1585), .Q(n320) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[3]  ( .D(
        \fpu_add_exp_dp/n622 ), .CLK(n1585), .Q(n319) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[2]  ( .D(
        \fpu_add_exp_dp/n623 ), .CLK(n1585), .Q(n309) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[1]  ( .D(
        \fpu_add_exp_dp/n624 ), .CLK(n1585), .Q(n56) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in2/q_reg[0]  ( .D(
        \fpu_add_exp_dp/n625 ), .CLK(n1585), .Q(n491) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[10]  ( .D(
        \fpu_add_exp_dp/n626 ), .CLK(n1585), .Q(n961), .QN(
        \fpu_add_exp_dp/n45 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[9]  ( .D(
        \fpu_add_exp_dp/n627 ), .CLK(n1584), .Q(n1000) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[8]  ( .D(
        \fpu_add_exp_dp/n628 ), .CLK(n1584), .Q(n999) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[7]  ( .D(
        \fpu_add_exp_dp/n629 ), .CLK(n1584), .Q(n998) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[6]  ( .D(
        \fpu_add_exp_dp/n630 ), .CLK(n1584), .Q(n997) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[5]  ( .D(
        \fpu_add_exp_dp/n631 ), .CLK(n1584), .Q(n996) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[4]  ( .D(
        \fpu_add_exp_dp/n632 ), .CLK(n1584), .Q(n995) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[3]  ( .D(
        \fpu_add_exp_dp/n633 ), .CLK(n1584), .Q(n994) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[2]  ( .D(
        \fpu_add_exp_dp/n634 ), .CLK(n1584), .Q(n993) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[1]  ( .D(
        \fpu_add_exp_dp/n635 ), .CLK(n1584), .Q(n138) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_expadd3_in1/q_reg[0]  ( .D(
        \fpu_add_exp_dp/n636 ), .CLK(n1584), .Q(n992) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_op_7/q_reg[3]  ( .D(\fpu_add_exp_dp/n637 ), 
        .CLK(n1584), .Q(n1241), .QN(\fpu_add_exp_dp/n170 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_op_7/q_reg[2]  ( .D(\fpu_add_exp_dp/n638 ), 
        .CLK(n1584), .Q(n1240), .QN(\fpu_add_exp_dp/n171 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_op_7/q_reg[1]  ( .D(\fpu_add_exp_dp/n639 ), 
        .CLK(n1583), .Q(n1239), .QN(\fpu_add_exp_dp/n172 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_op_7/q_reg[0]  ( .D(\fpu_add_exp_dp/n640 ), 
        .CLK(n1583), .Q(n13) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[10]  ( .D(
        \fpu_add_exp_dp/n641 ), .CLK(n1583), .Q(n1148), .QN(
        \fpu_add_exp_dp/n174 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[9]  ( .D(\fpu_add_exp_dp/n642 ), .CLK(n1583), .Q(n559), .QN(\fpu_add_exp_dp/n175 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[8]  ( .D(\fpu_add_exp_dp/n643 ), .CLK(n1583), .Q(n1163), .QN(\fpu_add_exp_dp/n176 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[7]  ( .D(\fpu_add_exp_dp/n644 ), .CLK(n1583), .Q(n1171), .QN(\fpu_add_exp_dp/n177 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[6]  ( .D(\fpu_add_exp_dp/n645 ), .CLK(n1583), .Q(n1168), .QN(\fpu_add_exp_dp/n178 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[5]  ( .D(\fpu_add_exp_dp/n646 ), .CLK(n1583), .Q(n1155), .QN(\fpu_add_exp_dp/n179 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[4]  ( .D(\fpu_add_exp_dp/n647 ), .CLK(n1583), .Q(n1167), .QN(\fpu_add_exp_dp/n180 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[3]  ( .D(\fpu_add_exp_dp/n648 ), .CLK(n1583), .Q(n1166), .QN(\fpu_add_exp_dp/n181 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[2]  ( .D(\fpu_add_exp_dp/n649 ), .CLK(n1583), .Q(n1179), .QN(\fpu_add_exp_dp/n182 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[1]  ( .D(\fpu_add_exp_dp/n650 ), .CLK(n1583), .Q(n558), .QN(\fpu_add_exp_dp/n183 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblopa/q_reg[0]  ( .D(\fpu_add_exp_dp/n651 ), .CLK(n1582), .Q(n151), .QN(\fpu_add_exp_dp/n184 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[10]  ( .D(\fpu_add_exp_dp/n652 ), .CLK(n1582), .Q(n928), .QN(\fpu_add_exp_dp/n185 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[9]  ( .D(\fpu_add_exp_dp/n653 ), 
        .CLK(n1582), .Q(n1150), .QN(\fpu_add_exp_dp/n186 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[8]  ( .D(\fpu_add_exp_dp/n654 ), 
        .CLK(n1582), .Q(n1147), .QN(\fpu_add_exp_dp/n187 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[7]  ( .D(\fpu_add_exp_dp/n655 ), 
        .CLK(n1582), .Q(n545), .QN(\fpu_add_exp_dp/n188 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[6]  ( .D(\fpu_add_exp_dp/n656 ), 
        .CLK(n1582), .Q(n546), .QN(\fpu_add_exp_dp/n189 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[5]  ( .D(\fpu_add_exp_dp/n657 ), 
        .CLK(n1582), .Q(n516), .QN(\fpu_add_exp_dp/n190 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[4]  ( .D(\fpu_add_exp_dp/n658 ), 
        .CLK(n1582), .Q(n515), .QN(\fpu_add_exp_dp/n191 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[3]  ( .D(\fpu_add_exp_dp/n659 ), 
        .CLK(n1582), .Q(n514), .QN(\fpu_add_exp_dp/n192 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[2]  ( .D(\fpu_add_exp_dp/n660 ), 
        .CLK(n1582), .Q(n1165), .QN(\fpu_add_exp_dp/n193 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[1]  ( .D(\fpu_add_exp_dp/n661 ), 
        .CLK(n1582), .Q(n1154), .QN(\fpu_add_exp_dp/n194 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_dblop/q_reg[0]  ( .D(\fpu_add_exp_dp/n662 ), 
        .CLK(n1582), .Q(n1164), .QN(\fpu_add_exp_dp/n195 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngopa/q_reg[7]  ( .D(\fpu_add_exp_dp/n663 ), .CLK(n1581), .Q(n1178), .QN(\fpu_add_exp_dp/n196 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngopa/q_reg[6]  ( .D(\fpu_add_exp_dp/n664 ), .CLK(n1581), .Q(n1177), .QN(\fpu_add_exp_dp/n197 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngopa/q_reg[5]  ( .D(\fpu_add_exp_dp/n665 ), .CLK(n1581), .Q(n1170), .QN(\fpu_add_exp_dp/n198 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngopa/q_reg[4]  ( .D(\fpu_add_exp_dp/n666 ), .CLK(n1581), .Q(n1176), .QN(\fpu_add_exp_dp/n199 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngopa/q_reg[3]  ( .D(\fpu_add_exp_dp/n667 ), .CLK(n1581), .Q(n1175), .QN(\fpu_add_exp_dp/n200 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngopa/q_reg[2]  ( .D(\fpu_add_exp_dp/n668 ), .CLK(n1581), .Q(n1174), .QN(\fpu_add_exp_dp/n201 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngopa/q_reg[1]  ( .D(\fpu_add_exp_dp/n669 ), .CLK(n1581), .Q(n61), .QN(\fpu_add_exp_dp/n202 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngopa/q_reg[0]  ( .D(\fpu_add_exp_dp/n670 ), .CLK(n1581), .Q(n510), .QN(\fpu_add_exp_dp/n203 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngop/q_reg[7]  ( .D(\fpu_add_exp_dp/n671 ), 
        .CLK(n1581), .Q(n936), .QN(\fpu_add_exp_dp/n204 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngop/q_reg[6]  ( .D(\fpu_add_exp_dp/n672 ), 
        .CLK(n1581), .Q(n937), .QN(\fpu_add_exp_dp/n205 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngop/q_reg[5]  ( .D(\fpu_add_exp_dp/n673 ), 
        .CLK(n1581), .Q(n960), .QN(\fpu_add_exp_dp/n206 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngop/q_reg[4]  ( .D(\fpu_add_exp_dp/n674 ), 
        .CLK(n1581), .Q(n959), .QN(\fpu_add_exp_dp/n207 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngop/q_reg[3]  ( .D(\fpu_add_exp_dp/n675 ), 
        .CLK(n1580), .Q(n958), .QN(\fpu_add_exp_dp/n208 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngop/q_reg[2]  ( .D(\fpu_add_exp_dp/n676 ), 
        .CLK(n1580), .Q(n1160), .QN(\fpu_add_exp_dp/n209 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngop/q_reg[1]  ( .D(\fpu_add_exp_dp/n677 ), 
        .CLK(n1580), .Q(n1169), .QN(\fpu_add_exp_dp/n210 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_dp_sngop/q_reg[0]  ( .D(\fpu_add_exp_dp/n678 ), 
        .CLK(n1580), .Q(n1159), .QN(\fpu_add_exp_dp/n211 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[10]  ( .D(\fpu_add_exp_dp/n679 ), 
        .CLK(n1580), .Q(n1181), .QN(\fpu_add_exp_dp/n212 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[9]  ( .D(\fpu_add_exp_dp/n680 ), 
        .CLK(n1580), .Q(n1075), .QN(\fpu_add_exp_dp/n213 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[8]  ( .D(\fpu_add_exp_dp/n681 ), 
        .CLK(n1580), .Q(n1180), .QN(\fpu_add_exp_dp/n214 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[7]  ( .D(\fpu_add_exp_dp/n682 ), 
        .CLK(n1577), .Q(\fpu_add_exp_dp/a1stg_in2a[59] ), .QN(
        \fpu_add_exp_dp/n215 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[6]  ( .D(\fpu_add_exp_dp/n683 ), 
        .CLK(n1577), .Q(\fpu_add_exp_dp/a1stg_in2a[58] ), .QN(
        \fpu_add_exp_dp/n216 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[5]  ( .D(\fpu_add_exp_dp/n684 ), 
        .CLK(n1577), .Q(\fpu_add_exp_dp/a1stg_in2a[57] ), .QN(
        \fpu_add_exp_dp/n217 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[4]  ( .D(\fpu_add_exp_dp/n685 ), 
        .CLK(n1577), .Q(\fpu_add_exp_dp/a1stg_in2a[56] ), .QN(
        \fpu_add_exp_dp/n218 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[3]  ( .D(\fpu_add_exp_dp/n686 ), 
        .CLK(n1577), .Q(\fpu_add_exp_dp/a1stg_in2a[55] ), .QN(
        \fpu_add_exp_dp/n219 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[2]  ( .D(\fpu_add_exp_dp/n687 ), 
        .CLK(n1576), .Q(\fpu_add_exp_dp/a1stg_in2a[54] ), .QN(
        \fpu_add_exp_dp/n220 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[1]  ( .D(\fpu_add_exp_dp/n688 ), 
        .CLK(n1576), .Q(\fpu_add_exp_dp/a1stg_in2a[53] ), .QN(
        \fpu_add_exp_dp/n221 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2a/q_reg[0]  ( .D(\fpu_add_exp_dp/n689 ), 
        .CLK(n1576), .Q(\fpu_add_exp_dp/a1stg_in2a[52] ), .QN(
        \fpu_add_exp_dp/n222 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[10]  ( .D(\fpu_add_exp_dp/n690 ), 
        .CLK(n1580), .Q(n105) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[9]  ( .D(\fpu_add_exp_dp/n691 ), 
        .CLK(n1580), .Q(n127), .QN(\fpu_add_exp_dp/n224 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[8]  ( .D(\fpu_add_exp_dp/n692 ), 
        .CLK(n1580), .Q(n126), .QN(\fpu_add_exp_dp/n225 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[7]  ( .D(\fpu_add_exp_dp/n693 ), 
        .CLK(n1580), .Q(n41) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[6]  ( .D(\fpu_add_exp_dp/n694 ), 
        .CLK(n1580), .Q(n42) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[5]  ( .D(\fpu_add_exp_dp/n695 ), 
        .CLK(n1579), .Q(n49), .QN(\fpu_add_exp_dp/n228 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[4]  ( .D(\fpu_add_exp_dp/n696 ), 
        .CLK(n1579), .Q(n110), .QN(\fpu_add_exp_dp/n229 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[3]  ( .D(\fpu_add_exp_dp/n697 ), 
        .CLK(n1579), .Q(n109), .QN(\fpu_add_exp_dp/n230 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[2]  ( .D(\fpu_add_exp_dp/n698 ), 
        .CLK(n1579), .Q(n1005), .QN(\fpu_add_exp_dp/n231 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[1]  ( .D(\fpu_add_exp_dp/n699 ), 
        .CLK(n1579), .Q(n991), .QN(\fpu_add_exp_dp/n232 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in2/q_reg[0]  ( .D(\fpu_add_exp_dp/n700 ), 
        .CLK(n1579), .Q(n990), .QN(\fpu_add_exp_dp/n233 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[10]  ( .D(\fpu_add_exp_dp/n701 ), 
        .CLK(n1579), .Q(n657), .QN(\fpu_add_exp_dp/n234 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[9]  ( .D(\fpu_add_exp_dp/n702 ), 
        .CLK(n1579), .Q(n656), .QN(\fpu_add_exp_dp/n235 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[8]  ( .D(\fpu_add_exp_dp/n703 ), 
        .CLK(n1579), .Q(n658), .QN(\fpu_add_exp_dp/n236 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[7]  ( .D(\fpu_add_exp_dp/n704 ), 
        .CLK(n1579), .Q(n669), .QN(\fpu_add_exp_dp/n237 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[6]  ( .D(\fpu_add_exp_dp/n705 ), 
        .CLK(n1579), .Q(n668), .QN(\fpu_add_exp_dp/n238 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[5]  ( .D(\fpu_add_exp_dp/n706 ), 
        .CLK(n1579), .Q(n675), .QN(\fpu_add_exp_dp/n239 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[4]  ( .D(\fpu_add_exp_dp/n707 ), 
        .CLK(n1578), .Q(n674), .QN(\fpu_add_exp_dp/n240 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[3]  ( .D(\fpu_add_exp_dp/n708 ), 
        .CLK(n1578), .Q(n672), .QN(\fpu_add_exp_dp/n241 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[2]  ( .D(\fpu_add_exp_dp/n709 ), 
        .CLK(n1578), .Q(n508), .QN(\fpu_add_exp_dp/n242 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[1]  ( .D(\fpu_add_exp_dp/n710 ), 
        .CLK(n1578), .Q(n507), .QN(\fpu_add_exp_dp/n243 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1a/q_reg[0]  ( .D(\fpu_add_exp_dp/n711 ), 
        .CLK(n1578), .Q(n509), .QN(\fpu_add_exp_dp/n244 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[10]  ( .D(\fpu_add_exp_dp/n712 ), 
        .CLK(n1578), .Q(n1156), .QN(\fpu_add_exp_dp/n245 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[9]  ( .D(\fpu_add_exp_dp/n713 ), 
        .CLK(n1578), .Q(n1183), .QN(\fpu_add_exp_dp/n246 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[8]  ( .D(\fpu_add_exp_dp/n714 ), 
        .CLK(n1578), .Q(n1182), .QN(\fpu_add_exp_dp/n247 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[7]  ( .D(\fpu_add_exp_dp/n715 ), 
        .CLK(n1578), .Q(n1172), .QN(\fpu_add_exp_dp/n248 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[6]  ( .D(\fpu_add_exp_dp/n716 ), 
        .CLK(n1578), .Q(n1162), .QN(\fpu_add_exp_dp/n249 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[5]  ( .D(\fpu_add_exp_dp/n717 ), 
        .CLK(n1578), .Q(n1161), .QN(\fpu_add_exp_dp/n250 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[4]  ( .D(\fpu_add_exp_dp/n718 ), 
        .CLK(n1578), .Q(n152), .QN(\fpu_add_exp_dp/n251 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[3]  ( .D(\fpu_add_exp_dp/n719 ), 
        .CLK(n1577), .Q(n60), .QN(\fpu_add_exp_dp/n252 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[2]  ( .D(\fpu_add_exp_dp/n720 ), 
        .CLK(n1577), .Q(n1223), .QN(\fpu_add_exp_dp/n253 ) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[1]  ( .D(\fpu_add_exp_dp/n721 ), 
        .CLK(n1577), .Q(n1066) );
  DFFX1 \fpu_add_exp_dp/i_a1stg_in1/q_reg[0]  ( .D(\fpu_add_exp_dp/n722 ), 
        .CLK(n1577), .Q(n1033) );
  LATCHX1 \fpu_add_exp_dp/ckbuf_add_exp_dp/clken_reg  ( .CLK(
        \fpu_add_frac_dp/n2189 ), .D(\fpu_add_exp_dp/ckbuf_add_exp_dp/N1 ), 
        .Q(\fpu_add_exp_dp/ckbuf_add_exp_dp/clken ), .QN(\fpu_add_exp_dp/n256 ) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[63]  ( .D(\fpu_add_frac_dp/n3375 ), 
        .CLK(n1529), .Q(n467) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[62]  ( .D(\fpu_add_frac_dp/n3376 ), 
        .CLK(n1529), .Q(n468) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[61]  ( .D(\fpu_add_frac_dp/n3377 ), 
        .CLK(n1529), .Q(n963) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[60]  ( .D(\fpu_add_frac_dp/n3378 ), 
        .CLK(n1528), .Q(n466) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[59]  ( .D(\fpu_add_frac_dp/n3379 ), 
        .CLK(n1528), .Q(n933) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[58]  ( .D(\fpu_add_frac_dp/n3380 ), 
        .CLK(n1529), .Q(n1034) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[57]  ( .D(\fpu_add_frac_dp/n3381 ), 
        .CLK(n1528), .Q(n906) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[56]  ( .D(\fpu_add_frac_dp/n3382 ), 
        .CLK(n1530), .Q(n1064) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[55]  ( .D(\fpu_add_frac_dp/n3383 ), 
        .CLK(n1536), .Q(n918) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[54]  ( .D(\fpu_add_frac_dp/n3384 ), 
        .CLK(n1536), .Q(n909) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[53]  ( .D(\fpu_add_frac_dp/n3385 ), 
        .CLK(n1530), .Q(n910) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[52]  ( .D(\fpu_add_frac_dp/n3386 ), 
        .CLK(n1531), .Q(n911) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[51]  ( .D(\fpu_add_frac_dp/n3387 ), 
        .CLK(n1531), .Q(n912) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[50]  ( .D(\fpu_add_frac_dp/n3388 ), 
        .CLK(n1531), .Q(n913) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[49]  ( .D(\fpu_add_frac_dp/n3389 ), 
        .CLK(n1526), .Q(n469) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[48]  ( .D(\fpu_add_frac_dp/n3390 ), 
        .CLK(n1525), .Q(n470) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[47]  ( .D(\fpu_add_frac_dp/n3391 ), 
        .CLK(n1525), .Q(n471) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[46]  ( .D(\fpu_add_frac_dp/n3392 ), 
        .CLK(n1525), .Q(n472) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[45]  ( .D(\fpu_add_frac_dp/n3393 ), 
        .CLK(n1525), .Q(n473) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[44]  ( .D(\fpu_add_frac_dp/n3394 ), 
        .CLK(n1524), .Q(n474) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[43]  ( .D(\fpu_add_frac_dp/n3395 ), 
        .CLK(n1524), .Q(n475) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[42]  ( .D(\fpu_add_frac_dp/n3396 ), 
        .CLK(n1524), .Q(n476) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[41]  ( .D(\fpu_add_frac_dp/n3397 ), 
        .CLK(n1524), .Q(n477) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[40]  ( .D(\fpu_add_frac_dp/n3398 ), 
        .CLK(n1524), .Q(n478) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[39]  ( .D(\fpu_add_frac_dp/n3399 ), 
        .CLK(n1523), .Q(n479) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[38]  ( .D(\fpu_add_frac_dp/n3400 ), 
        .CLK(n1523), .Q(n480) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[37]  ( .D(\fpu_add_frac_dp/n3401 ), 
        .CLK(n1523), .Q(n481) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[36]  ( .D(\fpu_add_frac_dp/n3402 ), 
        .CLK(n1523), .Q(n482) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[35]  ( .D(\fpu_add_frac_dp/n3403 ), 
        .CLK(n1522), .Q(n483) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[34]  ( .D(\fpu_add_frac_dp/n3404 ), 
        .CLK(n1522), .Q(n484) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[33]  ( .D(\fpu_add_frac_dp/n3405 ), 
        .CLK(n1521), .Q(n485) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[32]  ( .D(\fpu_add_frac_dp/n3406 ), 
        .CLK(n1521), .Q(n486) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[31]  ( .D(\fpu_add_frac_dp/n3407 ), 
        .CLK(n1521), .Q(n487) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[30]  ( .D(\fpu_add_frac_dp/n3408 ), 
        .CLK(n1521), .Q(n488) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[29]  ( .D(\fpu_add_frac_dp/n3409 ), 
        .CLK(n1521), .Q(n489) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[28]  ( .D(\fpu_add_frac_dp/n3410 ), 
        .CLK(n1520), .Q(n517) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[27]  ( .D(\fpu_add_frac_dp/n3411 ), 
        .CLK(n1520), .Q(n518) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[26]  ( .D(\fpu_add_frac_dp/n3412 ), 
        .CLK(n1520), .Q(n519) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[25]  ( .D(\fpu_add_frac_dp/n3413 ), 
        .CLK(n1520), .Q(n520) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[24]  ( .D(\fpu_add_frac_dp/n3414 ), 
        .CLK(n1537), .Q(n521) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[23]  ( .D(\fpu_add_frac_dp/n3415 ), 
        .CLK(n1538), .Q(n522) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[22]  ( .D(\fpu_add_frac_dp/n3416 ), 
        .CLK(n1538), .Q(n523) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[21]  ( .D(\fpu_add_frac_dp/n3417 ), 
        .CLK(n1518), .Q(n524) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[20]  ( .D(\fpu_add_frac_dp/n3418 ), 
        .CLK(n1519), .Q(n525) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[19]  ( .D(\fpu_add_frac_dp/n3419 ), 
        .CLK(n1519), .Q(n526) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[18]  ( .D(\fpu_add_frac_dp/n3420 ), 
        .CLK(n1519), .Q(n527) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[17]  ( .D(\fpu_add_frac_dp/n3421 ), 
        .CLK(n1537), .Q(n528) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[16]  ( .D(\fpu_add_frac_dp/n3422 ), 
        .CLK(n1537), .Q(n529) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[15]  ( .D(\fpu_add_frac_dp/n3423 ), 
        .CLK(n1532), .Q(n530) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[14]  ( .D(\fpu_add_frac_dp/n3424 ), 
        .CLK(n1535), .Q(n531) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[13]  ( .D(\fpu_add_frac_dp/n3425 ), 
        .CLK(n1535), .Q(n532) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[12]  ( .D(\fpu_add_frac_dp/n3426 ), 
        .CLK(n1536), .Q(n533) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[11]  ( .D(\fpu_add_frac_dp/n3427 ), 
        .CLK(n1519), .Q(n534) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[10]  ( .D(\fpu_add_frac_dp/n3428 ), 
        .CLK(n1519), .Q(n535) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[9]  ( .D(\fpu_add_frac_dp/n3429 ), 
        .CLK(n1537), .Q(n1002) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[8]  ( .D(\fpu_add_frac_dp/n3430 ), 
        .CLK(n1537), .Q(n1003) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[7]  ( .D(\fpu_add_frac_dp/n3431 ), 
        .CLK(n1531), .Q(n919) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[6]  ( .D(\fpu_add_frac_dp/n3432 ), 
        .CLK(n1535), .Q(n920) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[5]  ( .D(\fpu_add_frac_dp/n3433 ), 
        .CLK(n1535), .Q(n921) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[4]  ( .D(\fpu_add_frac_dp/n3434 ), 
        .CLK(n1536), .Q(n922) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[3]  ( .D(\fpu_add_frac_dp/n3435 ), 
        .CLK(n1522), .Q(n923) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[2]  ( .D(\fpu_add_frac_dp/n3436 ), 
        .CLK(n1522), .Q(n924) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[1]  ( .D(\fpu_add_frac_dp/n3437 ), 
        .CLK(n1522), .Q(n551) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_shl/q_reg[0]  ( .D(\fpu_add_frac_dp/n3438 ), 
        .CLK(n1522), .Q(n925) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[63]  ( .D(
        \fpu_add_frac_dp/n3439 ), .CLK(n1529), .Q(n859) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[62]  ( .D(
        \fpu_add_frac_dp/n3440 ), .CLK(n1529), .Q(n907) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[61]  ( .D(
        \fpu_add_frac_dp/n3441 ), .CLK(n1530), .Q(n493) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[60]  ( .D(
        \fpu_add_frac_dp/n3442 ), .CLK(n1533), .Q(n860) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[59]  ( .D(
        \fpu_add_frac_dp/n3443 ), .CLK(n1529), .Q(n494) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[58]  ( .D(
        \fpu_add_frac_dp/n3444 ), .CLK(n1529), .Q(n495) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[57]  ( .D(
        \fpu_add_frac_dp/n3445 ), .CLK(n1530), .Q(n496) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[56]  ( .D(
        \fpu_add_frac_dp/n3446 ), .CLK(n1530), .Q(n497) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[55]  ( .D(
        \fpu_add_frac_dp/n3447 ), .CLK(n1536), .Q(n498) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[54]  ( .D(
        \fpu_add_frac_dp/n3448 ), .CLK(n1536), .Q(n499) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[53]  ( .D(
        \fpu_add_frac_dp/n3449 ), .CLK(n1530), .Q(n500) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[52]  ( .D(
        \fpu_add_frac_dp/n3450 ), .CLK(n1531), .Q(n501) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[51]  ( .D(
        \fpu_add_frac_dp/n3451 ), .CLK(n1531), .Q(n502) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[50]  ( .D(
        \fpu_add_frac_dp/n3452 ), .CLK(n1531), .Q(n503) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[49]  ( .D(
        \fpu_add_frac_dp/n3453 ), .CLK(n1526), .Q(n861) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[48]  ( .D(
        \fpu_add_frac_dp/n3454 ), .CLK(n1525), .Q(n862) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[47]  ( .D(
        \fpu_add_frac_dp/n3455 ), .CLK(n1525), .Q(n863) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[46]  ( .D(
        \fpu_add_frac_dp/n3456 ), .CLK(n1525), .Q(n864) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[45]  ( .D(
        \fpu_add_frac_dp/n3457 ), .CLK(n1525), .Q(n865) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[44]  ( .D(
        \fpu_add_frac_dp/n3458 ), .CLK(n1525), .Q(n866) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[43]  ( .D(
        \fpu_add_frac_dp/n3459 ), .CLK(n1524), .Q(n867) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[42]  ( .D(
        \fpu_add_frac_dp/n3460 ), .CLK(n1524), .Q(n868) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[41]  ( .D(
        \fpu_add_frac_dp/n3461 ), .CLK(n1524), .Q(n869) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[40]  ( .D(
        \fpu_add_frac_dp/n3462 ), .CLK(n1524), .Q(n870) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[39]  ( .D(
        \fpu_add_frac_dp/n3463 ), .CLK(n1523), .Q(n871) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[38]  ( .D(
        \fpu_add_frac_dp/n3464 ), .CLK(n1523), .Q(n872) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[37]  ( .D(
        \fpu_add_frac_dp/n3465 ), .CLK(n1523), .Q(n873) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[36]  ( .D(
        \fpu_add_frac_dp/n3466 ), .CLK(n1523), .Q(n874) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[35]  ( .D(
        \fpu_add_frac_dp/n3467 ), .CLK(n1523), .Q(n875) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[34]  ( .D(
        \fpu_add_frac_dp/n3468 ), .CLK(n1522), .Q(n876) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[33]  ( .D(
        \fpu_add_frac_dp/n3469 ), .CLK(n1521), .Q(n877) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[32]  ( .D(
        \fpu_add_frac_dp/n3470 ), .CLK(n1521), .Q(n878) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[31]  ( .D(
        \fpu_add_frac_dp/n3471 ), .CLK(n1521), .Q(n879) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[30]  ( .D(
        \fpu_add_frac_dp/n3472 ), .CLK(n1521), .Q(n880) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[29]  ( .D(
        \fpu_add_frac_dp/n3473 ), .CLK(n1521), .Q(n881) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[28]  ( .D(
        \fpu_add_frac_dp/n3474 ), .CLK(n1520), .Q(n938) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[27]  ( .D(
        \fpu_add_frac_dp/n3475 ), .CLK(n1520), .Q(n939) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[26]  ( .D(
        \fpu_add_frac_dp/n3476 ), .CLK(n1520), .Q(n940) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[25]  ( .D(
        \fpu_add_frac_dp/n3477 ), .CLK(n1520), .Q(n941) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[24]  ( .D(
        \fpu_add_frac_dp/n3478 ), .CLK(n1537), .Q(n942) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[23]  ( .D(
        \fpu_add_frac_dp/n3479 ), .CLK(n1538), .Q(n943) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[22]  ( .D(
        \fpu_add_frac_dp/n3480 ), .CLK(n1523), .Q(n944) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[21]  ( .D(
        \fpu_add_frac_dp/n3481 ), .CLK(n1518), .Q(n945) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[20]  ( .D(
        \fpu_add_frac_dp/n3482 ), .CLK(n1519), .Q(n946) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[19]  ( .D(
        \fpu_add_frac_dp/n3483 ), .CLK(n1519), .Q(n947) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[18]  ( .D(
        \fpu_add_frac_dp/n3484 ), .CLK(n1519), .Q(n948) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[17]  ( .D(
        \fpu_add_frac_dp/n3485 ), .CLK(n1537), .Q(n949) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[16]  ( .D(
        \fpu_add_frac_dp/n3486 ), .CLK(n1537), .Q(n950) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[15]  ( .D(
        \fpu_add_frac_dp/n3487 ), .CLK(n1532), .Q(n951) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[14]  ( .D(
        \fpu_add_frac_dp/n3488 ), .CLK(n1535), .Q(n952) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[13]  ( .D(
        \fpu_add_frac_dp/n3489 ), .CLK(n1535), .Q(n953) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[12]  ( .D(
        \fpu_add_frac_dp/n3490 ), .CLK(n1536), .Q(n954) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[11]  ( .D(
        \fpu_add_frac_dp/n3491 ), .CLK(n1536), .Q(n955) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[10]  ( .D(
        \fpu_add_frac_dp/n3492 ), .CLK(n1519), .Q(n908) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[9]  ( .D(
        \fpu_add_frac_dp/n3493 ), .CLK(n1537), .Q(n536) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[8]  ( .D(
        \fpu_add_frac_dp/n3494 ), .CLK(n1537), .Q(n537) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[7]  ( .D(
        \fpu_add_frac_dp/n3495 ), .CLK(n1532), .Q(n538) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[6]  ( .D(
        \fpu_add_frac_dp/n3496 ), .CLK(n1535), .Q(n539) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[5]  ( .D(
        \fpu_add_frac_dp/n3497 ), .CLK(n1535), .Q(n540) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[4]  ( .D(
        \fpu_add_frac_dp/n3498 ), .CLK(n1536), .Q(n541) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[3]  ( .D(
        \fpu_add_frac_dp/n3499 ), .CLK(n1522), .Q(n542) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[2]  ( .D(
        \fpu_add_frac_dp/n3500 ), .CLK(n1522), .Q(n543) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[1]  ( .D(
        \fpu_add_frac_dp/n3501 ), .CLK(n1522), .Q(n978) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rnd_frac/q_reg[0]  ( .D(
        \fpu_add_frac_dp/n3502 ), .CLK(n1522), .Q(n544) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[57]  ( .D(
        \fpu_add_frac_dp/n3503 ), .CLK(n1528), .Q(n1248), .QN(
        \fpu_add_frac_dp/n129 ) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[56]  ( .D(
        \fpu_add_frac_dp/n3504 ), .CLK(n1532), .Q(n579) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[55]  ( .D(
        \fpu_add_frac_dp/n3505 ), .CLK(n1532), .Q(n66), .QN(
        \fpu_add_frac_dp/n5617 ) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[54]  ( .D(
        \fpu_add_frac_dp/n3506 ), .CLK(n1520), .Q(
        \fpu_add_frac_dp/a5stg_in_of ), .QN(\fpu_add_frac_dp/n132 ) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[53]  ( .D(
        \fpu_add_frac_dp/n3507 ), .CLK(n1520), .Q(n65), .QN(
        \fpu_add_frac_dp/n5616 ) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[52]  ( .D(
        \fpu_add_frac_dp/n3508 ), .CLK(n1555), .Q(n1186), .QN(
        \fpu_add_frac_dp/n134 ) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[51]  ( .D(
        \fpu_add_frac_dp/n3509 ), .CLK(n1528), .Q(n1006) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[50]  ( .D(
        \fpu_add_frac_dp/n3510 ), .CLK(n1538), .Q(n1035) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[49]  ( .D(
        \fpu_add_frac_dp/n3511 ), .CLK(n1481), .Q(n1036) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[48]  ( .D(
        \fpu_add_frac_dp/n3512 ), .CLK(n1529), .Q(n1037) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[47]  ( .D(
        \fpu_add_frac_dp/n3513 ), .CLK(n1529), .Q(n1038) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[46]  ( .D(
        \fpu_add_frac_dp/n3514 ), .CLK(n1530), .Q(n1039) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[45]  ( .D(
        \fpu_add_frac_dp/n3515 ), .CLK(n1530), .Q(n1040) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[44]  ( .D(
        \fpu_add_frac_dp/n3516 ), .CLK(n1530), .Q(n1041) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[43]  ( .D(
        \fpu_add_frac_dp/n3517 ), .CLK(n1530), .Q(n964) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[42]  ( .D(
        \fpu_add_frac_dp/n3518 ), .CLK(n1530), .Q(n965) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[41]  ( .D(
        \fpu_add_frac_dp/n3519 ), .CLK(n1531), .Q(n966) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[40]  ( .D(
        \fpu_add_frac_dp/n3520 ), .CLK(n1531), .Q(n967) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[39]  ( .D(
        \fpu_add_frac_dp/n3521 ), .CLK(n1531), .Q(n968) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[38]  ( .D(
        \fpu_add_frac_dp/n3522 ), .CLK(n1534), .Q(n1042) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[37]  ( .D(
        \fpu_add_frac_dp/n3523 ), .CLK(n1534), .Q(n1043) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[36]  ( .D(
        \fpu_add_frac_dp/n3524 ), .CLK(n1534), .Q(n1044) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[35]  ( .D(
        \fpu_add_frac_dp/n3525 ), .CLK(n1534), .Q(n1045) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[34]  ( .D(
        \fpu_add_frac_dp/n3526 ), .CLK(n1534), .Q(n1046) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[33]  ( .D(
        \fpu_add_frac_dp/n3527 ), .CLK(n1534), .Q(n1047) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[32]  ( .D(
        \fpu_add_frac_dp/n3528 ), .CLK(n1534), .Q(n1048) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[31]  ( .D(
        \fpu_add_frac_dp/n3529 ), .CLK(n1534), .Q(n1049) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[30]  ( .D(
        \fpu_add_frac_dp/n3530 ), .CLK(n1534), .Q(n1050) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[29]  ( .D(
        \fpu_add_frac_dp/n3531 ), .CLK(n1534), .Q(n1051) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[28]  ( .D(
        \fpu_add_frac_dp/n3532 ), .CLK(n1534), .Q(n1052) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[27]  ( .D(
        \fpu_add_frac_dp/n3533 ), .CLK(n1534), .Q(n1053) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[26]  ( .D(
        \fpu_add_frac_dp/n3534 ), .CLK(n1533), .Q(n1054) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[25]  ( .D(
        \fpu_add_frac_dp/n3535 ), .CLK(n1534), .Q(n1055) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[24]  ( .D(
        \fpu_add_frac_dp/n3536 ), .CLK(n1533), .Q(n1056) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[23]  ( .D(
        \fpu_add_frac_dp/n3537 ), .CLK(n1533), .Q(n1057) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[22]  ( .D(
        \fpu_add_frac_dp/n3538 ), .CLK(n1533), .Q(n1058) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[21]  ( .D(
        \fpu_add_frac_dp/n3539 ), .CLK(n1533), .Q(n1059) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[20]  ( .D(
        \fpu_add_frac_dp/n3540 ), .CLK(n1533), .Q(n1060) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[19]  ( .D(
        \fpu_add_frac_dp/n3541 ), .CLK(n1533), .Q(n1061) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[18]  ( .D(
        \fpu_add_frac_dp/n3542 ), .CLK(n1533), .Q(n1062) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[17]  ( .D(
        \fpu_add_frac_dp/n3543 ), .CLK(n1533), .Q(n969) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[16]  ( .D(
        \fpu_add_frac_dp/n3544 ), .CLK(n1533), .Q(n970) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[15]  ( .D(
        \fpu_add_frac_dp/n3545 ), .CLK(n1533), .Q(n971) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[14]  ( .D(
        \fpu_add_frac_dp/n3546 ), .CLK(n1533), .Q(n972) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[13]  ( .D(
        \fpu_add_frac_dp/n3547 ), .CLK(n1533), .Q(n973) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[12]  ( .D(
        \fpu_add_frac_dp/n3548 ), .CLK(n1532), .Q(n974) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[11]  ( .D(
        \fpu_add_frac_dp/n3549 ), .CLK(n1532), .Q(n975) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[10]  ( .D(
        \fpu_add_frac_dp/n3550 ), .CLK(n1532), .Q(n976) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[9]  ( .D(\fpu_add_frac_dp/n3551 ), .CLK(n1532), .Q(n977) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[8]  ( .D(\fpu_add_frac_dp/n3552 ), .CLK(n1532), .Q(n979) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[7]  ( .D(\fpu_add_frac_dp/n3553 ), .CLK(n1532), .Q(n980) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[6]  ( .D(\fpu_add_frac_dp/n3554 ), .CLK(n1532), .Q(n981) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[5]  ( .D(\fpu_add_frac_dp/n3555 ), .CLK(n1532), .Q(n982) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[4]  ( .D(\fpu_add_frac_dp/n3556 ), .CLK(n1532), .Q(n983) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[3]  ( .D(\fpu_add_frac_dp/n3557 ), .CLK(n1535), .Q(n984) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[2]  ( .D(\fpu_add_frac_dp/n3558 ), .CLK(n1535), .Q(n985) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[1]  ( .D(\fpu_add_frac_dp/n3559 ), .CLK(n1536), .Q(n986) );
  DFFX1 \fpu_add_frac_dp/i_a5stg_rndadd/q_reg[0]  ( .D(\fpu_add_frac_dp/n3560 ), .CLK(n1536), .Q(n987) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[63]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N66 ), .CLK(n1529), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[63] ), .QN(\fpu_add_frac_dp/n187 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[63]  ( .D(
        \fpu_add_frac_dp/n3561 ), .CLK(n1551), .Q(n846), .QN(
        \fpu_add_frac_dp/n188 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[62]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N65 ), .CLK(n1529), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[62] ), .QN(\fpu_add_frac_dp/n189 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[62]  ( .D(
        \fpu_add_frac_dp/n3562 ), .CLK(n1551), .Q(n831), .QN(
        \fpu_add_frac_dp/n190 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[61]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N64 ), .CLK(n1530), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[61] ), .QN(\fpu_add_frac_dp/n191 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[61]  ( .D(
        \fpu_add_frac_dp/n3563 ), .CLK(n1551), .Q(n832), .QN(
        \fpu_add_frac_dp/n192 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[60]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N63 ), .CLK(n1528), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[60] ), .QN(\fpu_add_frac_dp/n193 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[60]  ( .D(
        \fpu_add_frac_dp/n3564 ), .CLK(n1550), .Q(n843), .QN(
        \fpu_add_frac_dp/n194 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[59]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N62 ), .CLK(n1529), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[59] ), .QN(\fpu_add_frac_dp/n195 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[59]  ( .D(
        \fpu_add_frac_dp/n3565 ), .CLK(n1550), .Q(n840), .QN(
        \fpu_add_frac_dp/n196 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[58]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N61 ), .CLK(n1529), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[58] ), .QN(\fpu_add_frac_dp/n197 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[58]  ( .D(
        \fpu_add_frac_dp/n3566 ), .CLK(n1550), .Q(n833), .QN(
        \fpu_add_frac_dp/n198 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[57]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N60 ), .CLK(n1530), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[57] ), .QN(\fpu_add_frac_dp/n199 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[57]  ( .D(
        \fpu_add_frac_dp/n3567 ), .CLK(n1550), .Q(n834), .QN(
        \fpu_add_frac_dp/n200 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[56]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N59 ), .CLK(n1530), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[56] ), .QN(\fpu_add_frac_dp/n201 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[56]  ( .D(
        \fpu_add_frac_dp/n3568 ), .CLK(n1550), .Q(n844), .QN(
        \fpu_add_frac_dp/n202 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[55]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N58 ), .CLK(n1536), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[55] ), .QN(\fpu_add_frac_dp/n203 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[55]  ( .D(
        \fpu_add_frac_dp/n3569 ), .CLK(n1550), .Q(n841), .QN(
        \fpu_add_frac_dp/n204 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[54]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N57 ), .CLK(n1537), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[54] ), .QN(\fpu_add_frac_dp/n205 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[54]  ( .D(
        \fpu_add_frac_dp/n3570 ), .CLK(n1550), .Q(n835), .QN(
        \fpu_add_frac_dp/n206 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[53]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N56 ), .CLK(n1531), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[53] ), .QN(\fpu_add_frac_dp/n207 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[53]  ( .D(
        \fpu_add_frac_dp/n3571 ), .CLK(n1550), .Q(n836), .QN(
        \fpu_add_frac_dp/n208 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[52]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N55 ), .CLK(n1531), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[52] ), .QN(\fpu_add_frac_dp/n209 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[52]  ( .D(
        \fpu_add_frac_dp/n3572 ), .CLK(n1550), .Q(n845), .QN(
        \fpu_add_frac_dp/n210 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[51]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N54 ), .CLK(n1531), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[51] ), .QN(\fpu_add_frac_dp/n211 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[51]  ( .D(
        \fpu_add_frac_dp/n3573 ), .CLK(n1550), .Q(n842), .QN(
        \fpu_add_frac_dp/n212 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[50]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N53 ), .CLK(n1531), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[50] ), .QN(\fpu_add_frac_dp/n213 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[50]  ( .D(
        \fpu_add_frac_dp/n3574 ), .CLK(n1550), .Q(n837), .QN(
        \fpu_add_frac_dp/n214 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[49]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N52 ), .CLK(n1526), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[49] ), .QN(\fpu_add_frac_dp/n215 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[49]  ( .D(
        \fpu_add_frac_dp/n3575 ), .CLK(n1550), .Q(n838), .QN(
        \fpu_add_frac_dp/n216 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[48]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N51 ), .CLK(n1525), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[48] ), .QN(\fpu_add_frac_dp/n217 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[48]  ( .D(
        \fpu_add_frac_dp/n3576 ), .CLK(n1550), .Q(n914), .QN(
        \fpu_add_frac_dp/n218 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[47]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N50 ), .CLK(n1525), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[47] ), .QN(\fpu_add_frac_dp/n219 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[47]  ( .D(
        \fpu_add_frac_dp/n3577 ), .CLK(n1550), .Q(n451), .QN(
        \fpu_add_frac_dp/n220 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[46]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N49 ), .CLK(n1525), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[46] ), .QN(\fpu_add_frac_dp/n221 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[46]  ( .D(
        \fpu_add_frac_dp/n3578 ), .CLK(n1549), .Q(n456), .QN(
        \fpu_add_frac_dp/n222 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[45]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N48 ), .CLK(n1525), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[45] ), .QN(\fpu_add_frac_dp/n223 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[45]  ( .D(
        \fpu_add_frac_dp/n3579 ), .CLK(n1549), .Q(n457), .QN(
        \fpu_add_frac_dp/n224 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[44]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N47 ), .CLK(n1525), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[44] ), .QN(\fpu_add_frac_dp/n225 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[44]  ( .D(
        \fpu_add_frac_dp/n3580 ), .CLK(n1549), .Q(n464), .QN(
        \fpu_add_frac_dp/n226 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[43]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N46 ), .CLK(n1524), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[43] ), .QN(\fpu_add_frac_dp/n227 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[43]  ( .D(
        \fpu_add_frac_dp/n3581 ), .CLK(n1549), .Q(n461), .QN(
        \fpu_add_frac_dp/n228 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[42]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N45 ), .CLK(n1524), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[42] ), .QN(\fpu_add_frac_dp/n229 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[42]  ( .D(
        \fpu_add_frac_dp/n3582 ), .CLK(n1549), .Q(n766), .QN(
        \fpu_add_frac_dp/n230 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[41]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N44 ), .CLK(n1524), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[41] ), .QN(\fpu_add_frac_dp/n231 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[41]  ( .D(
        \fpu_add_frac_dp/n3583 ), .CLK(n1549), .Q(n462), .QN(
        \fpu_add_frac_dp/n232 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[40]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N43 ), .CLK(n1524), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[40] ), .QN(\fpu_add_frac_dp/n233 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[40]  ( .D(
        \fpu_add_frac_dp/n3584 ), .CLK(n1549), .Q(n458), .QN(
        \fpu_add_frac_dp/n234 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[39]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N42 ), .CLK(n1524), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[39] ), .QN(\fpu_add_frac_dp/n235 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[39]  ( .D(
        \fpu_add_frac_dp/n3585 ), .CLK(n1549), .Q(n459), .QN(
        \fpu_add_frac_dp/n236 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[38]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N41 ), .CLK(n1523), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[38] ), .QN(\fpu_add_frac_dp/n237 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[38]  ( .D(
        \fpu_add_frac_dp/n3586 ), .CLK(n1549), .Q(n767), .QN(
        \fpu_add_frac_dp/n238 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[37]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N40 ), .CLK(n1523), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[37] ), .QN(\fpu_add_frac_dp/n239 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[37]  ( .D(
        \fpu_add_frac_dp/n3587 ), .CLK(n1549), .Q(n765), .QN(
        \fpu_add_frac_dp/n240 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[36]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N39 ), .CLK(n1523), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[36] ), .QN(\fpu_add_frac_dp/n241 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[36]  ( .D(
        \fpu_add_frac_dp/n3588 ), .CLK(n1549), .Q(n742), .QN(
        \fpu_add_frac_dp/n242 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[35]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N38 ), .CLK(n1523), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[35] ), .QN(\fpu_add_frac_dp/n243 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[35]  ( .D(
        \fpu_add_frac_dp/n3589 ), .CLK(n1549), .Q(n741), .QN(
        \fpu_add_frac_dp/n244 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[34]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N37 ), .CLK(n1522), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[34] ), .QN(\fpu_add_frac_dp/n245 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[34]  ( .D(
        \fpu_add_frac_dp/n3590 ), .CLK(n1549), .Q(n739), .QN(
        \fpu_add_frac_dp/n246 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[33]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N36 ), .CLK(n1522), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[33] ), .QN(\fpu_add_frac_dp/n247 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[33]  ( .D(
        \fpu_add_frac_dp/n3591 ), .CLK(n1549), .Q(n740), .QN(
        \fpu_add_frac_dp/n248 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[32]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N35 ), .CLK(n1521), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[32] ), .QN(\fpu_add_frac_dp/n249 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[32]  ( .D(
        \fpu_add_frac_dp/n3592 ), .CLK(n1548), .Q(n1090), .QN(
        \fpu_add_frac_dp/n250 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[31]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N34 ), .CLK(n1521), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[31] ), .QN(\fpu_add_frac_dp/n251 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[31]  ( .D(
        \fpu_add_frac_dp/n3593 ), .CLK(n1548), .Q(n729), .QN(
        \fpu_add_frac_dp/n252 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[30]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N33 ), .CLK(n1521), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[30] ), .QN(\fpu_add_frac_dp/n253 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[30]  ( .D(
        \fpu_add_frac_dp/n3594 ), .CLK(n1548), .Q(n726), .QN(
        \fpu_add_frac_dp/n254 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[29]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N32 ), .CLK(n1521), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[29] ), .QN(\fpu_add_frac_dp/n255 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[29]  ( .D(
        \fpu_add_frac_dp/n3595 ), .CLK(n1548), .Q(n727), .QN(
        \fpu_add_frac_dp/n256 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[28]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N31 ), .CLK(n1520), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[28] ), .QN(\fpu_add_frac_dp/n257 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[28]  ( .D(
        \fpu_add_frac_dp/n3596 ), .CLK(n1548), .Q(n751), .QN(
        \fpu_add_frac_dp/n258 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[27]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N30 ), .CLK(n1520), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[27] ), .QN(\fpu_add_frac_dp/n259 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[27]  ( .D(
        \fpu_add_frac_dp/n3597 ), .CLK(n1548), .Q(n749), .QN(
        \fpu_add_frac_dp/n260 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[26]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N29 ), .CLK(n1520), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[26] ), .QN(\fpu_add_frac_dp/n261 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[26]  ( .D(
        \fpu_add_frac_dp/n3598 ), .CLK(n1548), .Q(n448), .QN(
        \fpu_add_frac_dp/n262 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[25]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N28 ), .CLK(n1520), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[25] ), .QN(\fpu_add_frac_dp/n263 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[25]  ( .D(
        \fpu_add_frac_dp/n3599 ), .CLK(n1548), .Q(n748), .QN(
        \fpu_add_frac_dp/n264 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[24]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N27 ), .CLK(n1537), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[24] ), .QN(\fpu_add_frac_dp/n265 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[24]  ( .D(
        \fpu_add_frac_dp/n3600 ), .CLK(n1548), .Q(n752), .QN(
        \fpu_add_frac_dp/n266 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[23]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N26 ), .CLK(n1538), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[23] ), .QN(\fpu_add_frac_dp/n267 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[23]  ( .D(
        \fpu_add_frac_dp/n3601 ), .CLK(n1548), .Q(n750), .QN(
        \fpu_add_frac_dp/n268 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[22]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N25 ), .CLK(n1518), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[22] ), .QN(\fpu_add_frac_dp/n269 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[22]  ( .D(
        \fpu_add_frac_dp/n3602 ), .CLK(n1548), .Q(n449), .QN(
        \fpu_add_frac_dp/n270 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[21]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N24 ), .CLK(n1519), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[21] ), .QN(\fpu_add_frac_dp/n271 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[21]  ( .D(
        \fpu_add_frac_dp/n3603 ), .CLK(n1548), .Q(n450), .QN(
        \fpu_add_frac_dp/n272 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[20]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N23 ), .CLK(n1519), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[20] ), .QN(\fpu_add_frac_dp/n273 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[20]  ( .D(
        \fpu_add_frac_dp/n3604 ), .CLK(n1552), .Q(n432), .QN(
        \fpu_add_frac_dp/n274 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[19]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N22 ), .CLK(n1519), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[19] ), .QN(\fpu_add_frac_dp/n275 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[19]  ( .D(
        \fpu_add_frac_dp/n3605 ), .CLK(n1528), .Q(n431), .QN(
        \fpu_add_frac_dp/n276 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[18]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N21 ), .CLK(n1519), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[18] ), .QN(\fpu_add_frac_dp/n277 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[18]  ( .D(
        \fpu_add_frac_dp/n3606 ), .CLK(n1528), .Q(n429), .QN(
        \fpu_add_frac_dp/n278 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[17]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N20 ), .CLK(n1537), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[17] ), .QN(\fpu_add_frac_dp/n279 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[17]  ( .D(
        \fpu_add_frac_dp/n3607 ), .CLK(n1528), .Q(n430), .QN(
        \fpu_add_frac_dp/n280 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[16]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N19 ), .CLK(n1537), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[16] ), .QN(\fpu_add_frac_dp/n281 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[16]  ( .D(
        \fpu_add_frac_dp/n3608 ), .CLK(n1528), .Q(n756), .QN(
        \fpu_add_frac_dp/n282 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[15]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N18 ), .CLK(n1534), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[15] ), .QN(\fpu_add_frac_dp/n283 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[15]  ( .D(
        \fpu_add_frac_dp/n3609 ), .CLK(n1528), .Q(n130), .QN(
        \fpu_add_frac_dp/n2417 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[14]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N17 ), .CLK(n1535), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[14] ), .QN(\fpu_add_frac_dp/n285 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[14]  ( .D(
        \fpu_add_frac_dp/n3610 ), .CLK(n1528), .Q(n45), .QN(
        \fpu_add_frac_dp/n2291 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[13]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N16 ), .CLK(n1535), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[13] ), .QN(\fpu_add_frac_dp/n287 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[13]  ( .D(
        \fpu_add_frac_dp/n3611 ), .CLK(n1528), .Q(n257), .QN(
        \fpu_add_frac_dp/n2358 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[12]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N15 ), .CLK(n1536), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[12] ), .QN(\fpu_add_frac_dp/n289 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[12]  ( .D(
        \fpu_add_frac_dp/n3612 ), .CLK(n1528), .Q(n107), .QN(
        \fpu_add_frac_dp/n2292 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[11]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N14 ), .CLK(n1536), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[11] ), .QN(\fpu_add_frac_dp/n291 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[11]  ( .D(
        \fpu_add_frac_dp/n3613 ), .CLK(n1527), .Q(n264), .QN(
        \fpu_add_frac_dp/n2360 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[10]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N13 ), .CLK(n1519), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[10] ), .QN(\fpu_add_frac_dp/n293 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[10]  ( .D(
        \fpu_add_frac_dp/n3614 ), .CLK(n1527), .Q(n119), .QN(
        \fpu_add_frac_dp/n2293 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[9]  ( .D(
        \fpu_add_frac_dp/n1566 ), .RSTB(\fpu_add_frac_dp/n1509 ), .SETB(
        \fpu_add_frac_dp/n1005 ), .CLK(n1476), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[9] ), .QN(\fpu_add_frac_dp/n295 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[9]  ( .D(
        \fpu_add_frac_dp/n3615 ), .CLK(n1527), .Q(n285), .QN(
        \fpu_add_frac_dp/n2410 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[8]  ( .D(
        \fpu_add_frac_dp/n1567 ), .RSTB(\fpu_add_frac_dp/n1509 ), .SETB(
        \fpu_add_frac_dp/n1006 ), .CLK(n1476), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[8] ), .QN(\fpu_add_frac_dp/n297 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[8]  ( .D(
        \fpu_add_frac_dp/n3616 ), .CLK(n1527), .Q(n123), .QN(
        \fpu_add_frac_dp/n2346 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[7]  ( .D(
        \fpu_add_frac_dp/n1568 ), .RSTB(\fpu_add_frac_dp/n1509 ), .SETB(
        \fpu_add_frac_dp/n1007 ), .CLK(n1478), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[7] ), .QN(\fpu_add_frac_dp/n299 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[7]  ( .D(
        \fpu_add_frac_dp/n3617 ), .CLK(n1527), .Q(n286), .QN(
        \fpu_add_frac_dp/n2413 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[6]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N9 ), .CLK(n1535), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[6] ), .QN(\fpu_add_frac_dp/n301 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[6]  ( .D(
        \fpu_add_frac_dp/n3618 ), .CLK(n1527), .Q(n124), .QN(
        \fpu_add_frac_dp/n2349 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[5]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N8 ), .CLK(n1535), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[5] ), .QN(\fpu_add_frac_dp/n303 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[5]  ( .D(
        \fpu_add_frac_dp/n3619 ), .CLK(n1527), .Q(n51), .QN(
        \fpu_add_frac_dp/n2294 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[4]  ( .D(
        \fpu_add_frac_dp/n1571 ), .RSTB(\fpu_add_frac_dp/n1509 ), .SETB(
        \fpu_add_frac_dp/n1001 ), .CLK(n1478), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[4] ), .QN(\fpu_add_frac_dp/n305 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[4]  ( .D(
        \fpu_add_frac_dp/n3620 ), .CLK(n1527), .Q(n284), .QN(
        \fpu_add_frac_dp/n2414 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[3]  ( .D(
        \fpu_add_frac_dp/n1572 ), .RSTB(\fpu_add_frac_dp/n1509 ), .SETB(
        \fpu_add_frac_dp/n1002 ), .CLK(n1477), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[3] ), .QN(\fpu_add_frac_dp/n307 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[3]  ( .D(
        \fpu_add_frac_dp/n3621 ), .CLK(n1527), .Q(n50), .QN(
        \fpu_add_frac_dp/n2347 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[2]  ( .D(
        \fpu_add_frac_dp/n1573 ), .RSTB(\fpu_add_frac_dp/n1509 ), .SETB(
        \fpu_add_frac_dp/n1003 ), .CLK(n1477), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[2] ), .QN(\fpu_add_frac_dp/n309 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[2]  ( .D(
        \fpu_add_frac_dp/n3622 ), .CLK(n1527), .Q(n115), .QN(
        \fpu_add_frac_dp/n2412 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[1]  ( .D(
        \fpu_add_frac_dp/n1574 ), .RSTB(\fpu_add_frac_dp/n1509 ), .SETB(
        \fpu_add_frac_dp/n1004 ), .CLK(n1477), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre2[1] ), .QN(\fpu_add_frac_dp/n311 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[1]  ( .D(
        \fpu_add_frac_dp/n3623 ), .CLK(n1527), .Q(n48), .QN(
        \fpu_add_frac_dp/n2348 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/q_reg[0]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N3 ), .CLK(n1522), .Q(n956), 
        .QN(\fpu_add_frac_dp/n313 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_shl_data/q_reg[0]  ( .D(
        \fpu_add_frac_dp/n3624 ), .CLK(n1527), .Q(n219), .QN(
        \fpu_add_frac_dp/n2401 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[63]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N66 ), .CLK(n1541), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[63] ), .QN(\fpu_add_frac_dp/n315 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[62]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N65 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[62] ), .QN(\fpu_add_frac_dp/n316 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[61]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N64 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[61] ), .QN(\fpu_add_frac_dp/n317 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[60]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N63 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[60] ), .QN(\fpu_add_frac_dp/n318 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[59]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N62 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[59] ), .QN(\fpu_add_frac_dp/n319 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[58]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N61 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[58] ), .QN(\fpu_add_frac_dp/n320 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[57]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N60 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[57] ), .QN(\fpu_add_frac_dp/n321 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[56]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N59 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[56] ), .QN(\fpu_add_frac_dp/n322 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[55]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N58 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[55] ), .QN(\fpu_add_frac_dp/n323 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[54]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N57 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[54] ), .QN(\fpu_add_frac_dp/n324 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[53]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N56 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[53] ), .QN(\fpu_add_frac_dp/n325 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[52]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N55 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[52] ), .QN(\fpu_add_frac_dp/n326 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[51]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N54 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[51] ), .QN(\fpu_add_frac_dp/n327 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[50]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N53 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[50] ), .QN(\fpu_add_frac_dp/n328 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[49]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N52 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[49] ), .QN(\fpu_add_frac_dp/n329 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[48]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N51 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[48] ), .QN(\fpu_add_frac_dp/n330 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[47]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N50 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[47] ), .QN(\fpu_add_frac_dp/n331 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[46]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N49 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[46] ), .QN(\fpu_add_frac_dp/n332 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[45]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N48 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[45] ), .QN(\fpu_add_frac_dp/n333 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[44]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N47 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[44] ), .QN(\fpu_add_frac_dp/n334 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[43]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N46 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[43] ), .QN(\fpu_add_frac_dp/n335 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[42]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N45 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[42] ), .QN(\fpu_add_frac_dp/n336 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[41]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N44 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[41] ), .QN(\fpu_add_frac_dp/n337 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[40]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N43 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[40] ), .QN(\fpu_add_frac_dp/n338 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[39]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N42 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[39] ), .QN(\fpu_add_frac_dp/n339 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[38]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N41 ), .CLK(n1539), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[38] ), .QN(\fpu_add_frac_dp/n340 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[37]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N40 ), .CLK(n1538), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[37] ), .QN(\fpu_add_frac_dp/n341 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[36]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N39 ), .CLK(n1538), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[36] ), .QN(\fpu_add_frac_dp/n342 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[35]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N38 ), .CLK(n1538), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[35] ), .QN(\fpu_add_frac_dp/n343 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[34]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N37 ), .CLK(n1538), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[34] ), .QN(\fpu_add_frac_dp/n344 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[33]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N36 ), .CLK(n1538), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[33] ), .QN(\fpu_add_frac_dp/n345 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[32]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N35 ), .CLK(n1538), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[32] ), .QN(\fpu_add_frac_dp/n346 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[31]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N34 ), .CLK(n1538), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[31] ), .QN(\fpu_add_frac_dp/n347 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[30]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N33 ), .CLK(n1538), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[30] ), .QN(\fpu_add_frac_dp/n348 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[29]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N32 ), .CLK(n1538), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[29] ), .QN(\fpu_add_frac_dp/n349 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[28]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N31 ), .CLK(n1543), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[28] ), .QN(\fpu_add_frac_dp/n350 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[27]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N30 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[27] ), .QN(\fpu_add_frac_dp/n351 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[26]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N29 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[26] ), .QN(\fpu_add_frac_dp/n352 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[25]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N28 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[25] ), .QN(\fpu_add_frac_dp/n353 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[24]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N27 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[24] ), .QN(\fpu_add_frac_dp/n354 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[23]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N26 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[23] ), .QN(\fpu_add_frac_dp/n355 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[22]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N25 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[22] ), .QN(\fpu_add_frac_dp/n356 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[21]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N24 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[21] ), .QN(\fpu_add_frac_dp/n357 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[20]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N23 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[20] ), .QN(\fpu_add_frac_dp/n358 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[19]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N22 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[19] ), .QN(\fpu_add_frac_dp/n359 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[18]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N21 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[18] ), .QN(\fpu_add_frac_dp/n360 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[17]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N20 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[17] ), .QN(\fpu_add_frac_dp/n361 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[16]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N19 ), .CLK(n1557), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[16] ), .QN(\fpu_add_frac_dp/n362 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[15]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N18 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[15] ), .QN(\fpu_add_frac_dp/n363 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[14]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N17 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[14] ), .QN(\fpu_add_frac_dp/n364 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[13]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N16 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[13] ), .QN(\fpu_add_frac_dp/n365 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[12]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N15 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[12] ), .QN(\fpu_add_frac_dp/n366 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[11]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N14 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[11] ), .QN(\fpu_add_frac_dp/n367 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[10]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N13 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[10] ), .QN(\fpu_add_frac_dp/n368 ) );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[9]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N12 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[9] ), .QN(\fpu_add_frac_dp/n369 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[8]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N11 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[8] ), .QN(\fpu_add_frac_dp/n370 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[7]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N10 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[7] ), .QN(\fpu_add_frac_dp/n371 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[6]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N9 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[6] ), .QN(\fpu_add_frac_dp/n372 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[5]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N8 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[5] ), .QN(\fpu_add_frac_dp/n373 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[4]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N7 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[4] ), .QN(\fpu_add_frac_dp/n374 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[3]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N6 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[3] ), .QN(\fpu_add_frac_dp/n375 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[2]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N5 ), .CLK(n1556), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[2] ), .QN(\fpu_add_frac_dp/n376 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/q_reg[1]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N4 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre3[1] ), .QN(\fpu_add_frac_dp/n377 )
         );
  DFFX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[63]  ( .D(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .CLK(n1540), .Q(
        \fpu_add_frac_dp/a4stg_rnd_frac_pre1[63] ), .QN(\fpu_add_frac_dp/n378 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[62]  ( .D(
        \fpu_add_frac_dp/n1515 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1479), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[62] ), .QN(
        \fpu_add_frac_dp/n380 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[61]  ( .D(
        \fpu_add_frac_dp/n1516 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1479), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[61] ), .QN(
        \fpu_add_frac_dp/n382 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[60]  ( .D(
        \fpu_add_frac_dp/n1517 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1478), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[60] ), .QN(
        \fpu_add_frac_dp/n384 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[59]  ( .D(
        \fpu_add_frac_dp/n1518 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1478), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[59] ), .QN(
        \fpu_add_frac_dp/n386 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[58]  ( .D(
        \fpu_add_frac_dp/n1519 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1478), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[58] ), .QN(
        \fpu_add_frac_dp/n388 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[57]  ( .D(
        \fpu_add_frac_dp/n1520 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1478), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[57] ), .QN(
        \fpu_add_frac_dp/n390 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[56]  ( .D(
        \fpu_add_frac_dp/n1521 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1477), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[56] ), .QN(
        \fpu_add_frac_dp/n392 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[55]  ( .D(
        \fpu_add_frac_dp/n1522 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1477), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[55] ), .QN(
        \fpu_add_frac_dp/n394 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[54]  ( .D(
        \fpu_add_frac_dp/n1523 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1477), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[54] ), .QN(
        \fpu_add_frac_dp/n396 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[53]  ( .D(
        \fpu_add_frac_dp/n1524 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1477), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[53] ), .QN(
        \fpu_add_frac_dp/n398 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[52]  ( .D(
        \fpu_add_frac_dp/n1525 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1476), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[52] ), .QN(
        \fpu_add_frac_dp/n400 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[51]  ( .D(
        \fpu_add_frac_dp/n1526 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1476), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[51] ), .QN(
        \fpu_add_frac_dp/n402 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[50]  ( .D(
        \fpu_add_frac_dp/n1527 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1477), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[50] ), .QN(
        \fpu_add_frac_dp/n404 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[49]  ( .D(
        \fpu_add_frac_dp/n1528 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1477), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[49] ), .QN(
        \fpu_add_frac_dp/n406 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[48]  ( .D(
        \fpu_add_frac_dp/n1529 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1476), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[48] ), .QN(
        \fpu_add_frac_dp/n408 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[47]  ( .D(
        \fpu_add_frac_dp/n1530 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1476), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[47] ), .QN(
        \fpu_add_frac_dp/n410 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[46]  ( .D(
        \fpu_add_frac_dp/n1531 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1476), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[46] ), .QN(
        \fpu_add_frac_dp/n412 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[45]  ( .D(
        \fpu_add_frac_dp/n1532 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1476), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[45] ), .QN(
        \fpu_add_frac_dp/n414 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[44]  ( .D(
        \fpu_add_frac_dp/n1533 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[44] ), .QN(
        \fpu_add_frac_dp/n416 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[43]  ( .D(
        \fpu_add_frac_dp/n1534 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1476), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[43] ), .QN(
        \fpu_add_frac_dp/n418 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[42]  ( .D(
        \fpu_add_frac_dp/n1535 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[42] ), .QN(
        \fpu_add_frac_dp/n420 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[41]  ( .D(
        \fpu_add_frac_dp/n1536 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[41] ), .QN(
        \fpu_add_frac_dp/n422 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[40]  ( .D(
        \fpu_add_frac_dp/n1537 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[40] ), .QN(
        \fpu_add_frac_dp/n424 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[39]  ( .D(
        \fpu_add_frac_dp/n1538 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[39] ), .QN(
        \fpu_add_frac_dp/n426 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[38]  ( .D(
        \fpu_add_frac_dp/n1539 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[38] ), .QN(
        \fpu_add_frac_dp/n428 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[37]  ( .D(
        \fpu_add_frac_dp/n1540 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[37] ), .QN(
        \fpu_add_frac_dp/n430 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[36]  ( .D(
        \fpu_add_frac_dp/n1541 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[36] ), .QN(
        \fpu_add_frac_dp/n432 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[35]  ( .D(
        \fpu_add_frac_dp/n1542 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[35] ), .QN(
        \fpu_add_frac_dp/n434 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[34]  ( .D(
        \fpu_add_frac_dp/n1543 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[34] ), .QN(
        \fpu_add_frac_dp/n436 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[33]  ( .D(
        \fpu_add_frac_dp/n1544 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[33] ), .QN(
        \fpu_add_frac_dp/n438 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[32]  ( .D(
        \fpu_add_frac_dp/n1545 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[32] ), .QN(
        \fpu_add_frac_dp/n440 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[31]  ( .D(
        \fpu_add_frac_dp/n1546 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[31] ), .QN(
        \fpu_add_frac_dp/n442 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[30]  ( .D(
        \fpu_add_frac_dp/n1547 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[30] ), .QN(
        \fpu_add_frac_dp/n444 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[29]  ( .D(
        \fpu_add_frac_dp/n1548 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[29] ), .QN(
        \fpu_add_frac_dp/n446 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[28]  ( .D(
        \fpu_add_frac_dp/n1549 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[28] ), .QN(
        \fpu_add_frac_dp/n448 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[27]  ( .D(
        \fpu_add_frac_dp/n1550 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[27] ), .QN(
        \fpu_add_frac_dp/n450 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[26]  ( .D(
        \fpu_add_frac_dp/n1551 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[26] ), .QN(
        \fpu_add_frac_dp/n452 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[25]  ( .D(
        \fpu_add_frac_dp/n1552 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[25] ), .QN(
        \fpu_add_frac_dp/n454 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[24]  ( .D(
        \fpu_add_frac_dp/n1553 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1474), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[24] ), .QN(
        \fpu_add_frac_dp/n456 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[23]  ( .D(
        \fpu_add_frac_dp/n1554 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[23] ), .QN(
        \fpu_add_frac_dp/n458 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[22]  ( .D(
        \fpu_add_frac_dp/n1555 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[22] ), .QN(
        \fpu_add_frac_dp/n460 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[21]  ( .D(
        \fpu_add_frac_dp/n1556 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[21] ), .QN(
        \fpu_add_frac_dp/n462 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[20]  ( .D(
        \fpu_add_frac_dp/n1557 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1475), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[20] ), .QN(
        \fpu_add_frac_dp/n464 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[19]  ( .D(
        \fpu_add_frac_dp/n1558 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1476), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[19] ), .QN(
        \fpu_add_frac_dp/n466 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[18]  ( .D(
        \fpu_add_frac_dp/n1559 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1476), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[18] ), .QN(
        \fpu_add_frac_dp/n468 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[17]  ( .D(
        \fpu_add_frac_dp/n1560 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1477), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[17] ), .QN(
        \fpu_add_frac_dp/n470 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[16]  ( .D(
        \fpu_add_frac_dp/n1561 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1478), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[16] ), .QN(
        \fpu_add_frac_dp/n472 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[15]  ( .D(
        \fpu_add_frac_dp/n1562 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1477), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[15] ), .QN(
        \fpu_add_frac_dp/n474 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[14]  ( .D(
        \fpu_add_frac_dp/n1563 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1478), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[14] ), .QN(
        \fpu_add_frac_dp/n476 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[13]  ( .D(
        \fpu_add_frac_dp/n1564 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1476), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[13] ), .QN(
        \fpu_add_frac_dp/n478 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[12]  ( .D(
        \fpu_add_frac_dp/n1565 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1478), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[12] ), .QN(
        \fpu_add_frac_dp/n480 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[11]  ( .D(
        \fpu_add_frac_dp/n1566 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1479), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[11] ), .QN(
        \fpu_add_frac_dp/n482 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[10]  ( .D(
        \fpu_add_frac_dp/n1567 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1478), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[10] ), .QN(
        \fpu_add_frac_dp/n484 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[9]  ( .D(
        \fpu_add_frac_dp/n1568 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1478), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[9] ), .QN(
        \fpu_add_frac_dp/n486 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[8]  ( .D(
        \fpu_add_frac_dp/n1569 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1479), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[8] ), .QN(
        \fpu_add_frac_dp/n488 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[7]  ( .D(
        \fpu_add_frac_dp/n1570 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1479), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[7] ), .QN(
        \fpu_add_frac_dp/n490 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[6]  ( .D(
        \fpu_add_frac_dp/n1571 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1477), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[6] ), .QN(
        \fpu_add_frac_dp/n492 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[5]  ( .D(
        \fpu_add_frac_dp/n1572 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1479), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[5] ), .QN(
        \fpu_add_frac_dp/n494 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[4]  ( .D(
        \fpu_add_frac_dp/n1573 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1479), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[4] ), .QN(
        \fpu_add_frac_dp/n496 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[3]  ( .D(
        \fpu_add_frac_dp/n1574 ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1479), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[3] ), .QN(
        \fpu_add_frac_dp/n498 ) );
  DFFSSRX1 \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/q_reg[2]  ( .D(
        \fpu_add_frac_dp/a3stg_fracadd[0] ), .RSTB(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ), .SETB(1'b1), .CLK(n1478), 
        .Q(\fpu_add_frac_dp/a4stg_rnd_frac_pre1[2] ), .QN(
        \fpu_add_frac_dp/n500 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[7]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N10 ), .CLK(n1545), .Q(n413), .QN(
        \fpu_add_frac_dp/n501 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[8]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N11 ), .CLK(n1545), .Q(n412), .QN(
        \fpu_add_frac_dp/n502 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[1]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N4 ), .CLK(n1543), .Q(n419), .QN(
        \fpu_add_frac_dp/n503 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[2]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N5 ), .CLK(n1542), .Q(n418), .QN(
        \fpu_add_frac_dp/n504 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[3]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N6 ), .CLK(n1541), .Q(n417), .QN(
        \fpu_add_frac_dp/n505 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[4]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N7 ), .CLK(n1541), .Q(n416), .QN(
        \fpu_add_frac_dp/n506 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[6]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N9 ), .CLK(n1541), .Q(n414), .QN(
        \fpu_add_frac_dp/n507 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[5]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N8 ), .CLK(n1541), .Q(n415), .QN(
        \fpu_add_frac_dp/n508 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[0]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N3 ), .CLK(n1544), .Q(n139), .QN(
        \fpu_add_frac_dp/n509 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[4]  ( .D(
        \fpu_add_frac_dp/n3735 ), .CLK(n1481), .Q(n1264), .QN(
        \fpu_add_frac_dp/n510 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[9]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N12 ), .CLK(n1545), .Q(n411), .QN(
        \fpu_add_frac_dp/n511 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[10]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N13 ), .CLK(n1545), .Q(n410), .QN(
        \fpu_add_frac_dp/n512 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[63]  ( .D(
        \fpu_add_frac_dp/n3738 ), .CLK(n1510), .Q(n1219), .QN(
        \fpu_add_frac_dp/n513 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[11]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N14 ), .CLK(n1545), .Q(n409), .QN(
        \fpu_add_frac_dp/n514 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[5]  ( .D(
        \fpu_add_frac_dp/n3734 ), .CLK(n1481), .Q(n1302), .QN(
        \fpu_add_frac_dp/n515 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[12]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N15 ), .CLK(n1545), .Q(n408), .QN(
        \fpu_add_frac_dp/n516 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[13]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N16 ), .CLK(n1545), .Q(n407), .QN(
        \fpu_add_frac_dp/n517 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[14]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N17 ), .CLK(n1545), .Q(n406), .QN(
        \fpu_add_frac_dp/n518 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[15]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N18 ), .CLK(n1545), .Q(n405), .QN(
        \fpu_add_frac_dp/n519 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[16]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N19 ), .CLK(n1545), .Q(n404), .QN(
        \fpu_add_frac_dp/n520 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[17]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N20 ), .CLK(n1545), .Q(n403), .QN(
        \fpu_add_frac_dp/n521 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[18]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N21 ), .CLK(n1544), .Q(n402), .QN(
        \fpu_add_frac_dp/n522 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[19]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N22 ), .CLK(n1544), .Q(n401), .QN(
        \fpu_add_frac_dp/n523 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[20]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N23 ), .CLK(n1544), .Q(n400), .QN(
        \fpu_add_frac_dp/n524 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[21]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N24 ), .CLK(n1544), .Q(n399), .QN(
        \fpu_add_frac_dp/n525 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[22]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N25 ), .CLK(n1544), .Q(n398), .QN(
        \fpu_add_frac_dp/n526 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[23]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N26 ), .CLK(n1544), .Q(n397), .QN(
        \fpu_add_frac_dp/n527 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[62]  ( .D(
        \fpu_add_frac_dp/n3625 ), .CLK(n1512), .Q(n20), .QN(
        \fpu_add_frac_dp/n528 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[24]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N27 ), .CLK(n1544), .Q(n396), .QN(
        \fpu_add_frac_dp/n529 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[25]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N28 ), .CLK(n1544), .Q(n395), .QN(
        \fpu_add_frac_dp/n530 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[26]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N29 ), .CLK(n1544), .Q(n394), .QN(
        \fpu_add_frac_dp/n531 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[27]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N30 ), .CLK(n1544), .Q(n393), .QN(
        \fpu_add_frac_dp/n532 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[28]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N31 ), .CLK(n1544), .Q(n392), .QN(
        \fpu_add_frac_dp/n533 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[29]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N32 ), .CLK(n1544), .Q(n391), .QN(
        \fpu_add_frac_dp/n534 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[30]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N33 ), .CLK(n1544), .Q(n390), .QN(
        \fpu_add_frac_dp/n535 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[31]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N34 ), .CLK(n1543), .Q(n389), .QN(
        \fpu_add_frac_dp/n536 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[32]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N35 ), .CLK(n1543), .Q(n388), .QN(
        \fpu_add_frac_dp/n537 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[33]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N36 ), .CLK(n1543), .Q(n387), .QN(
        \fpu_add_frac_dp/n538 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[34]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N37 ), .CLK(n1543), .Q(n386), .QN(
        \fpu_add_frac_dp/n539 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[35]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N38 ), .CLK(n1543), .Q(n385), .QN(
        \fpu_add_frac_dp/n540 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[36]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N39 ), .CLK(n1543), .Q(n384), .QN(
        \fpu_add_frac_dp/n541 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[37]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N40 ), .CLK(n1543), .Q(n383), .QN(
        \fpu_add_frac_dp/n542 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[38]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N41 ), .CLK(n1543), .Q(n382), .QN(
        \fpu_add_frac_dp/n543 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[39]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N42 ), .CLK(n1543), .Q(n381), .QN(
        \fpu_add_frac_dp/n544 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[61]  ( .D(
        \fpu_add_frac_dp/n3626 ), .CLK(n1512), .Q(n118), .QN(
        \fpu_add_frac_dp/n545 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[40]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N43 ), .CLK(n1543), .Q(n380), .QN(
        \fpu_add_frac_dp/n546 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[41]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N44 ), .CLK(n1543), .Q(n379), .QN(
        \fpu_add_frac_dp/n547 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[42]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N45 ), .CLK(n1543), .Q(n378), .QN(
        \fpu_add_frac_dp/n548 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[43]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N46 ), .CLK(n1542), .Q(n377), .QN(
        \fpu_add_frac_dp/n549 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[44]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N47 ), .CLK(n1542), .Q(n376), .QN(
        \fpu_add_frac_dp/n550 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[45]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N48 ), .CLK(n1542), .Q(n375), .QN(
        \fpu_add_frac_dp/n551 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[46]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N49 ), .CLK(n1542), .Q(n374), .QN(
        \fpu_add_frac_dp/n552 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[47]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N50 ), .CLK(n1542), .Q(n373), .QN(
        \fpu_add_frac_dp/n553 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[48]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N51 ), .CLK(n1542), .Q(n372), .QN(
        \fpu_add_frac_dp/n554 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[49]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N52 ), .CLK(n1542), .Q(n371), .QN(
        \fpu_add_frac_dp/n555 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[50]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N53 ), .CLK(n1542), .Q(n370), .QN(
        \fpu_add_frac_dp/n556 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[51]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N54 ), .CLK(n1542), .Q(n369), .QN(
        \fpu_add_frac_dp/n557 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[52]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N55 ), .CLK(n1542), .Q(n368), .QN(
        \fpu_add_frac_dp/n558 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[53]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N56 ), .CLK(n1542), .Q(n367), .QN(
        \fpu_add_frac_dp/n559 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[54]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N57 ), .CLK(n1542), .Q(n366), .QN(
        \fpu_add_frac_dp/n560 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[55]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N58 ), .CLK(n1542), .Q(n365), .QN(
        \fpu_add_frac_dp/n561 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[56]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N59 ), .CLK(n1541), .Q(n364), .QN(
        \fpu_add_frac_dp/n562 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[57]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N60 ), .CLK(n1541), .Q(n363), .QN(
        \fpu_add_frac_dp/n563 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[58]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N61 ), .CLK(n1541), .Q(n362), .QN(
        \fpu_add_frac_dp/n564 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[59]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N62 ), .CLK(n1541), .Q(n361), .QN(
        \fpu_add_frac_dp/n565 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[60]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N63 ), .CLK(n1541), .Q(n360), .QN(
        \fpu_add_frac_dp/n566 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[61]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N64 ), .CLK(n1541), .Q(n359), .QN(
        \fpu_add_frac_dp/n567 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[62]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N65 ), .CLK(n1541), .Q(n753), .QN(
        \fpu_add_frac_dp/n568 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac2/q_reg[63]  ( .D(
        \fpu_add_frac_dp/i_a3stg_frac2/N66 ), .CLK(n1541), .Q(
        \fpu_add_frac_dp/a3stg_frac2[63] ), .QN(\fpu_add_frac_dp/n569 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[60]  ( .D(
        \fpu_add_frac_dp/n3627 ), .CLK(n1512), .Q(n1124), .QN(
        \fpu_add_frac_dp/n570 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[59]  ( .D(
        \fpu_add_frac_dp/n3628 ), .CLK(n1512), .Q(n1222), .QN(
        \fpu_add_frac_dp/n571 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[58]  ( .D(
        \fpu_add_frac_dp/n3629 ), .CLK(n1512), .Q(n5), .QN(
        \fpu_add_frac_dp/n572 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[57]  ( .D(
        \fpu_add_frac_dp/n3630 ), .CLK(n1512), .Q(n47), .QN(
        \fpu_add_frac_dp/n573 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[52]  ( .D(
        \fpu_add_frac_dp/n3631 ), .CLK(n1512), .Q(\fpu_add_frac_dp/n2382 ), 
        .QN(\fpu_add_frac_dp/n1391 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[51]  ( .D(
        \fpu_add_frac_dp/n3632 ), .CLK(n1512), .Q(
        \fpu_add_frac_dp/a2stg_shr_cnt_4[3] ), .QN(\fpu_add_frac_dp/n574 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[50]  ( .D(
        \fpu_add_frac_dp/n3633 ), .CLK(n1512), .Q(n1126), .QN(
        \fpu_add_frac_dp/n575 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[49]  ( .D(
        \fpu_add_frac_dp/n3634 ), .CLK(n1511), .Q(n1221), .QN(
        \fpu_add_frac_dp/n576 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[48]  ( .D(
        \fpu_add_frac_dp/n3635 ), .CLK(n1511), .Q(n1220), .QN(
        \fpu_add_frac_dp/n577 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[47]  ( .D(
        \fpu_add_frac_dp/n3636 ), .CLK(n1511), .Q(\fpu_add_frac_dp/n2322 ), 
        .QN(n580) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[46]  ( .D(
        \fpu_add_frac_dp/n3637 ), .CLK(n1511), .Q(\fpu_add_frac_dp/n2397 ), 
        .QN(\fpu_add_frac_dp/n1384 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[45]  ( .D(
        \fpu_add_frac_dp/n3638 ), .CLK(n1511), .Q(n581), .QN(
        \fpu_add_frac_dp/n2375 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[44]  ( .D(
        \fpu_add_frac_dp/n3639 ), .CLK(n1511), .Q(\fpu_add_frac_dp/n2399 ), 
        .QN(\fpu_add_frac_dp/n1382 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[43]  ( .D(
        \fpu_add_frac_dp/n3640 ), .CLK(n1511), .Q(n1063) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[42]  ( .D(
        \fpu_add_frac_dp/n3641 ), .CLK(n1511), .Q(
        \fpu_add_frac_dp/a2stg_shr_cnt[5] ), .QN(\fpu_add_frac_dp/n579 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[41]  ( .D(
        \fpu_add_frac_dp/n3642 ), .CLK(n1511), .Q(\fpu_add_frac_dp/n2306 ), 
        .QN(n624) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[40]  ( .D(
        \fpu_add_frac_dp/n3643 ), .CLK(n1511), .Q(n693), .QN(
        \fpu_add_frac_dp/n2377 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[39]  ( .D(
        \fpu_add_frac_dp/n3644 ), .CLK(n1511), .Q(n755), .QN(
        \fpu_add_frac_dp/n580 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[38]  ( .D(
        \fpu_add_frac_dp/n3645 ), .CLK(n1511), .Q(n255), .QN(
        \fpu_add_frac_dp/n2308 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[37]  ( .D(
        \fpu_add_frac_dp/n3646 ), .CLK(n1511), .Q(n962), .QN(
        \fpu_add_frac_dp/n2448 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[36]  ( .D(
        \fpu_add_frac_dp/n3647 ), .CLK(n1540), .Q(n296), .QN(
        \fpu_add_frac_dp/n582 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[35]  ( .D(
        \fpu_add_frac_dp/n3648 ), .CLK(n1511), .Q(n746), .QN(
        \fpu_add_frac_dp/n583 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[34]  ( .D(
        \fpu_add_frac_dp/n3649 ), .CLK(n1510), .Q(n653), .QN(
        \fpu_add_frac_dp/n2370 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[33]  ( .D(
        \fpu_add_frac_dp/n3650 ), .CLK(n1510), .Q(n311), .QN(
        \fpu_add_frac_dp/n2465 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[32]  ( .D(
        \fpu_add_frac_dp/n3651 ), .CLK(n1510), .Q(n1145), .QN(
        \fpu_add_frac_dp/n584 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[31]  ( .D(
        \fpu_add_frac_dp/n3652 ), .CLK(n1510), .Q(n166), .QN(
        \fpu_add_frac_dp/n5641 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[30]  ( .D(
        \fpu_add_frac_dp/n3653 ), .CLK(n1510), .Q(n641), .QN(
        \fpu_add_frac_dp/n2385 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[29]  ( .D(
        \fpu_add_frac_dp/n3654 ), .CLK(n1527), .Q(n1144), .QN(
        \fpu_add_frac_dp/n586 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[28]  ( .D(
        \fpu_add_frac_dp/n3655 ), .CLK(n1527), .Q(n596), .QN(
        \fpu_add_frac_dp/n2271 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[27]  ( .D(
        \fpu_add_frac_dp/n3656 ), .CLK(n1526), .Q(\fpu_add_frac_dp/n2320 ), 
        .QN(\fpu_add_frac_dp/n5634 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[25]  ( .D(
        \fpu_add_frac_dp/n3657 ), .CLK(n1526), .Q(
        \fpu_add_frac_dp/a4stg_shl_cnt_dec54_1[1] ), .QN(
        \fpu_add_frac_dp/n589 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[24]  ( .D(
        \fpu_add_frac_dp/n3658 ), .CLK(n1526), .Q(n14), .QN(
        \fpu_add_frac_dp/n5633 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[21]  ( .D(
        \fpu_add_frac_dp/n3659 ), .CLK(n1526), .Q(\fpu_add_frac_dp/n2325 ), 
        .QN(\fpu_add_frac_dp/n5635 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[18]  ( .D(
        \fpu_add_frac_dp/n3660 ), .CLK(n1526), .Q(n2), .QN(
        \fpu_add_frac_dp/n592 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[17]  ( .D(
        \fpu_add_frac_dp/n3661 ), .CLK(n1526), .Q(\a4stg_shl_cnt[5] ), .QN(
        \fpu_add_frac_dp/n593 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[16]  ( .D(
        \fpu_add_frac_dp/n3662 ), .CLK(n1526), .Q(n762), .QN(
        \fpu_add_frac_dp/n594 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[15]  ( .D(
        \fpu_add_frac_dp/n3663 ), .CLK(n1526), .Q(n584), .QN(
        \fpu_add_frac_dp/n2307 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[14]  ( .D(
        \fpu_add_frac_dp/n3664 ), .CLK(n1526), .Q(n63), .QN(
        \fpu_add_frac_dp/n2471 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[13]  ( .D(
        \fpu_add_frac_dp/n3665 ), .CLK(n1526), .Q(n582), .QN(
        \fpu_add_frac_dp/n2460 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[12]  ( .D(
        \fpu_add_frac_dp/n3666 ), .CLK(n1526), .Q(n154), .QN(
        \fpu_add_frac_dp/n2449 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[8]  ( .D(
        \fpu_add_frac_dp/n3731 ), .CLK(n1545), .Q(n64), .QN(
        \fpu_add_frac_dp/n5614 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[7]  ( .D(
        \fpu_add_frac_dp/n3732 ), .CLK(n1510), .Q(\fpu_add_frac_dp/n2369 ), 
        .QN(\fpu_add_frac_dp/n2287 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[6]  ( .D(
        \fpu_add_frac_dp/n3733 ), .CLK(n1551), .Q(n1121), .QN(
        \fpu_add_frac_dp/n596 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[2]  ( .D(
        \fpu_add_frac_dp/n3736 ), .CLK(n1510), .Q(n926), .QN(
        \fpu_add_frac_dp/n2478 ) );
  DFFX1 \fpu_add_frac_dp/i_astg_xtra_regs/q_reg[0]  ( .D(
        \fpu_add_frac_dp/n3737 ), .CLK(n1541), .Q(n852), .QN(
        \fpu_add_frac_dp/n598 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[53]  ( .D(
        \fpu_add_frac_dp/n3739 ), .CLK(n1510), .Q(n1235), .QN(
        \fpu_add_frac_dp/n599 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[52]  ( .D(
        \fpu_add_frac_dp/n3740 ), .CLK(n1510), .Q(n1301), .QN(
        \fpu_add_frac_dp/n600 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[51]  ( .D(
        \fpu_add_frac_dp/n3741 ), .CLK(n1510), .Q(n1300), .QN(
        \fpu_add_frac_dp/n601 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[50]  ( .D(
        \fpu_add_frac_dp/n3742 ), .CLK(n1510), .Q(n1263), .QN(
        \fpu_add_frac_dp/n602 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[49]  ( .D(
        \fpu_add_frac_dp/n3743 ), .CLK(n1510), .Q(n1270), .QN(
        \fpu_add_frac_dp/n603 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[48]  ( .D(
        \fpu_add_frac_dp/n3744 ), .CLK(n1510), .Q(n1299), .QN(
        \fpu_add_frac_dp/n604 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[47]  ( .D(
        \fpu_add_frac_dp/n3745 ), .CLK(n1509), .Q(n1298), .QN(
        \fpu_add_frac_dp/n605 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[46]  ( .D(
        \fpu_add_frac_dp/n3746 ), .CLK(n1509), .Q(n1262), .QN(
        \fpu_add_frac_dp/n606 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[45]  ( .D(
        \fpu_add_frac_dp/n3747 ), .CLK(n1509), .Q(n1244), .QN(
        \fpu_add_frac_dp/n607 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[44]  ( .D(
        \fpu_add_frac_dp/n3748 ), .CLK(n1509), .Q(n1297), .QN(
        \fpu_add_frac_dp/n608 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[43]  ( .D(
        \fpu_add_frac_dp/n3749 ), .CLK(n1509), .Q(n1296), .QN(
        \fpu_add_frac_dp/n609 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[42]  ( .D(
        \fpu_add_frac_dp/n3750 ), .CLK(n1509), .Q(n1261), .QN(
        \fpu_add_frac_dp/n610 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[41]  ( .D(
        \fpu_add_frac_dp/n3751 ), .CLK(n1509), .Q(n1224), .QN(
        \fpu_add_frac_dp/n611 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[40]  ( .D(
        \fpu_add_frac_dp/n3752 ), .CLK(n1509), .Q(n1295), .QN(
        \fpu_add_frac_dp/n612 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[39]  ( .D(
        \fpu_add_frac_dp/n3753 ), .CLK(n1509), .Q(n1294), .QN(
        \fpu_add_frac_dp/n613 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[38]  ( .D(
        \fpu_add_frac_dp/n3754 ), .CLK(n1509), .Q(n1260), .QN(
        \fpu_add_frac_dp/n614 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[37]  ( .D(
        \fpu_add_frac_dp/n3755 ), .CLK(n1509), .Q(n1293), .QN(
        \fpu_add_frac_dp/n615 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[36]  ( .D(
        \fpu_add_frac_dp/n3756 ), .CLK(n1509), .Q(n1259), .QN(
        \fpu_add_frac_dp/n616 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[35]  ( .D(
        \fpu_add_frac_dp/n3757 ), .CLK(n1509), .Q(n1292), .QN(
        \fpu_add_frac_dp/n617 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[34]  ( .D(
        \fpu_add_frac_dp/n3758 ), .CLK(n1509), .Q(n1258), .QN(
        \fpu_add_frac_dp/n618 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[33]  ( .D(
        \fpu_add_frac_dp/n3759 ), .CLK(n1508), .Q(n1291), .QN(
        \fpu_add_frac_dp/n619 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[32]  ( .D(
        \fpu_add_frac_dp/n3760 ), .CLK(n1508), .Q(n1290), .QN(
        \fpu_add_frac_dp/n620 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[31]  ( .D(
        \fpu_add_frac_dp/n3761 ), .CLK(n1508), .Q(n1289), .QN(
        \fpu_add_frac_dp/n621 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[30]  ( .D(
        \fpu_add_frac_dp/n3762 ), .CLK(n1508), .Q(n1257), .QN(
        \fpu_add_frac_dp/n622 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[29]  ( .D(
        \fpu_add_frac_dp/n3763 ), .CLK(n1508), .Q(n1288), .QN(
        \fpu_add_frac_dp/n623 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[28]  ( .D(
        \fpu_add_frac_dp/n3764 ), .CLK(n1508), .Q(n1287), .QN(
        \fpu_add_frac_dp/n624 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[27]  ( .D(
        \fpu_add_frac_dp/n3765 ), .CLK(n1508), .Q(n1256), .QN(
        \fpu_add_frac_dp/n625 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[26]  ( .D(
        \fpu_add_frac_dp/n3766 ), .CLK(n1508), .Q(n1286), .QN(
        \fpu_add_frac_dp/n626 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[25]  ( .D(
        \fpu_add_frac_dp/n3767 ), .CLK(n1508), .Q(n1255), .QN(
        \fpu_add_frac_dp/n627 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[24]  ( .D(
        \fpu_add_frac_dp/n3768 ), .CLK(n1508), .Q(n1243), .QN(
        \fpu_add_frac_dp/n628 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[23]  ( .D(
        \fpu_add_frac_dp/n3769 ), .CLK(n1508), .Q(n1285), .QN(
        \fpu_add_frac_dp/n629 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[22]  ( .D(
        \fpu_add_frac_dp/n3770 ), .CLK(n1508), .Q(n1254), .QN(
        \fpu_add_frac_dp/n630 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[21]  ( .D(
        \fpu_add_frac_dp/n3771 ), .CLK(n1508), .Q(n1269), .QN(
        \fpu_add_frac_dp/n631 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[20]  ( .D(
        \fpu_add_frac_dp/n3772 ), .CLK(n1508), .Q(n1268), .QN(
        \fpu_add_frac_dp/n632 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[19]  ( .D(
        \fpu_add_frac_dp/n3773 ), .CLK(n1507), .Q(n1284), .QN(
        \fpu_add_frac_dp/n633 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[18]  ( .D(
        \fpu_add_frac_dp/n3774 ), .CLK(n1513), .Q(n1253), .QN(
        \fpu_add_frac_dp/n634 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[17]  ( .D(
        \fpu_add_frac_dp/n3775 ), .CLK(n1487), .Q(n1267), .QN(
        \fpu_add_frac_dp/n635 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[16]  ( .D(
        \fpu_add_frac_dp/n3776 ), .CLK(n1480), .Q(n1283), .QN(
        \fpu_add_frac_dp/n636 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[15]  ( .D(
        \fpu_add_frac_dp/n3777 ), .CLK(n1487), .Q(n1282), .QN(
        \fpu_add_frac_dp/n637 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[14]  ( .D(
        \fpu_add_frac_dp/n3778 ), .CLK(n1487), .Q(n1252), .QN(
        \fpu_add_frac_dp/n638 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[13]  ( .D(
        \fpu_add_frac_dp/n3779 ), .CLK(n1487), .Q(n1281), .QN(
        \fpu_add_frac_dp/n639 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[12]  ( .D(
        \fpu_add_frac_dp/n3780 ), .CLK(n1487), .Q(n1280), .QN(
        \fpu_add_frac_dp/n640 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[11]  ( .D(
        \fpu_add_frac_dp/n3781 ), .CLK(n1486), .Q(n1279), .QN(
        \fpu_add_frac_dp/n641 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[10]  ( .D(
        \fpu_add_frac_dp/n3782 ), .CLK(n1486), .Q(n1278), .QN(
        \fpu_add_frac_dp/n642 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[9]  ( .D(\fpu_add_frac_dp/n3783 ), .CLK(n1486), .Q(n1247), .QN(\fpu_add_frac_dp/n643 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[8]  ( .D(\fpu_add_frac_dp/n3784 ), .CLK(n1486), .Q(n1266), .QN(\fpu_add_frac_dp/n644 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[7]  ( .D(\fpu_add_frac_dp/n3785 ), .CLK(n1486), .Q(n1277), .QN(\fpu_add_frac_dp/n645 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[6]  ( .D(\fpu_add_frac_dp/n3786 ), .CLK(n1486), .Q(n1251), .QN(\fpu_add_frac_dp/n646 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[5]  ( .D(\fpu_add_frac_dp/n3787 ), .CLK(n1486), .Q(n1273), .QN(\fpu_add_frac_dp/n647 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[4]  ( .D(\fpu_add_frac_dp/n3788 ), .CLK(n1486), .Q(n1276), .QN(\fpu_add_frac_dp/n648 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[3]  ( .D(\fpu_add_frac_dp/n3789 ), .CLK(n1486), .Q(n1275), .QN(\fpu_add_frac_dp/n649 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[2]  ( .D(\fpu_add_frac_dp/n3790 ), .CLK(n1486), .Q(n1250), .QN(\fpu_add_frac_dp/n650 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[1]  ( .D(\fpu_add_frac_dp/n3791 ), .CLK(n1486), .Q(n1081) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_expdec/q_reg[0]  ( .D(\fpu_add_frac_dp/n3792 ), .CLK(n1486), .Q(n1274), .QN(\fpu_add_frac_dp/n652 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[63]  ( .D(
        \fpu_add_frac_dp/n3667 ), .CLK(n1551), .Q(n87), .QN(
        \fpu_add_frac_dp/n2440 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[62]  ( .D(
        \fpu_add_frac_dp/n3668 ), .CLK(n1551), .Q(n266), .QN(
        \fpu_add_frac_dp/n5618 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[61]  ( .D(
        \fpu_add_frac_dp/n3669 ), .CLK(n1551), .Q(n94), .QN(
        \fpu_add_frac_dp/n2288 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[60]  ( .D(
        \fpu_add_frac_dp/n3670 ), .CLK(n1551), .Q(\fpu_add_frac_dp/n2337 ), 
        .QN(n654) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[59]  ( .D(
        \fpu_add_frac_dp/n3671 ), .CLK(n1551), .Q(n82), .QN(
        \fpu_add_frac_dp/n2394 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[58]  ( .D(
        \fpu_add_frac_dp/n3672 ), .CLK(n1551), .Q(n171), .QN(
        \fpu_add_frac_dp/n654 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[57]  ( .D(
        \fpu_add_frac_dp/n3673 ), .CLK(n1551), .Q(\fpu_add_frac_dp/n2343 ), 
        .QN(\fpu_add_frac_dp/n1355 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[56]  ( .D(
        \fpu_add_frac_dp/n3674 ), .CLK(n1551), .Q(\fpu_add_frac_dp/n2407 ), 
        .QN(\fpu_add_frac_dp/n1354 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[55]  ( .D(
        \fpu_add_frac_dp/n3675 ), .CLK(n1551), .Q(\fpu_add_frac_dp/n2338 ), 
        .QN(\fpu_add_frac_dp/n1352 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[54]  ( .D(
        \fpu_add_frac_dp/n3676 ), .CLK(n1551), .Q(n265), .QN(
        \fpu_add_frac_dp/n2290 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[53]  ( .D(
        \fpu_add_frac_dp/n3677 ), .CLK(n1552), .Q(n92), .QN(
        \fpu_add_frac_dp/n2345 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[52]  ( .D(
        \fpu_add_frac_dp/n3678 ), .CLK(n1552), .Q(n313), .QN(
        \fpu_add_frac_dp/n2416 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[51]  ( .D(
        \fpu_add_frac_dp/n3679 ), .CLK(n1552), .Q(n85), .QN(
        \fpu_add_frac_dp/n2378 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[50]  ( .D(
        \fpu_add_frac_dp/n3680 ), .CLK(n1552), .Q(n22), .QN(
        \fpu_add_frac_dp/n5631 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[49]  ( .D(
        \fpu_add_frac_dp/n3681 ), .CLK(n1552), .Q(n175), .QN(
        \fpu_add_frac_dp/n2386 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[48]  ( .D(
        \fpu_add_frac_dp/n3682 ), .CLK(n1552), .Q(n104), .QN(
        \fpu_add_frac_dp/n5630 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[47]  ( .D(
        \fpu_add_frac_dp/n3683 ), .CLK(n1552), .Q(n40), .QN(
        \fpu_add_frac_dp/n2333 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[46]  ( .D(
        \fpu_add_frac_dp/n3684 ), .CLK(n1552), .Q(n667), .QN(
        \fpu_add_frac_dp/n5632 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[45]  ( .D(
        \fpu_add_frac_dp/n3685 ), .CLK(n1552), .Q(n100), .QN(
        \fpu_add_frac_dp/n2387 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[44]  ( .D(
        \fpu_add_frac_dp/n3686 ), .CLK(n1552), .Q(n665), .QN(
        \fpu_add_frac_dp/n5609 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[43]  ( .D(
        \fpu_add_frac_dp/n3687 ), .CLK(n1552), .Q(n83), .QN(
        \fpu_add_frac_dp/n2537 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[42]  ( .D(
        \fpu_add_frac_dp/n3688 ), .CLK(n1552), .Q(n38), .QN(
        \fpu_add_frac_dp/n2481 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[41]  ( .D(
        \fpu_add_frac_dp/n3689 ), .CLK(n1552), .Q(n117), .QN(
        \fpu_add_frac_dp/n2361 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[40]  ( .D(
        \fpu_add_frac_dp/n3690 ), .CLK(n1553), .Q(n673), .QN(
        \fpu_add_frac_dp/n658 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[39]  ( .D(
        \fpu_add_frac_dp/n3691 ), .CLK(n1553), .Q(n19), .QN(
        \fpu_add_frac_dp/n2404 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[38]  ( .D(
        \fpu_add_frac_dp/n3692 ), .CLK(n1553), .Q(n86), .QN(
        \fpu_add_frac_dp/n2336 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[37]  ( .D(
        \fpu_add_frac_dp/n3693 ), .CLK(n1553), .Q(n177), .QN(
        \fpu_add_frac_dp/n659 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[36]  ( .D(
        \fpu_add_frac_dp/n3694 ), .CLK(n1553), .Q(\fpu_add_frac_dp/n2332 ), 
        .QN(n716) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[35]  ( .D(
        \fpu_add_frac_dp/n3695 ), .CLK(n1553), .Q(\fpu_add_frac_dp/n2406 ), 
        .QN(\fpu_add_frac_dp/n1335 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[34]  ( .D(
        \fpu_add_frac_dp/n3696 ), .CLK(n1553), .Q(\fpu_add_frac_dp/n2289 ), 
        .QN(n1271) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[33]  ( .D(
        \fpu_add_frac_dp/n3697 ), .CLK(n1553), .Q(\fpu_add_frac_dp/n2342 ), 
        .QN(\fpu_add_frac_dp/n1333 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[32]  ( .D(
        \fpu_add_frac_dp/n3698 ), .CLK(n1553), .Q(\fpu_add_frac_dp/n2403 ), 
        .QN(\fpu_add_frac_dp/n1332 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[31]  ( .D(
        \fpu_add_frac_dp/n3699 ), .CLK(n1553), .Q(\fpu_add_frac_dp/n2335 ), 
        .QN(n839) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[30]  ( .D(
        \fpu_add_frac_dp/n3700 ), .CLK(n1553), .Q(n262), .QN(
        \fpu_add_frac_dp/n2363 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[29]  ( .D(
        \fpu_add_frac_dp/n3701 ), .CLK(n1553), .Q(n101), .QN(
        \fpu_add_frac_dp/n2496 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[28]  ( .D(
        \fpu_add_frac_dp/n3702 ), .CLK(n1553), .Q(n329), .QN(
        \fpu_add_frac_dp/n660 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[27]  ( .D(
        \fpu_add_frac_dp/n3703 ), .CLK(n1553), .Q(\fpu_add_frac_dp/n2313 ), 
        .QN(n346) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[26]  ( .D(
        \fpu_add_frac_dp/n3704 ), .CLK(n1554), .Q(\fpu_add_frac_dp/n2402 ), 
        .QN(n710) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[25]  ( .D(
        \fpu_add_frac_dp/n3705 ), .CLK(n1554), .Q(n116), .QN(
        \fpu_add_frac_dp/n2470 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[24]  ( .D(
        \fpu_add_frac_dp/n3706 ), .CLK(n1554), .Q(n331), .QN(
        \fpu_add_frac_dp/n5619 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[23]  ( .D(
        \fpu_add_frac_dp/n3707 ), .CLK(n1554), .Q(n74), .QN(
        \fpu_add_frac_dp/n2409 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[22]  ( .D(
        \fpu_add_frac_dp/n3708 ), .CLK(n1554), .Q(n594), .QN(
        \fpu_add_frac_dp/n662 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[21]  ( .D(
        \fpu_add_frac_dp/n3709 ), .CLK(n1554), .Q(\fpu_add_frac_dp/n2405 ), 
        .QN(n1087) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[20]  ( .D(
        \fpu_add_frac_dp/n3710 ), .CLK(n1554), .Q(\fpu_add_frac_dp/n2339 ), 
        .QN(n447) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[19]  ( .D(
        \fpu_add_frac_dp/n3711 ), .CLK(n1554), .Q(n664), .QN(
        \fpu_add_frac_dp/n2411 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[18]  ( .D(
        \fpu_add_frac_dp/n3712 ), .CLK(n1554), .Q(n111), .QN(
        \fpu_add_frac_dp/n2344 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[17]  ( .D(
        \fpu_add_frac_dp/n3713 ), .CLK(n1554), .Q(n43), .QN(
        \fpu_add_frac_dp/n2495 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[16]  ( .D(
        \fpu_add_frac_dp/n3714 ), .CLK(n1554), .Q(n328), .QN(
        \fpu_add_frac_dp/n664 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[15]  ( .D(
        \fpu_add_frac_dp/n3715 ), .CLK(n1554), .Q(\fpu_add_frac_dp/n2400 ), 
        .QN(\fpu_add_frac_dp/n1315 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[14]  ( .D(
        \fpu_add_frac_dp/n3716 ), .CLK(n1554), .Q(\fpu_add_frac_dp/n2330 ), 
        .QN(\fpu_add_frac_dp/n1314 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[13]  ( .D(
        \fpu_add_frac_dp/n3717 ), .CLK(n1554), .Q(n597), .QN(
        \fpu_add_frac_dp/n2437 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[12]  ( .D(
        \fpu_add_frac_dp/n3718 ), .CLK(n1555), .Q(n37) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[11]  ( .D(
        \fpu_add_frac_dp/n3719 ), .CLK(n1555), .Q(n691), .QN(
        \fpu_add_frac_dp/n2519 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[10]  ( .D(
        \fpu_add_frac_dp/n3720 ), .CLK(n1555), .Q(n12), .QN(
        \fpu_add_frac_dp/n5610 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[9]  ( .D(
        \fpu_add_frac_dp/n3721 ), .CLK(n1555), .Q(n34), .QN(
        \fpu_add_frac_dp/n2494 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[8]  ( .D(
        \fpu_add_frac_dp/n3722 ), .CLK(n1555), .Q(n623), .QN(
        \fpu_add_frac_dp/n666 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[7]  ( .D(
        \fpu_add_frac_dp/n3723 ), .CLK(n1555), .Q(n33), .QN(
        \fpu_add_frac_dp/n2513 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[6]  ( .D(
        \fpu_add_frac_dp/n3724 ), .CLK(n1555), .Q(n173), .QN(
        \fpu_add_frac_dp/n668 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[5]  ( .D(
        \fpu_add_frac_dp/n3725 ), .CLK(n1555), .Q(n626), .QN(
        \fpu_add_frac_dp/n2520 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[4]  ( .D(
        \fpu_add_frac_dp/n3726 ), .CLK(n1555), .Q(n90) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[3]  ( .D(
        \fpu_add_frac_dp/n3727 ), .CLK(n1555), .Q(n671), .QN(
        \fpu_add_frac_dp/n670 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[2]  ( .D(
        \fpu_add_frac_dp/n3728 ), .CLK(n1555), .Q(n282), .QN(
        \fpu_add_frac_dp/n2447 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[1]  ( .D(
        \fpu_add_frac_dp/n3729 ), .CLK(n1555), .Q(n103), .QN(
        \fpu_add_frac_dp/n5642 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_ld0_frac/q_reg[0]  ( .D(
        \fpu_add_frac_dp/n3730 ), .CLK(n1555), .Q(n652) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[62]  ( .D(\fpu_add_frac_dp/n3794 ), .CLK(n1493), .Q(n453), .QN(\fpu_add_frac_dp/n673 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[61]  ( .D(\fpu_add_frac_dp/n3795 ), .CLK(n1493), .Q(n768), .QN(\fpu_add_frac_dp/n674 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[60]  ( .D(\fpu_add_frac_dp/n3796 ), .CLK(n1493), .Q(n769), .QN(\fpu_add_frac_dp/n675 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[59]  ( .D(\fpu_add_frac_dp/n3797 ), .CLK(n1493), .Q(n770), .QN(\fpu_add_frac_dp/n676 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[58]  ( .D(\fpu_add_frac_dp/n3798 ), .CLK(n1493), .Q(n771), .QN(\fpu_add_frac_dp/n677 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[57]  ( .D(\fpu_add_frac_dp/n3799 ), .CLK(n1493), .Q(n772), .QN(\fpu_add_frac_dp/n678 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[56]  ( .D(\fpu_add_frac_dp/n3800 ), .CLK(n1493), .Q(n773), .QN(\fpu_add_frac_dp/n679 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[55]  ( .D(\fpu_add_frac_dp/n3801 ), .CLK(n1492), .Q(n774), .QN(\fpu_add_frac_dp/n680 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[54]  ( .D(\fpu_add_frac_dp/n3802 ), .CLK(n1492), .Q(n775), .QN(\fpu_add_frac_dp/n681 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[53]  ( .D(\fpu_add_frac_dp/n3803 ), .CLK(n1492), .Q(n776), .QN(\fpu_add_frac_dp/n682 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[52]  ( .D(\fpu_add_frac_dp/n3804 ), .CLK(n1492), .Q(n777), .QN(\fpu_add_frac_dp/n683 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[51]  ( .D(\fpu_add_frac_dp/n3805 ), .CLK(n1492), .Q(n778), .QN(\fpu_add_frac_dp/n684 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[50]  ( .D(\fpu_add_frac_dp/n3806 ), .CLK(n1492), .Q(n779), .QN(\fpu_add_frac_dp/n685 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[49]  ( .D(\fpu_add_frac_dp/n3807 ), .CLK(n1492), .Q(n780), .QN(\fpu_add_frac_dp/n686 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[48]  ( .D(\fpu_add_frac_dp/n3808 ), .CLK(n1491), .Q(n781), .QN(\fpu_add_frac_dp/n687 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[47]  ( .D(\fpu_add_frac_dp/n3809 ), .CLK(n1491), .Q(n782), .QN(\fpu_add_frac_dp/n688 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[46]  ( .D(\fpu_add_frac_dp/n3810 ), .CLK(n1491), .Q(n783), .QN(\fpu_add_frac_dp/n689 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[45]  ( .D(\fpu_add_frac_dp/n3811 ), .CLK(n1491), .Q(n784), .QN(\fpu_add_frac_dp/n690 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[44]  ( .D(\fpu_add_frac_dp/n3812 ), .CLK(n1491), .Q(n785), .QN(\fpu_add_frac_dp/n691 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[43]  ( .D(\fpu_add_frac_dp/n3813 ), .CLK(n1491), .Q(n786), .QN(\fpu_add_frac_dp/n692 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[42]  ( .D(\fpu_add_frac_dp/n3814 ), .CLK(n1491), .Q(n787), .QN(\fpu_add_frac_dp/n693 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[41]  ( .D(\fpu_add_frac_dp/n3815 ), .CLK(n1490), .Q(n788), .QN(\fpu_add_frac_dp/n694 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[40]  ( .D(\fpu_add_frac_dp/n3816 ), .CLK(n1490), .Q(n789), .QN(\fpu_add_frac_dp/n695 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[39]  ( .D(\fpu_add_frac_dp/n3817 ), .CLK(n1490), .Q(n790), .QN(\fpu_add_frac_dp/n696 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[38]  ( .D(\fpu_add_frac_dp/n3818 ), .CLK(n1490), .Q(n791), .QN(\fpu_add_frac_dp/n697 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[37]  ( .D(\fpu_add_frac_dp/n3819 ), .CLK(n1490), .Q(n792), .QN(\fpu_add_frac_dp/n698 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[36]  ( .D(\fpu_add_frac_dp/n3820 ), .CLK(n1490), .Q(n793), .QN(\fpu_add_frac_dp/n699 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[35]  ( .D(\fpu_add_frac_dp/n3821 ), .CLK(n1490), .Q(n794), .QN(\fpu_add_frac_dp/n700 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[34]  ( .D(\fpu_add_frac_dp/n3822 ), .CLK(n1489), .Q(n795), .QN(\fpu_add_frac_dp/n701 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[33]  ( .D(\fpu_add_frac_dp/n3823 ), .CLK(n1489), .Q(n796), .QN(\fpu_add_frac_dp/n702 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[32]  ( .D(\fpu_add_frac_dp/n3824 ), .CLK(n1489), .Q(n797), .QN(\fpu_add_frac_dp/n703 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[31]  ( .D(\fpu_add_frac_dp/n3825 ), .CLK(n1489), .Q(n798), .QN(\fpu_add_frac_dp/n704 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[30]  ( .D(\fpu_add_frac_dp/n3826 ), .CLK(n1489), .Q(n799), .QN(\fpu_add_frac_dp/n705 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[29]  ( .D(\fpu_add_frac_dp/n3827 ), .CLK(n1489), .Q(n800), .QN(\fpu_add_frac_dp/n706 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[28]  ( .D(\fpu_add_frac_dp/n3828 ), .CLK(n1489), .Q(n801), .QN(\fpu_add_frac_dp/n707 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[27]  ( .D(\fpu_add_frac_dp/n3829 ), .CLK(n1488), .Q(n802), .QN(\fpu_add_frac_dp/n708 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[26]  ( .D(\fpu_add_frac_dp/n3830 ), .CLK(n1488), .Q(n803), .QN(\fpu_add_frac_dp/n709 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[25]  ( .D(\fpu_add_frac_dp/n3831 ), .CLK(n1488), .Q(n804), .QN(\fpu_add_frac_dp/n710 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[24]  ( .D(\fpu_add_frac_dp/n3832 ), .CLK(n1488), .Q(n805), .QN(\fpu_add_frac_dp/n711 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[23]  ( .D(\fpu_add_frac_dp/n3833 ), .CLK(n1488), .Q(n806), .QN(\fpu_add_frac_dp/n712 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[22]  ( .D(\fpu_add_frac_dp/n3834 ), .CLK(n1488), .Q(n807), .QN(\fpu_add_frac_dp/n713 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[21]  ( .D(\fpu_add_frac_dp/n3835 ), .CLK(n1488), .Q(n808), .QN(\fpu_add_frac_dp/n714 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[20]  ( .D(\fpu_add_frac_dp/n3836 ), .CLK(n1487), .Q(n809), .QN(\fpu_add_frac_dp/n715 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[19]  ( .D(\fpu_add_frac_dp/n3837 ), .CLK(n1487), .Q(n810), .QN(\fpu_add_frac_dp/n716 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[18]  ( .D(\fpu_add_frac_dp/n3838 ), .CLK(n1487), .Q(n811), .QN(\fpu_add_frac_dp/n717 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[17]  ( .D(\fpu_add_frac_dp/n3839 ), .CLK(n1487), .Q(n812), .QN(\fpu_add_frac_dp/n718 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[16]  ( .D(\fpu_add_frac_dp/n3840 ), .CLK(n1492), .Q(n813), .QN(\fpu_add_frac_dp/n719 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[15]  ( .D(\fpu_add_frac_dp/n3841 ), .CLK(n1548), .Q(n814), .QN(\fpu_add_frac_dp/n720 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[14]  ( .D(\fpu_add_frac_dp/n3842 ), .CLK(n1547), .Q(n815), .QN(\fpu_add_frac_dp/n721 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[13]  ( .D(\fpu_add_frac_dp/n3843 ), .CLK(n1547), .Q(n816), .QN(\fpu_add_frac_dp/n722 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[12]  ( .D(\fpu_add_frac_dp/n3844 ), .CLK(n1547), .Q(n817), .QN(\fpu_add_frac_dp/n723 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[11]  ( .D(\fpu_add_frac_dp/n3845 ), .CLK(n1547), .Q(n818), .QN(\fpu_add_frac_dp/n724 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[10]  ( .D(\fpu_add_frac_dp/n3846 ), .CLK(n1547), .Q(n819), .QN(\fpu_add_frac_dp/n725 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[9]  ( .D(\fpu_add_frac_dp/n3847 ), 
        .CLK(n1547), .Q(n820), .QN(\fpu_add_frac_dp/n726 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[8]  ( .D(\fpu_add_frac_dp/n3848 ), 
        .CLK(n1547), .Q(n821), .QN(\fpu_add_frac_dp/n727 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[7]  ( .D(\fpu_add_frac_dp/n3849 ), 
        .CLK(n1546), .Q(n822), .QN(\fpu_add_frac_dp/n728 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[6]  ( .D(\fpu_add_frac_dp/n3850 ), 
        .CLK(n1546), .Q(n823), .QN(\fpu_add_frac_dp/n729 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[5]  ( .D(\fpu_add_frac_dp/n3851 ), 
        .CLK(n1546), .Q(n824), .QN(\fpu_add_frac_dp/n730 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[4]  ( .D(\fpu_add_frac_dp/n3852 ), 
        .CLK(n1546), .Q(n825), .QN(\fpu_add_frac_dp/n731 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[3]  ( .D(\fpu_add_frac_dp/n3853 ), 
        .CLK(n1546), .Q(n826), .QN(\fpu_add_frac_dp/n732 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[2]  ( .D(\fpu_add_frac_dp/n3854 ), 
        .CLK(n1546), .Q(n827), .QN(\fpu_add_frac_dp/n733 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[1]  ( .D(\fpu_add_frac_dp/n3855 ), 
        .CLK(n1546), .Q(n828), .QN(\fpu_add_frac_dp/n734 ) );
  DFFX1 \fpu_add_frac_dp/i_a3stg_frac1/q_reg[0]  ( .D(\fpu_add_frac_dp/n3856 ), 
        .CLK(n1545), .Q(n465), .QN(\fpu_add_frac_dp/n735 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[63]  ( .D(
        \fpu_add_frac_dp/n3857 ), .CLK(n1486), .Q(n15), .QN(
        \fpu_add_frac_dp/n2262 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[62]  ( .D(
        \fpu_add_frac_dp/n3858 ), .CLK(n1486), .Q(n16), .QN(
        \fpu_add_frac_dp/n2270 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[61]  ( .D(
        \fpu_add_frac_dp/n3859 ), .CLK(n1485), .Q(n3), .QN(
        \fpu_add_frac_dp/n2282 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[60]  ( .D(
        \fpu_add_frac_dp/n3860 ), .CLK(n1485), .Q(n156), .QN(
        \fpu_add_frac_dp/n2317 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[59]  ( .D(
        \fpu_add_frac_dp/n3861 ), .CLK(n1485), .Q(n68), .QN(
        \fpu_add_frac_dp/n2269 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[58]  ( .D(
        \fpu_add_frac_dp/n3862 ), .CLK(n1485), .Q(
        \fpu_add_frac_dp/a2stg_frac2a[58] ), .QN(\fpu_add_frac_dp/n2281 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[57]  ( .D(
        \fpu_add_frac_dp/n3863 ), .CLK(n1485), .Q(n157), .QN(
        \fpu_add_frac_dp/n2314 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[56]  ( .D(
        \fpu_add_frac_dp/n3864 ), .CLK(n1485), .Q(n4), .QN(
        \fpu_add_frac_dp/n2331 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[55]  ( .D(
        \fpu_add_frac_dp/n3865 ), .CLK(n1485), .Q(n98), .QN(
        \fpu_add_frac_dp/n2430 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[54]  ( .D(
        \fpu_add_frac_dp/n3866 ), .CLK(n1485), .Q(n97), .QN(
        \fpu_add_frac_dp/n2429 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[53]  ( .D(
        \fpu_add_frac_dp/n3867 ), .CLK(n1485), .Q(n613), .QN(
        \fpu_add_frac_dp/n2428 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[52]  ( .D(
        \fpu_add_frac_dp/n3868 ), .CLK(n1485), .Q(n95), .QN(
        \fpu_add_frac_dp/n2427 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[51]  ( .D(
        \fpu_add_frac_dp/n3869 ), .CLK(n1485), .Q(n632), .QN(
        \fpu_add_frac_dp/n2341 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[50]  ( .D(
        \fpu_add_frac_dp/n3870 ), .CLK(n1485), .Q(n630), .QN(
        \fpu_add_frac_dp/n2395 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[49]  ( .D(
        \fpu_add_frac_dp/n3871 ), .CLK(n1485), .Q(n631), .QN(
        \fpu_add_frac_dp/n2426 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[48]  ( .D(
        \fpu_add_frac_dp/n3872 ), .CLK(n1485), .Q(n96), .QN(
        \fpu_add_frac_dp/n2425 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[47]  ( .D(
        \fpu_add_frac_dp/n3873 ), .CLK(n1484), .Q(n217), .QN(
        \fpu_add_frac_dp/n2518 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[46]  ( .D(
        \fpu_add_frac_dp/n3874 ), .CLK(n1484), .Q(n280), .QN(
        \fpu_add_frac_dp/n2517 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[45]  ( .D(
        \fpu_add_frac_dp/n3875 ), .CLK(n1484), .Q(n281), .QN(
        \fpu_add_frac_dp/n2516 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[44]  ( .D(
        \fpu_add_frac_dp/n3876 ), .CLK(n1484), .Q(n638), .QN(
        \fpu_add_frac_dp/n2515 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[43]  ( .D(
        \fpu_add_frac_dp/n3877 ), .CLK(n1484), .Q(n174), .QN(
        \fpu_add_frac_dp/n2480 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[42]  ( .D(
        \fpu_add_frac_dp/n3878 ), .CLK(n1484), .Q(n70), .QN(
        \fpu_add_frac_dp/n2479 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[41]  ( .D(
        \fpu_add_frac_dp/n3879 ), .CLK(n1484), .Q(\fpu_add_frac_dp/n2380 ), 
        .QN(\fpu_add_frac_dp/n1215 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[40]  ( .D(
        \fpu_add_frac_dp/n3880 ), .CLK(n1484), .Q(n168), .QN(
        \fpu_add_frac_dp/n2497 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[39]  ( .D(
        \fpu_add_frac_dp/n3881 ), .CLK(n1484), .Q(n271), .QN(
        \fpu_add_frac_dp/n736 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[38]  ( .D(
        \fpu_add_frac_dp/n3882 ), .CLK(n1484), .Q(n23) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[37]  ( .D(
        \fpu_add_frac_dp/n3883 ), .CLK(n1484), .Q(n162) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[36]  ( .D(
        \fpu_add_frac_dp/n3884 ), .CLK(n1484), .Q(n6) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[35]  ( .D(
        \fpu_add_frac_dp/n3885 ), .CLK(n1484), .Q(n205), .QN(
        \fpu_add_frac_dp/n2424 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[34]  ( .D(
        \fpu_add_frac_dp/n3886 ), .CLK(n1484), .Q(\fpu_add_frac_dp/n2393 ), 
        .QN(\fpu_add_frac_dp/n1213 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[33]  ( .D(
        \fpu_add_frac_dp/n3887 ), .CLK(n1483), .Q(n278), .QN(
        \fpu_add_frac_dp/n741 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[32]  ( .D(
        \fpu_add_frac_dp/n3888 ), .CLK(n1483), .Q(n218) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[31]  ( .D(
        \fpu_add_frac_dp/n3889 ), .CLK(n1483), .Q(n696), .QN(
        \fpu_add_frac_dp/n743 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[30]  ( .D(
        \fpu_add_frac_dp/n3890 ), .CLK(n1483), .Q(n678), .QN(
        \fpu_add_frac_dp/n744 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[29]  ( .D(
        \fpu_add_frac_dp/n3891 ), .CLK(n1483), .Q(n679), .QN(
        \fpu_add_frac_dp/n745 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[28]  ( .D(
        \fpu_add_frac_dp/n3892 ), .CLK(n1483), .Q(n106) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[27]  ( .D(
        \fpu_add_frac_dp/n3893 ), .CLK(n1483), .Q(n720), .QN(
        \fpu_add_frac_dp/n747 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[26]  ( .D(
        \fpu_add_frac_dp/n3894 ), .CLK(n1483), .Q(n312) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[25]  ( .D(
        \fpu_add_frac_dp/n3895 ), .CLK(n1483), .Q(n932), .QN(
        \fpu_add_frac_dp/n749 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[24]  ( .D(
        \fpu_add_frac_dp/n3896 ), .CLK(n1483), .Q(n929), .QN(
        \fpu_add_frac_dp/n750 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[23]  ( .D(
        \fpu_add_frac_dp/n3897 ), .CLK(n1483), .Q(n931), .QN(
        \fpu_add_frac_dp/n751 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[22]  ( .D(
        \fpu_add_frac_dp/n3898 ), .CLK(n1483), .Q(n934), .QN(
        \fpu_add_frac_dp/n752 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[21]  ( .D(
        \fpu_add_frac_dp/n3899 ), .CLK(n1483), .Q(n131) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[20]  ( .D(
        \fpu_add_frac_dp/n3900 ), .CLK(n1483), .Q(n314) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[19]  ( .D(
        \fpu_add_frac_dp/n3901 ), .CLK(n1482), .Q(n717), .QN(
        \fpu_add_frac_dp/n755 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[18]  ( .D(
        \fpu_add_frac_dp/n3902 ), .CLK(n1482), .Q(n1152), .QN(
        \fpu_add_frac_dp/n756 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[17]  ( .D(
        \fpu_add_frac_dp/n3903 ), .CLK(n1482), .Q(n1151), .QN(
        \fpu_add_frac_dp/n757 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[16]  ( .D(
        \fpu_add_frac_dp/n3904 ), .CLK(n1482), .Q(n930), .QN(
        \fpu_add_frac_dp/n758 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[15]  ( .D(
        \fpu_add_frac_dp/n3905 ), .CLK(n1482), .Q(n935), .QN(
        \fpu_add_frac_dp/n759 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[14]  ( .D(
        \fpu_add_frac_dp/n3906 ), .CLK(n1482), .Q(n425), .QN(
        \fpu_add_frac_dp/n760 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[13]  ( .D(
        \fpu_add_frac_dp/n3907 ), .CLK(n1482), .Q(n721), .QN(
        \fpu_add_frac_dp/n761 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[12]  ( .D(
        \fpu_add_frac_dp/n3908 ), .CLK(n1482), .Q(n150), .QN(
        \fpu_add_frac_dp/n762 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[11]  ( .D(
        \fpu_add_frac_dp/n3909 ), .CLK(n1482), .Q(n627), .QN(
        \fpu_add_frac_dp/n763 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[10]  ( .D(
        \fpu_add_frac_dp/n3910 ), .CLK(n1482), .Q(n161) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[9]  ( .D(\fpu_add_frac_dp/n3911 ), .CLK(n1482), .Q(n75) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[8]  ( .D(\fpu_add_frac_dp/n3912 ), .CLK(n1482), .Q(n659), .QN(\fpu_add_frac_dp/n766 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[7]  ( .D(\fpu_add_frac_dp/n3913 ), .CLK(n1482), .Q(n901), .QN(\fpu_add_frac_dp/n767 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[6]  ( .D(\fpu_add_frac_dp/n3914 ), .CLK(n1482), .Q(n655), .QN(\fpu_add_frac_dp/n768 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[5]  ( .D(\fpu_add_frac_dp/n3915 ), .CLK(n1481), .Q(n898), .QN(\fpu_add_frac_dp/n769 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[4]  ( .D(\fpu_add_frac_dp/n3916 ), .CLK(n1481), .Q(n660), .QN(\fpu_add_frac_dp/n770 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[3]  ( .D(\fpu_add_frac_dp/n3917 ), .CLK(n1481), .Q(n899), .QN(\fpu_add_frac_dp/n771 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[2]  ( .D(\fpu_add_frac_dp/n3918 ), .CLK(n1481), .Q(n690), .QN(\fpu_add_frac_dp/n772 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[1]  ( .D(\fpu_add_frac_dp/n3919 ), .CLK(n1481), .Q(n902), .QN(\fpu_add_frac_dp/n773 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2a/q_reg[0]  ( .D(\fpu_add_frac_dp/n3920 ), .CLK(n1481), .Q(n896), .QN(\fpu_add_frac_dp/n774 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[63]  ( .D(\fpu_add_frac_dp/n3921 ), .CLK(n1481), .Q(n1101), .QN(\fpu_add_frac_dp/n2498 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[62]  ( .D(\fpu_add_frac_dp/n3922 ), .CLK(n1481), .Q(n142), .QN(\fpu_add_frac_dp/n2502 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[61]  ( .D(\fpu_add_frac_dp/n3923 ), .CLK(n1481), .Q(n706), .QN(\fpu_add_frac_dp/n2506 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[60]  ( .D(\fpu_add_frac_dp/n3924 ), .CLK(n1480), .Q(\fpu_add_frac_dp/n2384 ), .QN(n1009) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[59]  ( .D(\fpu_add_frac_dp/n3925 ), .CLK(n1480), .Q(\fpu_add_frac_dp/n2391 ), .QN(n153) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[58]  ( .D(\fpu_add_frac_dp/n3926 ), .CLK(n1480), .Q(\fpu_add_frac_dp/n2390 ), .QN(n561) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[57]  ( .D(\fpu_add_frac_dp/n3927 ), .CLK(n1480), .Q(\fpu_add_frac_dp/n2392 ), .QN(n62) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[56]  ( .D(\fpu_add_frac_dp/n3928 ), .CLK(n1480), .Q(n343), .QN(\fpu_add_frac_dp/n2357 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[55]  ( .D(\fpu_add_frac_dp/n3929 ), .CLK(n1480), .Q(n1118), .QN(\fpu_add_frac_dp/n2431 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[54]  ( .D(\fpu_add_frac_dp/n3930 ), .CLK(n1480), .Q(n1103), .QN(\fpu_add_frac_dp/n2418 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[53]  ( .D(\fpu_add_frac_dp/n3931 ), .CLK(n1480), .Q(n1100), .QN(\fpu_add_frac_dp/n2351 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[52]  ( .D(\fpu_add_frac_dp/n3932 ), .CLK(n1481), .Q(n1110), .QN(\fpu_add_frac_dp/n2505 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[51]  ( .D(\fpu_add_frac_dp/n3933 ), .CLK(n1480), .Q(n708), .QN(\fpu_add_frac_dp/n2501 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[50]  ( .D(\fpu_add_frac_dp/n3934 ), .CLK(n1480), .Q(n345), .QN(\fpu_add_frac_dp/n2512 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[49]  ( .D(\fpu_add_frac_dp/n3935 ), .CLK(n1481), .Q(n144), .QN(\fpu_add_frac_dp/n2509 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[48]  ( .D(\fpu_add_frac_dp/n3936 ), .CLK(n1480), .Q(n59), .QN(\fpu_add_frac_dp/n2500 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[47]  ( .D(\fpu_add_frac_dp/n3937 ), .CLK(n1479), .Q(n707), .QN(\fpu_add_frac_dp/n2303 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[46]  ( .D(\fpu_add_frac_dp/n3938 ), .CLK(n1480), .Q(n344), .QN(\fpu_add_frac_dp/n2356 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[45]  ( .D(\fpu_add_frac_dp/n3939 ), .CLK(n1479), .Q(n143), .QN(\fpu_add_frac_dp/n2508 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[44]  ( .D(\fpu_add_frac_dp/n3940 ), .CLK(n1479), .Q(n58), .QN(\fpu_add_frac_dp/n2504 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[43]  ( .D(\fpu_add_frac_dp/n3941 ), .CLK(n1480), .Q(n1117), .QN(\fpu_add_frac_dp/n2276 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[42]  ( .D(\fpu_add_frac_dp/n3942 ), .CLK(n1479), .Q(n1102), .QN(\fpu_add_frac_dp/n2302 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[41]  ( .D(\fpu_add_frac_dp/n3943 ), .CLK(n1479), .Q(n1099), .QN(\fpu_add_frac_dp/n2422 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[40]  ( .D(\fpu_add_frac_dp/n3944 ), .CLK(n1496), .Q(n1109), .QN(\fpu_add_frac_dp/n2355 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[39]  ( .D(\fpu_add_frac_dp/n3945 ), .CLK(n1496), .Q(n1116), .QN(\fpu_add_frac_dp/n2275 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[38]  ( .D(\fpu_add_frac_dp/n3946 ), .CLK(n1496), .Q(n1098), .QN(\fpu_add_frac_dp/n2301 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[37]  ( .D(\fpu_add_frac_dp/n3947 ), .CLK(n1496), .Q(n1097), .QN(\fpu_add_frac_dp/n2421 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[36]  ( .D(\fpu_add_frac_dp/n3948 ), .CLK(n1496), .Q(n1108), .QN(\fpu_add_frac_dp/n2511 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[35]  ( .D(\fpu_add_frac_dp/n3949 ), .CLK(n1496), .Q(n1115), .QN(\fpu_add_frac_dp/n2435 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[34]  ( .D(\fpu_add_frac_dp/n3950 ), .CLK(n1496), .Q(n1096), .QN(\fpu_add_frac_dp/n2354 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[33]  ( .D(\fpu_add_frac_dp/n3951 ), .CLK(n1496), .Q(n1095), .QN(\fpu_add_frac_dp/n2274 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[32]  ( .D(\fpu_add_frac_dp/n3952 ), .CLK(n1496), .Q(n1107), .QN(\fpu_add_frac_dp/n2300 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[31]  ( .D(\fpu_add_frac_dp/n3953 ), .CLK(n1496), .Q(n1114), .QN(\fpu_add_frac_dp/n2510 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[30]  ( .D(\fpu_add_frac_dp/n3954 ), .CLK(n1496), .Q(n1094), .QN(\fpu_add_frac_dp/n2503 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[29]  ( .D(\fpu_add_frac_dp/n3955 ), .CLK(n1496), .Q(n1106), .QN(\fpu_add_frac_dp/n2499 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[28]  ( .D(\fpu_add_frac_dp/n3956 ), .CLK(n1496), .Q(n424), .QN(\fpu_add_frac_dp/n2507 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[27]  ( .D(\fpu_add_frac_dp/n3957 ), .CLK(n1496), .Q(n723), .QN(\fpu_add_frac_dp/n2419 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[26]  ( .D(\fpu_add_frac_dp/n3958 ), .CLK(n1495), .Q(n1113), .QN(\fpu_add_frac_dp/n2299 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[25]  ( .D(\fpu_add_frac_dp/n3959 ), .CLK(n1495), .Q(n1093), .QN(\fpu_add_frac_dp/n2420 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[24]  ( .D(\fpu_add_frac_dp/n3960 ), .CLK(n1495), .Q(n1105), .QN(\fpu_add_frac_dp/n2273 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[23]  ( .D(\fpu_add_frac_dp/n3961 ), .CLK(n1495), .Q(n426), .QN(\fpu_add_frac_dp/n2352 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[22]  ( .D(\fpu_add_frac_dp/n3962 ), .CLK(n1495), .Q(n724), .QN(\fpu_add_frac_dp/n2353 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[21]  ( .D(\fpu_add_frac_dp/n3963 ), .CLK(n1495), .Q(n1112), .QN(\fpu_add_frac_dp/n2434 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[20]  ( .D(\fpu_add_frac_dp/n3964 ), .CLK(n1495), .Q(n1092), .QN(\fpu_add_frac_dp/n2433 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[19]  ( .D(\fpu_add_frac_dp/n3965 ), .CLK(n1495), .Q(n1104), .QN(\fpu_add_frac_dp/n2297 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[18]  ( .D(\fpu_add_frac_dp/n3966 ), .CLK(n1495), .Q(n423), .QN(\fpu_add_frac_dp/n2272 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[17]  ( .D(\fpu_add_frac_dp/n3967 ), .CLK(n1495), .Q(n722), .QN(\fpu_add_frac_dp/n2298 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[16]  ( .D(\fpu_add_frac_dp/n3968 ), .CLK(n1495), .Q(n1123), .QN(\fpu_add_frac_dp/n2359 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[15]  ( .D(\fpu_add_frac_dp/n3969 ), .CLK(n1495), .Q(n1125), .QN(\fpu_add_frac_dp/n2432 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[14]  ( .D(\fpu_add_frac_dp/n3970 ), .CLK(n1495), .Q(n1122), .QN(\fpu_add_frac_dp/n2362 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[13]  ( .D(\fpu_add_frac_dp/n3971 ), .CLK(n1495), .Q(n1091), .QN(\fpu_add_frac_dp/n2304 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[12]  ( .D(\fpu_add_frac_dp/n3972 ), .CLK(n1494), .Q(\fpu_add_frac_dp/n2389 ), .QN(n904) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[11]  ( .D(\fpu_add_frac_dp/n3973 ), .CLK(n1494), .Q(n1111), .QN(\fpu_add_frac_dp/n2277 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[10]  ( .D(\fpu_add_frac_dp/n3974 ), .CLK(n1494), .Q(n1142), .QN(\fpu_add_frac_dp/n2531 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[9]  ( .D(\fpu_add_frac_dp/n3975 ), 
        .CLK(n1494), .Q(n1141), .QN(\fpu_add_frac_dp/n2530 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[8]  ( .D(\fpu_add_frac_dp/n3976 ), 
        .CLK(n1494), .Q(n1140), .QN(\fpu_add_frac_dp/n2529 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[7]  ( .D(\fpu_add_frac_dp/n3977 ), 
        .CLK(n1494), .Q(n1139), .QN(\fpu_add_frac_dp/n2528 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[6]  ( .D(\fpu_add_frac_dp/n3978 ), 
        .CLK(n1494), .Q(n1138), .QN(\fpu_add_frac_dp/n2527 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[5]  ( .D(\fpu_add_frac_dp/n3979 ), 
        .CLK(n1494), .Q(n1149), .QN(\fpu_add_frac_dp/n2526 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[4]  ( .D(\fpu_add_frac_dp/n3980 ), 
        .CLK(n1494), .Q(n1137), .QN(\fpu_add_frac_dp/n2525 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[3]  ( .D(\fpu_add_frac_dp/n3981 ), 
        .CLK(n1494), .Q(n1136), .QN(\fpu_add_frac_dp/n2524 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[2]  ( .D(\fpu_add_frac_dp/n3982 ), 
        .CLK(n1494), .Q(n1135), .QN(\fpu_add_frac_dp/n2523 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[1]  ( .D(\fpu_add_frac_dp/n3983 ), 
        .CLK(n1494), .Q(n1134), .QN(\fpu_add_frac_dp/n2522 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac2/q_reg[0]  ( .D(\fpu_add_frac_dp/n3984 ), 
        .CLK(n1494), .Q(n1196), .QN(\fpu_add_frac_dp/n2539 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[63]  ( .D(\fpu_add_frac_dp/n3985 ), .CLK(n1494), .Q(n850), .QN(\fpu_add_frac_dp/n5640 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[62]  ( .D(\fpu_add_frac_dp/n3986 ), .CLK(n1493), .Q(n226) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[61]  ( .D(\fpu_add_frac_dp/n3987 ), .CLK(n1493), .Q(n195) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[60]  ( .D(\fpu_add_frac_dp/n3988 ), .CLK(n1493), .Q(n317), .QN(\fpu_add_frac_dp/n777 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[59]  ( .D(\fpu_add_frac_dp/n3989 ), .CLK(n1493), .Q(n293), .QN(\fpu_add_frac_dp/n778 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[58]  ( .D(\fpu_add_frac_dp/n3990 ), .CLK(n1493), .Q(n334), .QN(\fpu_add_frac_dp/n779 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[57]  ( .D(\fpu_add_frac_dp/n3991 ), .CLK(n1493), .Q(n332), .QN(\fpu_add_frac_dp/n780 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[56]  ( .D(\fpu_add_frac_dp/n3992 ), .CLK(n1493), .Q(n294), .QN(\fpu_add_frac_dp/n781 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[55]  ( .D(\fpu_add_frac_dp/n3993 ), .CLK(n1492), .Q(n196) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[54]  ( .D(\fpu_add_frac_dp/n3994 ), .CLK(n1492), .Q(n227) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[53]  ( .D(\fpu_add_frac_dp/n3995 ), .CLK(n1492), .Q(n228) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[52]  ( .D(\fpu_add_frac_dp/n3996 ), .CLK(n1492), .Q(n229) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[51]  ( .D(\fpu_add_frac_dp/n3997 ), .CLK(n1492), .Q(n230) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[50]  ( .D(\fpu_add_frac_dp/n3998 ), .CLK(n1492), .Q(n231) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[49]  ( .D(\fpu_add_frac_dp/n3999 ), .CLK(n1491), .Q(n232) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[48]  ( .D(\fpu_add_frac_dp/n4000 ), .CLK(n1491), .Q(n233) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[47]  ( .D(\fpu_add_frac_dp/n4001 ), .CLK(n1491), .Q(n197) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[46]  ( .D(\fpu_add_frac_dp/n4002 ), .CLK(n1491), .Q(n198) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[45]  ( .D(\fpu_add_frac_dp/n4003 ), .CLK(n1491), .Q(n234) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[44]  ( .D(\fpu_add_frac_dp/n4004 ), .CLK(n1491), .Q(n235) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[43]  ( .D(\fpu_add_frac_dp/n4005 ), .CLK(n1491), .Q(n236) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[42]  ( .D(\fpu_add_frac_dp/n4006 ), .CLK(n1490), .Q(n199) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[41]  ( .D(\fpu_add_frac_dp/n4007 ), .CLK(n1490), .Q(n237) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[40]  ( .D(\fpu_add_frac_dp/n4008 ), .CLK(n1490), .Q(n259) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[39]  ( .D(\fpu_add_frac_dp/n4009 ), .CLK(n1490), .Q(n200) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[38]  ( .D(\fpu_add_frac_dp/n4010 ), .CLK(n1490), .Q(n238) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[37]  ( .D(\fpu_add_frac_dp/n4011 ), .CLK(n1490), .Q(n201) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[36]  ( .D(\fpu_add_frac_dp/n4012 ), .CLK(n1490), .Q(n239) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[35]  ( .D(\fpu_add_frac_dp/n4013 ), .CLK(n1489), .Q(n202) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[34]  ( .D(\fpu_add_frac_dp/n4014 ), .CLK(n1489), .Q(n240) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[33]  ( .D(\fpu_add_frac_dp/n4015 ), .CLK(n1489), .Q(n241) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[32]  ( .D(\fpu_add_frac_dp/n4016 ), .CLK(n1489), .Q(n242) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[31]  ( .D(\fpu_add_frac_dp/n4017 ), .CLK(n1489), .Q(n243) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[30]  ( .D(\fpu_add_frac_dp/n4018 ), .CLK(n1489), .Q(n203) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[29]  ( .D(\fpu_add_frac_dp/n4019 ), .CLK(n1489), .Q(n244) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[28]  ( .D(\fpu_add_frac_dp/n4020 ), .CLK(n1488), .Q(n245) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[27]  ( .D(\fpu_add_frac_dp/n4021 ), .CLK(n1488), .Q(n204) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[26]  ( .D(\fpu_add_frac_dp/n4022 ), .CLK(n1488), .Q(n246) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[25]  ( .D(\fpu_add_frac_dp/n4023 ), .CLK(n1488), .Q(n247) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[24]  ( .D(\fpu_add_frac_dp/n4024 ), .CLK(n1488), .Q(n248) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[23]  ( .D(\fpu_add_frac_dp/n4025 ), .CLK(n1488), .Q(n318), .QN(\fpu_add_frac_dp/n814 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[22]  ( .D(\fpu_add_frac_dp/n4026 ), .CLK(n1488), .Q(n279), .QN(\fpu_add_frac_dp/n815 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[21]  ( .D(\fpu_add_frac_dp/n4027 ), .CLK(n1487), .Q(n267), .QN(\fpu_add_frac_dp/n816 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[20]  ( .D(\fpu_add_frac_dp/n4028 ), .CLK(n1487), .Q(n263), .QN(\fpu_add_frac_dp/n817 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[19]  ( .D(\fpu_add_frac_dp/n4029 ), .CLK(n1487), .Q(n249) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[18]  ( .D(\fpu_add_frac_dp/n4030 ), .CLK(n1487), .Q(n250) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[17]  ( .D(\fpu_add_frac_dp/n4031 ), .CLK(n1487), .Q(n251) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[16]  ( .D(\fpu_add_frac_dp/n4032 ), .CLK(n1497), .Q(n179) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[15]  ( .D(\fpu_add_frac_dp/n4033 ), .CLK(n1548), .Q(n268), .QN(\fpu_add_frac_dp/n822 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[14]  ( .D(\fpu_add_frac_dp/n4034 ), .CLK(n1547), .Q(n180), .QN(\fpu_add_frac_dp/n823 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[13]  ( .D(\fpu_add_frac_dp/n4035 ), .CLK(n1547), .Q(n327), .QN(\fpu_add_frac_dp/n824 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[12]  ( .D(\fpu_add_frac_dp/n4036 ), .CLK(n1547), .Q(n252) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[11]  ( .D(\fpu_add_frac_dp/n4037 ), .CLK(n1547), .Q(n253) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[10]  ( .D(\fpu_add_frac_dp/n4038 ), .CLK(n1547), .Q(n260) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[9]  ( .D(\fpu_add_frac_dp/n4039 ), 
        .CLK(n1547), .Q(n261) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[8]  ( .D(\fpu_add_frac_dp/n4040 ), 
        .CLK(n1547), .Q(n224) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[7]  ( .D(\fpu_add_frac_dp/n4041 ), 
        .CLK(n1546), .Q(n222) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[6]  ( .D(\fpu_add_frac_dp/n4042 ), 
        .CLK(n1546), .Q(n225) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[5]  ( .D(\fpu_add_frac_dp/n4043 ), 
        .CLK(n1546), .Q(n223) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[4]  ( .D(\fpu_add_frac_dp/n4044 ), 
        .CLK(n1546), .Q(n288), .QN(\fpu_add_frac_dp/n833 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[3]  ( .D(\fpu_add_frac_dp/n4045 ), 
        .CLK(n1546), .Q(n310), .QN(\fpu_add_frac_dp/n834 ) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[2]  ( .D(\fpu_add_frac_dp/n4046 ), 
        .CLK(n1546), .Q(n220) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[1]  ( .D(\fpu_add_frac_dp/n4047 ), 
        .CLK(n1546), .Q(n625) );
  DFFX1 \fpu_add_frac_dp/i_a2stg_frac1/q_reg[0]  ( .D(\fpu_add_frac_dp/n4048 ), 
        .CLK(n1545), .Q(n307), .QN(\fpu_add_frac_dp/n2477 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[54]  ( .D(\fpu_add_frac_dp/n4049 ), 
        .CLK(n1518), .Q(n1130), .QN(\fpu_add_frac_dp/n2364 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[53]  ( .D(\fpu_add_frac_dp/n4050 ), 
        .CLK(n1507), .Q(n650), .QN(\fpu_add_frac_dp/n2442 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[52]  ( .D(\fpu_add_frac_dp/n4051 ), 
        .CLK(n1507), .Q(\fpu_add_frac_dp/n5644 ), .QN(n1304) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[51]  ( .D(\fpu_add_frac_dp/n4052 ), 
        .CLK(n1507), .Q(\fpu_add_frac_dp/n2491 ), .QN(n1089) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[50]  ( .D(\fpu_add_frac_dp/n4053 ), 
        .CLK(n1507), .Q(n427), .QN(\fpu_add_frac_dp/n2535 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[49]  ( .D(\fpu_add_frac_dp/n4054 ), 
        .CLK(n1507), .Q(n1065), .QN(\fpu_add_frac_dp/n5625 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[48]  ( .D(\fpu_add_frac_dp/n4055 ), 
        .CLK(n1507), .Q(n1211), .QN(\fpu_add_frac_dp/n5626 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[47]  ( .D(\fpu_add_frac_dp/n4056 ), 
        .CLK(n1507), .Q(\fpu_add_frac_dp/n5624 ), .QN(\fpu_add_frac_dp/n1123 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[46]  ( .D(\fpu_add_frac_dp/n4057 ), 
        .CLK(n1507), .Q(\fpu_add_frac_dp/n5611 ), .QN(\fpu_add_frac_dp/n1122 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[45]  ( .D(\fpu_add_frac_dp/n4058 ), 
        .CLK(n1507), .Q(n1208), .QN(\fpu_add_frac_dp/n2538 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[44]  ( .D(\fpu_add_frac_dp/n4059 ), 
        .CLK(n1507), .Q(\fpu_add_frac_dp/n5621 ), .QN(n578) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[43]  ( .D(\fpu_add_frac_dp/n4060 ), 
        .CLK(n1507), .Q(n763), .QN(\fpu_add_frac_dp/n2543 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[42]  ( .D(\fpu_add_frac_dp/n4061 ), 
        .CLK(n1507), .Q(n1199), .QN(\fpu_add_frac_dp/n839 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[41]  ( .D(\fpu_add_frac_dp/n4062 ), 
        .CLK(n1507), .Q(\fpu_add_frac_dp/n5620 ), .QN(\fpu_add_frac_dp/n1119 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[40]  ( .D(\fpu_add_frac_dp/n4063 ), 
        .CLK(n1506), .Q(n463), .QN(\fpu_add_frac_dp/n2438 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[39]  ( .D(\fpu_add_frac_dp/n4064 ), 
        .CLK(n1506), .Q(n141) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[38]  ( .D(\fpu_add_frac_dp/n4065 ), 
        .CLK(n1506), .Q(\fpu_add_frac_dp/n5613 ), .QN(n306) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[37]  ( .D(\fpu_add_frac_dp/n4066 ), 
        .CLK(n1506), .Q(\fpu_add_frac_dp/n5612 ), .QN(n719) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[36]  ( .D(\fpu_add_frac_dp/n4067 ), 
        .CLK(n1506), .Q(n1207), .QN(\fpu_add_frac_dp/n841 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[35]  ( .D(\fpu_add_frac_dp/n4068 ), 
        .CLK(n1506), .Q(\fpu_add_frac_dp/n5623 ), .QN(\fpu_add_frac_dp/n1115 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[34]  ( .D(\fpu_add_frac_dp/n4069 ), 
        .CLK(n1506), .Q(n916), .QN(\fpu_add_frac_dp/n2365 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[33]  ( .D(\fpu_add_frac_dp/n4070 ), 
        .CLK(n1506), .Q(n326), .QN(\fpu_add_frac_dp/n2532 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[32]  ( .D(\fpu_add_frac_dp/n4071 ), 
        .CLK(n1506), .Q(\fpu_add_frac_dp/n5622 ), .QN(n358) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[31]  ( .D(\fpu_add_frac_dp/n4072 ), 
        .CLK(n1506), .Q(n1194), .QN(\fpu_add_frac_dp/n2441 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[30]  ( .D(\fpu_add_frac_dp/n4073 ), 
        .CLK(n1506), .Q(n132), .QN(\fpu_add_frac_dp/n843 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[29]  ( .D(\fpu_add_frac_dp/n4074 ), 
        .CLK(n1506), .Q(n1132), .QN(\fpu_add_frac_dp/n2514 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[28]  ( .D(\fpu_add_frac_dp/n4075 ), 
        .CLK(n1506), .Q(\fpu_add_frac_dp/n5605 ), .QN(n428) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[27]  ( .D(\fpu_add_frac_dp/n4076 ), 
        .CLK(n1506), .Q(\fpu_add_frac_dp/n5608 ), .QN(\fpu_add_frac_dp/n1109 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[26]  ( .D(\fpu_add_frac_dp/n4077 ), 
        .CLK(n1505), .Q(\fpu_add_frac_dp/n2482 ), .QN(n1303) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[25]  ( .D(\fpu_add_frac_dp/n4078 ), 
        .CLK(n1505), .Q(\fpu_add_frac_dp/n2486 ), .QN(\fpu_add_frac_dp/n1107 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[24]  ( .D(\fpu_add_frac_dp/n4079 ), 
        .CLK(n1505), .Q(n1127), .QN(\fpu_add_frac_dp/n844 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[23]  ( .D(\fpu_add_frac_dp/n4080 ), 
        .CLK(n1505), .Q(\fpu_add_frac_dp/n2458 ), .QN(\fpu_add_frac_dp/n1106 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[22]  ( .D(\fpu_add_frac_dp/n4081 ), 
        .CLK(n1505), .Q(\fpu_add_frac_dp/n2492 ), .QN(\fpu_add_frac_dp/n1105 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[21]  ( .D(\fpu_add_frac_dp/n4082 ), 
        .CLK(n1505), .Q(n335), .QN(\fpu_add_frac_dp/n845 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[20]  ( .D(\fpu_add_frac_dp/n4083 ), 
        .CLK(n1505), .Q(\fpu_add_frac_dp/n2487 ), .QN(\fpu_add_frac_dp/n1104 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[19]  ( .D(\fpu_add_frac_dp/n4084 ), 
        .CLK(n1505), .Q(\fpu_add_frac_dp/n2485 ), .QN(\fpu_add_frac_dp/n1103 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[18]  ( .D(\fpu_add_frac_dp/n4085 ), 
        .CLK(n1505), .Q(n1192), .QN(\fpu_add_frac_dp/n846 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[17]  ( .D(\fpu_add_frac_dp/n4086 ), 
        .CLK(n1505), .Q(n1131), .QN(\fpu_add_frac_dp/n2536 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[16]  ( .D(\fpu_add_frac_dp/n4087 ), 
        .CLK(n1505), .Q(n1193), .QN(\fpu_add_frac_dp/n5629 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[15]  ( .D(\fpu_add_frac_dp/n4088 ), 
        .CLK(n1505), .Q(n1203), .QN(\fpu_add_frac_dp/n847 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[14]  ( .D(\fpu_add_frac_dp/n4089 ), 
        .CLK(n1505), .Q(n1007), .QN(\fpu_add_frac_dp/n5627 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[13]  ( .D(\fpu_add_frac_dp/n4090 ), 
        .CLK(n1505), .Q(n330) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[12]  ( .D(\fpu_add_frac_dp/n4091 ), 
        .CLK(n1504), .Q(n670), .QN(\fpu_add_frac_dp/n848 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[11]  ( .D(\fpu_add_frac_dp/n4092 ), 
        .CLK(n1504), .Q(\fpu_add_frac_dp/n2457 ), .QN(n357) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[10]  ( .D(\fpu_add_frac_dp/n4093 ), 
        .CLK(n1504), .Q(\fpu_add_frac_dp/n2483 ), .QN(n1088) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[9]  ( .D(\fpu_add_frac_dp/n4094 ), 
        .CLK(n1504), .Q(n697), .QN(\fpu_add_frac_dp/n2374 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[8]  ( .D(\fpu_add_frac_dp/n4095 ), 
        .CLK(n1504), .Q(\fpu_add_frac_dp/n2472 ), .QN(\fpu_add_frac_dp/n1096 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[7]  ( .D(\fpu_add_frac_dp/n4096 ), 
        .CLK(n1504), .Q(\fpu_add_frac_dp/n2489 ), .QN(\fpu_add_frac_dp/n1095 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[6]  ( .D(\fpu_add_frac_dp/n4097 ), 
        .CLK(n1504), .Q(\fpu_add_frac_dp/n2490 ), .QN(\fpu_add_frac_dp/n1094 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[5]  ( .D(\fpu_add_frac_dp/n4098 ), 
        .CLK(n1504), .Q(\fpu_add_frac_dp/n2459 ), .QN(\fpu_add_frac_dp/n1093 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[4]  ( .D(\fpu_add_frac_dp/n4099 ), 
        .CLK(n1504), .Q(n900), .QN(\fpu_add_frac_dp/n2366 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[3]  ( .D(\fpu_add_frac_dp/n4100 ), 
        .CLK(n1504), .Q(n1205), .QN(\fpu_add_frac_dp/n2533 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[2]  ( .D(\fpu_add_frac_dp/n4101 ), 
        .CLK(n1504), .Q(n337), .QN(\fpu_add_frac_dp/n2436 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[1]  ( .D(\fpu_add_frac_dp/n4102 ), 
        .CLK(n1504), .Q(\fpu_add_frac_dp/n2455 ), .QN(\fpu_add_frac_dp/n1090 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2a/q_reg[0]  ( .D(\fpu_add_frac_dp/n4103 ), 
        .CLK(n1504), .Q(n702), .QN(\fpu_add_frac_dp/n851 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[63]  ( .D(\fpu_add_frac_dp/n4104 ), 
        .CLK(n1504), .Q(n1080) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[62]  ( .D(\fpu_add_frac_dp/n4105 ), 
        .CLK(n1503), .Q(\fpu_add_frac_dp/n2469 ), .QN(\fpu_add_frac_dp/n1089 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[61]  ( .D(\fpu_add_frac_dp/n4106 ), 
        .CLK(n1503), .Q(\fpu_add_frac_dp/n2468 ), .QN(\fpu_add_frac_dp/n1088 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[60]  ( .D(\fpu_add_frac_dp/n4107 ), 
        .CLK(n1503), .Q(\fpu_add_frac_dp/n2475 ), .QN(\fpu_add_frac_dp/n1087 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[59]  ( .D(\fpu_add_frac_dp/n4108 ), 
        .CLK(n1503), .Q(\fpu_add_frac_dp/n2467 ), .QN(\fpu_add_frac_dp/n1086 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[58]  ( .D(\fpu_add_frac_dp/n4109 ), 
        .CLK(n1503), .Q(\fpu_add_frac_dp/n2474 ), .QN(\fpu_add_frac_dp/n1085 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[57]  ( .D(\fpu_add_frac_dp/n4110 ), 
        .CLK(n1503), .Q(\fpu_add_frac_dp/n2466 ), .QN(\fpu_add_frac_dp/n1084 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[56]  ( .D(\fpu_add_frac_dp/n4111 ), 
        .CLK(n1503), .Q(\fpu_add_frac_dp/n2473 ), .QN(\fpu_add_frac_dp/n1083 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[55]  ( .D(\fpu_add_frac_dp/n4112 ), 
        .CLK(n1503), .Q(\fpu_add_frac_dp/n2446 ), .QN(\fpu_add_frac_dp/n1082 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[54]  ( .D(\fpu_add_frac_dp/n4113 ), 
        .CLK(n1503), .Q(n593), .QN(\fpu_add_frac_dp/n2340 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[53]  ( .D(\fpu_add_frac_dp/n4114 ), 
        .CLK(n1503), .Q(n592), .QN(\fpu_add_frac_dp/n2285 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[52]  ( .D(\fpu_add_frac_dp/n4115 ), 
        .CLK(n1503), .Q(n591), .QN(\fpu_add_frac_dp/n2309 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[51]  ( .D(\fpu_add_frac_dp/n4116 ), 
        .CLK(n1503), .Q(n169), .QN(\fpu_add_frac_dp/n2398 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[50]  ( .D(\fpu_add_frac_dp/n4117 ), 
        .CLK(n1503), .Q(n165), .QN(\fpu_add_frac_dp/n2396 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[49]  ( .D(\fpu_add_frac_dp/n4118 ), 
        .CLK(n1503), .Q(n78), .QN(\fpu_add_frac_dp/n2376 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[48]  ( .D(\fpu_add_frac_dp/n4119 ), 
        .CLK(n1502), .Q(n589), .QN(\fpu_add_frac_dp/n2334 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[47]  ( .D(\fpu_add_frac_dp/n4120 ), 
        .CLK(n1502), .Q(n588), .QN(\fpu_add_frac_dp/n2379 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[46]  ( .D(\fpu_add_frac_dp/n4121 ), 
        .CLK(n1502), .Q(n587), .QN(\fpu_add_frac_dp/n2280 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[45]  ( .D(\fpu_add_frac_dp/n4122 ), 
        .CLK(n1502), .Q(n164), .QN(\fpu_add_frac_dp/n2310 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[44]  ( .D(\fpu_add_frac_dp/n4123 ), 
        .CLK(n1502), .Q(n163), .QN(\fpu_add_frac_dp/n2278 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[43]  ( .D(\fpu_add_frac_dp/n4124 ), 
        .CLK(n1502), .Q(n29), .QN(\fpu_add_frac_dp/n2316 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[42]  ( .D(\fpu_add_frac_dp/n4125 ), 
        .CLK(n1502), .Q(n28), .QN(\fpu_add_frac_dp/n2279 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[41]  ( .D(\fpu_add_frac_dp/n4126 ), 
        .CLK(n1502), .Q(n27), .QN(\fpu_add_frac_dp/n2423 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[40]  ( .D(\fpu_add_frac_dp/n4127 ), 
        .CLK(n1502), .Q(n167), .QN(\fpu_add_frac_dp/n2381 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[39]  ( .D(\fpu_add_frac_dp/n4128 ), 
        .CLK(n1502), .Q(n77) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[38]  ( .D(\fpu_add_frac_dp/n4129 ), 
        .CLK(n1502), .Q(n76) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[37]  ( .D(\fpu_add_frac_dp/n4130 ), 
        .CLK(n1502), .Q(n26) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[36]  ( .D(\fpu_add_frac_dp/n4131 ), 
        .CLK(n1502), .Q(n25), .QN(\fpu_add_frac_dp/n2388 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[35]  ( .D(\fpu_add_frac_dp/n4132 ), 
        .CLK(n1501), .Q(n24) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[34]  ( .D(\fpu_add_frac_dp/n4133 ), 
        .CLK(n1501), .Q(n9) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[33]  ( .D(\fpu_add_frac_dp/n4134 ), 
        .CLK(n1501), .Q(n8) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[32]  ( .D(\fpu_add_frac_dp/n4135 ), 
        .CLK(n1501), .Q(n7) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[31]  ( .D(\fpu_add_frac_dp/n4136 ), 
        .CLK(n1501), .Q(n114) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[30]  ( .D(\fpu_add_frac_dp/n4137 ), 
        .CLK(n1501), .Q(n113) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[29]  ( .D(\fpu_add_frac_dp/n4138 ), 
        .CLK(n1501), .Q(n112) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[28]  ( .D(\fpu_add_frac_dp/n4139 ), 
        .CLK(n1501), .Q(n639) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[27]  ( .D(\fpu_add_frac_dp/n4140 ), 
        .CLK(n1501), .Q(n277) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[26]  ( .D(\fpu_add_frac_dp/n4141 ), 
        .CLK(n1501), .Q(n637) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[25]  ( .D(\fpu_add_frac_dp/n4142 ), 
        .CLK(n1501), .Q(n276) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[24]  ( .D(\fpu_add_frac_dp/n4143 ), 
        .CLK(n1501), .Q(n636) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[23]  ( .D(\fpu_add_frac_dp/n4144 ), 
        .CLK(n1501), .Q(n275) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[22]  ( .D(\fpu_add_frac_dp/n4145 ), 
        .CLK(n1501), .Q(n635) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[21]  ( .D(\fpu_add_frac_dp/n4146 ), 
        .CLK(n1500), .Q(n274) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[20]  ( .D(\fpu_add_frac_dp/n4147 ), 
        .CLK(n1500), .Q(n634) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[19]  ( .D(\fpu_add_frac_dp/n4148 ), 
        .CLK(n1500), .Q(n273) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[18]  ( .D(\fpu_add_frac_dp/n4149 ), 
        .CLK(n1500), .Q(n633) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[17]  ( .D(\fpu_add_frac_dp/n4150 ), 
        .CLK(n1500), .Q(n272) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[16]  ( .D(\fpu_add_frac_dp/n4151 ), 
        .CLK(n1500), .Q(n122) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[15]  ( .D(\fpu_add_frac_dp/n4152 ), 
        .CLK(n1500), .Q(n53) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[14]  ( .D(\fpu_add_frac_dp/n4153 ), 
        .CLK(n1500), .Q(n121) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[13]  ( .D(\fpu_add_frac_dp/n4154 ), 
        .CLK(n1500), .Q(n52) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[12]  ( .D(\fpu_add_frac_dp/n4155 ), 
        .CLK(n1500), .Q(n120) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[11]  ( .D(\fpu_add_frac_dp/n4156 ), 
        .CLK(n1500), .Q(n39) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[10]  ( .D(\fpu_add_frac_dp/n4157 ), 
        .CLK(n1500), .Q(n81) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[9]  ( .D(\fpu_add_frac_dp/n4158 ), 
        .CLK(n1500), .Q(n32) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[8]  ( .D(\fpu_add_frac_dp/n4159 ), 
        .CLK(n1500), .Q(n80) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[7]  ( .D(\fpu_add_frac_dp/n4160 ), 
        .CLK(n1499), .Q(n31) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[6]  ( .D(\fpu_add_frac_dp/n4161 ), 
        .CLK(n1499), .Q(n79) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[5]  ( .D(\fpu_add_frac_dp/n4162 ), 
        .CLK(n1499), .Q(n30) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[4]  ( .D(\fpu_add_frac_dp/n4163 ), 
        .CLK(n1499), .Q(n11) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[3]  ( .D(\fpu_add_frac_dp/n4164 ), 
        .CLK(n1499), .Q(\fpu_add_frac_dp/a1stg_in2[3] ), .QN(
        \fpu_add_frac_dp/n895 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[2]  ( .D(\fpu_add_frac_dp/n4165 ), 
        .CLK(n1499), .Q(n10) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[1]  ( .D(\fpu_add_frac_dp/n4166 ), 
        .CLK(n1499), .Q(n170) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in2/q_reg[0]  ( .D(\fpu_add_frac_dp/n4167 ), 
        .CLK(n1499), .Q(n36), .QN(\fpu_add_frac_dp/n898 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[54]  ( .D(\fpu_add_frac_dp/n4168 ), 
        .CLK(n1499), .Q(n283) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[53]  ( .D(\fpu_add_frac_dp/n4169 ), 
        .CLK(n1499), .Q(n747), .QN(\fpu_add_frac_dp/n900 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[52]  ( .D(\fpu_add_frac_dp/n4170 ), 
        .CLK(n1499), .Q(n548), .QN(\fpu_add_frac_dp/n5643 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[51]  ( .D(\fpu_add_frac_dp/n4171 ), 
        .CLK(n1499), .Q(n340), .QN(\fpu_add_frac_dp/n901 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[50]  ( .D(\fpu_add_frac_dp/n4172 ), 
        .CLK(n1499), .Q(\fpu_add_frac_dp/n2350 ), .QN(n1158) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[49]  ( .D(\fpu_add_frac_dp/n4173 ), 
        .CLK(n1499), .Q(n917), .QN(\fpu_add_frac_dp/n2415 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[48]  ( .D(\fpu_add_frac_dp/n4174 ), 
        .CLK(n1498), .Q(\fpu_add_frac_dp/n2476 ), .QN(\fpu_add_frac_dp/n1070 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[47]  ( .D(\fpu_add_frac_dp/n4175 ), 
        .CLK(n1498), .Q(n1202), .QN(\fpu_add_frac_dp/n903 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[46]  ( .D(\fpu_add_frac_dp/n4176 ), 
        .CLK(n1498), .Q(n1198), .QN(\fpu_add_frac_dp/n904 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[45]  ( .D(\fpu_add_frac_dp/n4177 ), 
        .CLK(n1498), .Q(n677), .QN(\fpu_add_frac_dp/n2373 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[44]  ( .D(\fpu_add_frac_dp/n4178 ), 
        .CLK(n1498), .Q(n57), .QN(\fpu_add_frac_dp/n905 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[43]  ( .D(\fpu_add_frac_dp/n4179 ), 
        .CLK(n1498), .Q(n848), .QN(\fpu_add_frac_dp/n2540 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[42]  ( .D(\fpu_add_frac_dp/n4180 ), 
        .CLK(n1498), .Q(\fpu_add_frac_dp/n2462 ), .QN(\fpu_add_frac_dp/n1067 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[41]  ( .D(\fpu_add_frac_dp/n4181 ), 
        .CLK(n1498), .Q(n1129), .QN(\fpu_add_frac_dp/n907 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[40]  ( .D(\fpu_add_frac_dp/n4182 ), 
        .CLK(n1498), .Q(n709), .QN(\fpu_add_frac_dp/n908 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[39]  ( .D(\fpu_add_frac_dp/n4183 ), 
        .CLK(n1498), .Q(\fpu_add_frac_dp/n2452 ), .QN(n1079) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[38]  ( .D(\fpu_add_frac_dp/n4184 ), 
        .CLK(n1498), .Q(n46) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[37]  ( .D(\fpu_add_frac_dp/n4185 ), 
        .CLK(n1498), .Q(n125) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[36]  ( .D(\fpu_add_frac_dp/n4186 ), 
        .CLK(n1498), .Q(n292), .QN(\fpu_add_frac_dp/n2408 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[35]  ( .D(\fpu_add_frac_dp/n4187 ), 
        .CLK(n1498), .Q(n1215), .QN(\fpu_add_frac_dp/n911 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[34]  ( .D(\fpu_add_frac_dp/n4188 ), 
        .CLK(n1497), .Q(n857), .QN(\fpu_add_frac_dp/n912 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[33]  ( .D(\fpu_add_frac_dp/n4189 ), 
        .CLK(n1497), .Q(\fpu_add_frac_dp/n2295 ), .QN(n1067) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[32]  ( .D(\fpu_add_frac_dp/n4190 ), 
        .CLK(n1497), .Q(n855), .QN(\fpu_add_frac_dp/n913 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[31]  ( .D(\fpu_add_frac_dp/n4191 ), 
        .CLK(n1497), .Q(n704) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[30]  ( .D(\fpu_add_frac_dp/n4192 ), 
        .CLK(n1497), .Q(\fpu_add_frac_dp/n2445 ), .QN(n989) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[29]  ( .D(\fpu_add_frac_dp/n4193 ), 
        .CLK(n1497), .Q(n856), .QN(\fpu_add_frac_dp/n2367 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[28]  ( .D(\fpu_add_frac_dp/n4194 ), 
        .CLK(n1497), .Q(n54) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[27]  ( .D(\fpu_add_frac_dp/n4195 ), 
        .CLK(n1497), .Q(n647) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[26]  ( .D(\fpu_add_frac_dp/n4196 ), 
        .CLK(n1497), .Q(n550), .QN(\fpu_add_frac_dp/n917 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[25]  ( .D(\fpu_add_frac_dp/n4197 ), 
        .CLK(n1497), .Q(n1209), .QN(\fpu_add_frac_dp/n918 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[24]  ( .D(\fpu_add_frac_dp/n4198 ), 
        .CLK(n1497), .Q(\fpu_add_frac_dp/n2488 ), .QN(\fpu_add_frac_dp/n1056 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[23]  ( .D(\fpu_add_frac_dp/n4199 ), 
        .CLK(n1497), .Q(n1206), .QN(\fpu_add_frac_dp/n919 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[22]  ( .D(\fpu_add_frac_dp/n4200 ), 
        .CLK(n1497), .Q(n1204), .QN(\fpu_add_frac_dp/n920 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[21]  ( .D(\fpu_add_frac_dp/n4201 ), 
        .CLK(n1502), .Q(\fpu_add_frac_dp/n2444 ), .QN(n1078) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[20]  ( .D(\fpu_add_frac_dp/n4202 ), 
        .CLK(n1518), .Q(n1143), .QN(\fpu_add_frac_dp/n921 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[19]  ( .D(\fpu_add_frac_dp/n4203 ), 
        .CLK(n1518), .Q(n1197), .QN(\fpu_add_frac_dp/n922 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[18]  ( .D(\fpu_add_frac_dp/n4204 ), 
        .CLK(n1518), .Q(n1153), .QN(\fpu_add_frac_dp/n2439 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[17]  ( .D(\fpu_add_frac_dp/n4205 ), 
        .CLK(n1518), .Q(n853), .QN(\fpu_add_frac_dp/n2372 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[16]  ( .D(\fpu_add_frac_dp/n4206 ), 
        .CLK(n1518), .Q(n703), .QN(\fpu_add_frac_dp/n2305 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[15]  ( .D(\fpu_add_frac_dp/n4207 ), 
        .CLK(n1518), .Q(\fpu_add_frac_dp/n2453 ), .QN(\fpu_add_frac_dp/n1050 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[14]  ( .D(\fpu_add_frac_dp/n4208 ), 
        .CLK(n1518), .Q(n988), .QN(\fpu_add_frac_dp/n2454 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[13]  ( .D(\fpu_add_frac_dp/n4209 ), 
        .CLK(n1518), .Q(n1184), .QN(\fpu_add_frac_dp/n2368 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[12]  ( .D(\fpu_add_frac_dp/n4210 ), 
        .CLK(n1518), .Q(\fpu_add_frac_dp/n2484 ), .QN(\fpu_add_frac_dp/n1048 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[11]  ( .D(\fpu_add_frac_dp/n4211 ), 
        .CLK(n1518), .Q(n854), .QN(\fpu_add_frac_dp/n927 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[10]  ( .D(\fpu_add_frac_dp/n4212 ), 
        .CLK(n1517), .Q(n145), .QN(\fpu_add_frac_dp/n928 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[9]  ( .D(\fpu_add_frac_dp/n4213 ), 
        .CLK(n1517), .Q(n577), .QN(\fpu_add_frac_dp/n2544 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[8]  ( .D(\fpu_add_frac_dp/n4214 ), 
        .CLK(n1517), .Q(n1146), .QN(\fpu_add_frac_dp/n929 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[7]  ( .D(\fpu_add_frac_dp/n4215 ), 
        .CLK(n1517), .Q(n1195), .QN(\fpu_add_frac_dp/n930 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[6]  ( .D(\fpu_add_frac_dp/n4216 ), 
        .CLK(n1517), .Q(n1133), .QN(\fpu_add_frac_dp/n931 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[5]  ( .D(\fpu_add_frac_dp/n4217 ), 
        .CLK(n1517), .Q(n1128), .QN(\fpu_add_frac_dp/n932 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[4]  ( .D(\fpu_add_frac_dp/n4218 ), 
        .CLK(n1517), .Q(n695), .QN(\fpu_add_frac_dp/n933 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[3]  ( .D(\fpu_add_frac_dp/n4219 ), 
        .CLK(n1517), .Q(\fpu_add_frac_dp/n2296 ), .QN(\fpu_add_frac_dp/n1045 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[2]  ( .D(\fpu_add_frac_dp/n4220 ), 
        .CLK(n1517), .Q(n745), .QN(\fpu_add_frac_dp/n934 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[1]  ( .D(\fpu_add_frac_dp/n4221 ), 
        .CLK(n1517), .Q(n1185), .QN(\fpu_add_frac_dp/n935 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1a/q_reg[0]  ( .D(\fpu_add_frac_dp/n4222 ), 
        .CLK(n1517), .Q(\fpu_add_frac_dp/n2493 ), .QN(\fpu_add_frac_dp/n1044 )
         );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[62]  ( .D(\fpu_add_frac_dp/n4223 ), 
        .CLK(n1517), .Q(n715) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[61]  ( .D(\fpu_add_frac_dp/n4224 ), 
        .CLK(n1517), .Q(n1191), .QN(\fpu_add_frac_dp/n937 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[60]  ( .D(\fpu_add_frac_dp/n4225 ), 
        .CLK(n1517), .Q(n712) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[59]  ( .D(\fpu_add_frac_dp/n4226 ), 
        .CLK(n1516), .Q(n713) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[58]  ( .D(\fpu_add_frac_dp/n4227 ), 
        .CLK(n1516), .Q(n1190), .QN(\fpu_add_frac_dp/n940 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[57]  ( .D(\fpu_add_frac_dp/n4228 ), 
        .CLK(n1516), .Q(n714) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[56]  ( .D(\fpu_add_frac_dp/n4229 ), 
        .CLK(n1516), .Q(n1189), .QN(\fpu_add_frac_dp/n942 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[55]  ( .D(\fpu_add_frac_dp/n4230 ), 
        .CLK(n1516), .Q(n1188), .QN(\fpu_add_frac_dp/n943 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[54]  ( .D(\fpu_add_frac_dp/n4231 ), 
        .CLK(n1516), .Q(n705), .QN(\fpu_add_frac_dp/n2534 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[53]  ( .D(\fpu_add_frac_dp/n4232 ), 
        .CLK(n1516), .Q(n689), .QN(\fpu_add_frac_dp/n945 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[52]  ( .D(\fpu_add_frac_dp/n4233 ), 
        .CLK(n1516), .Q(n688), .QN(\fpu_add_frac_dp/n2521 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[51]  ( .D(\fpu_add_frac_dp/n4234 ), 
        .CLK(n1516), .Q(n206) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[50]  ( .D(\fpu_add_frac_dp/n4235 ), 
        .CLK(n1516), .Q(n216) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[49]  ( .D(\fpu_add_frac_dp/n4236 ), 
        .CLK(n1516), .Q(n215) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[48]  ( .D(\fpu_add_frac_dp/n4237 ), 
        .CLK(n1516), .Q(n621) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[47]  ( .D(\fpu_add_frac_dp/n4238 ), 
        .CLK(n1516), .Q(n620) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[46]  ( .D(\fpu_add_frac_dp/n4239 ), 
        .CLK(n1516), .Q(n619) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[45]  ( .D(\fpu_add_frac_dp/n4240 ), 
        .CLK(n1515), .Q(n214) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[44]  ( .D(\fpu_add_frac_dp/n4241 ), 
        .CLK(n1515), .Q(n213) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[43]  ( .D(\fpu_add_frac_dp/n4242 ), 
        .CLK(n1515), .Q(n212) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[42]  ( .D(\fpu_add_frac_dp/n4243 ), 
        .CLK(n1515), .Q(n618) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[41]  ( .D(\fpu_add_frac_dp/n4244 ), 
        .CLK(n1515), .Q(n617) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[40]  ( .D(\fpu_add_frac_dp/n4245 ), 
        .CLK(n1515), .Q(n616) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[39]  ( .D(\fpu_add_frac_dp/n4246 ), 
        .CLK(n1515), .Q(n211) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[38]  ( .D(\fpu_add_frac_dp/n4247 ), 
        .CLK(n1515), .Q(n210) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[37]  ( .D(\fpu_add_frac_dp/n4248 ), 
        .CLK(n1515), .Q(n209) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[36]  ( .D(\fpu_add_frac_dp/n4249 ), 
        .CLK(n1515), .Q(n615) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[35]  ( .D(\fpu_add_frac_dp/n4250 ), 
        .CLK(n1515), .Q(n614) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[34]  ( .D(\fpu_add_frac_dp/n4251 ), 
        .CLK(n1515), .Q(n99) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[33]  ( .D(\fpu_add_frac_dp/n4252 ), 
        .CLK(n1515), .Q(n208) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[32]  ( .D(\fpu_add_frac_dp/n4253 ), 
        .CLK(n1515), .Q(n176), .QN(\fpu_add_frac_dp/n965 ) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[31]  ( .D(\fpu_add_frac_dp/n4254 ), 
        .CLK(n1514), .Q(n699) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[30]  ( .D(\fpu_add_frac_dp/n4255 ), 
        .CLK(n1514), .Q(n698) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[29]  ( .D(\fpu_add_frac_dp/n4256 ), 
        .CLK(n1514), .Q(n644) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[28]  ( .D(\fpu_add_frac_dp/n4257 ), 
        .CLK(n1514), .Q(n207) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[27]  ( .D(\fpu_add_frac_dp/n4258 ), 
        .CLK(n1514), .Q(n611) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[26]  ( .D(\fpu_add_frac_dp/n4259 ), 
        .CLK(n1514), .Q(n194) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[25]  ( .D(\fpu_add_frac_dp/n4260 ), 
        .CLK(n1514), .Q(n610) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[24]  ( .D(\fpu_add_frac_dp/n4261 ), 
        .CLK(n1514), .Q(n193) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[23]  ( .D(\fpu_add_frac_dp/n4262 ), 
        .CLK(n1514), .Q(n609) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[22]  ( .D(\fpu_add_frac_dp/n4263 ), 
        .CLK(n1514), .Q(n192) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[21]  ( .D(\fpu_add_frac_dp/n4264 ), 
        .CLK(n1514), .Q(n608) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[20]  ( .D(\fpu_add_frac_dp/n4265 ), 
        .CLK(n1514), .Q(n191) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[19]  ( .D(\fpu_add_frac_dp/n4266 ), 
        .CLK(n1514), .Q(n607) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[18]  ( .D(\fpu_add_frac_dp/n4267 ), 
        .CLK(n1514), .Q(n190) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[17]  ( .D(\fpu_add_frac_dp/n4268 ), 
        .CLK(n1513), .Q(n606) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[16]  ( .D(\fpu_add_frac_dp/n4269 ), 
        .CLK(n1513), .Q(n189) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[15]  ( .D(\fpu_add_frac_dp/n4270 ), 
        .CLK(n1513), .Q(n605) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[14]  ( .D(\fpu_add_frac_dp/n4271 ), 
        .CLK(n1513), .Q(n188) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[13]  ( .D(\fpu_add_frac_dp/n4272 ), 
        .CLK(n1513), .Q(n604) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[12]  ( .D(\fpu_add_frac_dp/n4273 ), 
        .CLK(n1513), .Q(n187) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[11]  ( .D(\fpu_add_frac_dp/n4274 ), 
        .CLK(n1513), .Q(n603) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[10]  ( .D(\fpu_add_frac_dp/n4275 ), 
        .CLK(n1513), .Q(n186) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[9]  ( .D(\fpu_add_frac_dp/n4276 ), 
        .CLK(n1513), .Q(n602) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[8]  ( .D(\fpu_add_frac_dp/n4277 ), 
        .CLK(n1513), .Q(n185) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[7]  ( .D(\fpu_add_frac_dp/n4278 ), 
        .CLK(n1513), .Q(n601) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[6]  ( .D(\fpu_add_frac_dp/n4279 ), 
        .CLK(n1513), .Q(n184) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[5]  ( .D(\fpu_add_frac_dp/n4280 ), 
        .CLK(n1513), .Q(n600) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[4]  ( .D(\fpu_add_frac_dp/n4281 ), 
        .CLK(n1512), .Q(n183) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[3]  ( .D(\fpu_add_frac_dp/n4282 ), 
        .CLK(n1512), .Q(n599) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[2]  ( .D(\fpu_add_frac_dp/n4283 ), 
        .CLK(n1512), .Q(n182) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[1]  ( .D(\fpu_add_frac_dp/n4284 ), 
        .CLK(n1512), .Q(n93) );
  DFFX1 \fpu_add_frac_dp/i_a1stg_in1/q_reg[0]  ( .D(\fpu_add_frac_dp/n4285 ), 
        .CLK(n1512), .Q(n612) );
  LATCHX1 \fpu_add_frac_dp/ckbuf_add_frac_dp/clken_reg  ( .CLK(
        \fpu_add_frac_dp/n2189 ), .D(\fpu_add_frac_dp/ckbuf_add_frac_dp/N1 ), 
        .Q(\fpu_add_frac_dp/ckbuf_add_frac_dp/clken ), .QN(
        \fpu_add_frac_dp/n998 ) );
  OR2X1 U2 ( .IN1(n4114), .IN2(\fpu_add_ctl/n210 ), .Q(n586) );
  OR2X1 U3 ( .IN1(n2590), .IN2(n1745), .Q(n590) );
  OR2X1 U4 ( .IN1(\fpu_add_frac_dp/n132 ), .IN2(\fpu_add_frac_dp/n134 ), .Q(
        n628) );
  INVX0 U5 ( .INP(\fpu_add_frac_dp/n5617 ), .ZN(n1305) );
  INVX0 U6 ( .INP(\fpu_add_frac_dp/n5617 ), .ZN(n1306) );
  INVX0 U7 ( .INP(\fpu_add_frac_dp/n5617 ), .ZN(n1307) );
  INVX0 U8 ( .INP(\fpu_add_frac_dp/n5616 ), .ZN(n1308) );
  INVX0 U9 ( .INP(\fpu_add_frac_dp/n5616 ), .ZN(n1309) );
  INVX0 U10 ( .INP(\fpu_add_frac_dp/n5616 ), .ZN(n1310) );
  INVX0 U11 ( .INP(n3973), .ZN(n1311) );
  INVX0 U12 ( .INP(n3973), .ZN(n1312) );
  INVX0 U13 ( .INP(n3973), .ZN(n1313) );
  INVX0 U14 ( .INP(n3973), .ZN(n1314) );
  INVX0 U15 ( .INP(n628), .ZN(n1315) );
  INVX0 U16 ( .INP(n628), .ZN(n1316) );
  INVX0 U17 ( .INP(n628), .ZN(n1317) );
  INVX0 U18 ( .INP(n628), .ZN(n1318) );
  INVX0 U19 ( .INP(n590), .ZN(n1319) );
  INVX0 U20 ( .INP(n590), .ZN(n1320) );
  INVX0 U21 ( .INP(n590), .ZN(n1321) );
  INVX0 U22 ( .INP(n590), .ZN(n1322) );
  INVX0 U23 ( .INP(\fpu_add_ctl/n1 ), .ZN(n1323) );
  INVX0 U24 ( .INP(\fpu_add_ctl/n1 ), .ZN(n1324) );
  INVX0 U25 ( .INP(\fpu_add_ctl/n1 ), .ZN(n1325) );
  INVX0 U26 ( .INP(\fpu_add_frac_dp/n5614 ), .ZN(n1326) );
  INVX0 U27 ( .INP(\fpu_add_frac_dp/n5614 ), .ZN(n1327) );
  INVX0 U28 ( .INP(\fpu_add_frac_dp/n5614 ), .ZN(n1328) );
  INVX0 U29 ( .INP(n1933), .ZN(n1329) );
  INVX0 U30 ( .INP(n1933), .ZN(n1330) );
  INVX0 U31 ( .INP(n1933), .ZN(n1331) );
  INVX0 U32 ( .INP(n1933), .ZN(n1332) );
  INVX0 U33 ( .INP(n586), .ZN(n1333) );
  INVX0 U34 ( .INP(n586), .ZN(n1334) );
  INVX0 U35 ( .INP(n586), .ZN(n1335) );
  INVX0 U36 ( .INP(n586), .ZN(n1336) );
  INVX0 U37 ( .INP(n4057), .ZN(n1337) );
  INVX0 U38 ( .INP(n4057), .ZN(n1338) );
  INVX0 U39 ( .INP(n4057), .ZN(n1339) );
  INVX0 U40 ( .INP(n4057), .ZN(n1340) );
  INVX2 U41 ( .INP(n1811), .ZN(n1594) );
  INVX2 U42 ( .INP(n1598), .ZN(n1597) );
  NOR2X1 U43 ( .IN1(n584), .IN2(n1745), .QN(n2994) );
  NOR2X1 U44 ( .IN1(n129), .IN2(n295), .QN(n1596) );
  INVX2 U45 ( .INP(n3071), .ZN(n3065) );
  NAND2X1 U46 ( .IN1(n3156), .IN2(n3157), .QN(\fpu_add_frac_dp/n1509 ) );
  INVX0 U47 ( .INP(n1450), .ZN(n1440) );
  INVX0 U48 ( .INP(n1450), .ZN(n1439) );
  INVX0 U49 ( .INP(n1450), .ZN(n1436) );
  INVX0 U50 ( .INP(n1450), .ZN(n1437) );
  INVX0 U51 ( .INP(n1450), .ZN(n1438) );
  INVX0 U52 ( .INP(n1450), .ZN(n1441) );
  INVX0 U53 ( .INP(n1473), .ZN(n1462) );
  INVX0 U54 ( .INP(n1450), .ZN(n1443) );
  INVX0 U55 ( .INP(n1450), .ZN(n1444) );
  INVX0 U56 ( .INP(n1450), .ZN(n1445) );
  INVX0 U57 ( .INP(n1450), .ZN(n1448) );
  INVX0 U58 ( .INP(n1450), .ZN(n1447) );
  INVX0 U59 ( .INP(n1450), .ZN(n1446) );
  INVX0 U60 ( .INP(n1450), .ZN(n1442) );
  INVX0 U61 ( .INP(n1450), .ZN(n1435) );
  INVX0 U62 ( .INP(n1473), .ZN(n1463) );
  INVX0 U63 ( .INP(n1473), .ZN(n1464) );
  INVX0 U64 ( .INP(n1473), .ZN(n1472) );
  INVX0 U65 ( .INP(n1473), .ZN(n1465) );
  INVX0 U66 ( .INP(n1473), .ZN(n1466) );
  INVX0 U67 ( .INP(n1473), .ZN(n1467) );
  INVX0 U68 ( .INP(n1473), .ZN(n1468) );
  INVX0 U69 ( .INP(n1473), .ZN(n1469) );
  INVX0 U70 ( .INP(n1473), .ZN(n1470) );
  INVX0 U71 ( .INP(n1473), .ZN(n1471) );
  INVX0 U72 ( .INP(n1431), .ZN(n1430) );
  INVX0 U73 ( .INP(n1434), .ZN(n1389) );
  INVX0 U74 ( .INP(n1432), .ZN(n1415) );
  INVX0 U75 ( .INP(n1434), .ZN(n1395) );
  INVX0 U76 ( .INP(n1434), .ZN(n1390) );
  INVX0 U77 ( .INP(n1434), .ZN(n1394) );
  INVX0 U78 ( .INP(n1434), .ZN(n1391) );
  INVX0 U79 ( .INP(n1434), .ZN(n1392) );
  INVX0 U80 ( .INP(n1434), .ZN(n1393) );
  INVX0 U81 ( .INP(n1433), .ZN(n1396) );
  INVX0 U82 ( .INP(n1433), .ZN(n1398) );
  INVX0 U83 ( .INP(n1433), .ZN(n1403) );
  INVX0 U84 ( .INP(n1433), .ZN(n1402) );
  INVX0 U85 ( .INP(n1433), .ZN(n1399) );
  INVX0 U86 ( .INP(n1433), .ZN(n1401) );
  INVX0 U87 ( .INP(n1433), .ZN(n1400) );
  INVX0 U88 ( .INP(n1433), .ZN(n1397) );
  INVX0 U89 ( .INP(n1433), .ZN(n1405) );
  INVX0 U90 ( .INP(n1433), .ZN(n1404) );
  INVX0 U91 ( .INP(n1433), .ZN(n1406) );
  INVX0 U92 ( .INP(n1432), .ZN(n1409) );
  INVX0 U93 ( .INP(n1432), .ZN(n1408) );
  INVX0 U94 ( .INP(n1433), .ZN(n1407) );
  INVX0 U95 ( .INP(n1432), .ZN(n1410) );
  INVX0 U96 ( .INP(n1432), .ZN(n1411) );
  INVX0 U97 ( .INP(n1432), .ZN(n1412) );
  INVX0 U98 ( .INP(n1432), .ZN(n1413) );
  INVX0 U99 ( .INP(n1432), .ZN(n1414) );
  INVX0 U100 ( .INP(n1432), .ZN(n1416) );
  INVX0 U101 ( .INP(n1434), .ZN(n1388) );
  INVX0 U102 ( .INP(n1434), .ZN(n1387) );
  INVX0 U103 ( .INP(n1434), .ZN(n1386) );
  INVX0 U104 ( .INP(n1434), .ZN(n1385) );
  INVX0 U105 ( .INP(n1434), .ZN(n1384) );
  INVX0 U106 ( .INP(n1432), .ZN(n1418) );
  INVX0 U107 ( .INP(n1431), .ZN(n1420) );
  INVX0 U108 ( .INP(n1431), .ZN(n1422) );
  INVX0 U109 ( .INP(n1431), .ZN(n1423) );
  INVX0 U110 ( .INP(n1431), .ZN(n1424) );
  INVX0 U111 ( .INP(n1431), .ZN(n1425) );
  INVX0 U112 ( .INP(n1431), .ZN(n1421) );
  INVX0 U113 ( .INP(n1431), .ZN(n1426) );
  INVX0 U114 ( .INP(n1431), .ZN(n1427) );
  INVX0 U115 ( .INP(n1431), .ZN(n1428) );
  INVX0 U116 ( .INP(n1431), .ZN(n1429) );
  INVX0 U117 ( .INP(n1432), .ZN(n1419) );
  INVX0 U118 ( .INP(n1432), .ZN(n1417) );
  INVX0 U119 ( .INP(n2046), .ZN(n1379) );
  INVX0 U120 ( .INP(n2046), .ZN(n1380) );
  INVX0 U121 ( .INP(n2046), .ZN(n1381) );
  INVX0 U122 ( .INP(n2046), .ZN(n1382) );
  INVX0 U123 ( .INP(n1431), .ZN(n1383) );
  INVX0 U124 ( .INP(n1450), .ZN(n1449) );
  INVX0 U125 ( .INP(n1473), .ZN(n1461) );
  INVX0 U126 ( .INP(n4000), .ZN(n1473) );
  INVX0 U127 ( .INP(n3986), .ZN(n1451) );
  INVX0 U128 ( .INP(n3986), .ZN(n1452) );
  INVX0 U129 ( .INP(n3986), .ZN(n1453) );
  INVX0 U130 ( .INP(n3986), .ZN(n1454) );
  INVX0 U131 ( .INP(n3986), .ZN(n1455) );
  INVX0 U132 ( .INP(n3986), .ZN(n1456) );
  INVX0 U133 ( .INP(n3986), .ZN(n1457) );
  INVX0 U134 ( .INP(n3986), .ZN(n1458) );
  INVX0 U135 ( .INP(n3986), .ZN(n1459) );
  INVX0 U136 ( .INP(n3986), .ZN(n1460) );
  INVX0 U137 ( .INP(n1746), .ZN(n1450) );
  INVX0 U138 ( .INP(n1379), .ZN(n1431) );
  INVX0 U139 ( .INP(n1380), .ZN(n1432) );
  INVX0 U140 ( .INP(n1381), .ZN(n1433) );
  INVX0 U141 ( .INP(n1382), .ZN(n1434) );
  INVX0 U142 ( .INP(n1357), .ZN(n1348) );
  INVX0 U143 ( .INP(n1357), .ZN(n1347) );
  INVX0 U144 ( .INP(n1357), .ZN(n1345) );
  INVX0 U145 ( .INP(n1357), .ZN(n1344) );
  INVX0 U146 ( .INP(n1357), .ZN(n1346) );
  INVX0 U147 ( .INP(n1357), .ZN(n1349) );
  INVX0 U148 ( .INP(n1357), .ZN(n1352) );
  INVX0 U149 ( .INP(n1357), .ZN(n1351) );
  INVX0 U150 ( .INP(n1357), .ZN(n1350) );
  INVX0 U151 ( .INP(n1357), .ZN(n1353) );
  INVX0 U152 ( .INP(n1357), .ZN(n1354) );
  INVX0 U153 ( .INP(n1357), .ZN(n1356) );
  INVX0 U154 ( .INP(n1357), .ZN(n1355) );
  INVX0 U155 ( .INP(n1357), .ZN(n1343) );
  INVX0 U156 ( .INP(n1377), .ZN(n1375) );
  INVX0 U157 ( .INP(n1377), .ZN(n1374) );
  INVX0 U158 ( .INP(n1377), .ZN(n1373) );
  INVX0 U159 ( .INP(n1377), .ZN(n1372) );
  INVX0 U160 ( .INP(n1377), .ZN(n1371) );
  INVX0 U161 ( .INP(n1377), .ZN(n1370) );
  INVX0 U162 ( .INP(n1377), .ZN(n1369) );
  INVX0 U163 ( .INP(n1377), .ZN(n1368) );
  INVX0 U164 ( .INP(n1377), .ZN(n1367) );
  INVX0 U165 ( .INP(n1377), .ZN(n1366) );
  INVX0 U166 ( .INP(n1378), .ZN(n1365) );
  INVX0 U167 ( .INP(n1378), .ZN(n1364) );
  INVX0 U168 ( .INP(n1378), .ZN(n1363) );
  INVX0 U169 ( .INP(n1378), .ZN(n1362) );
  INVX0 U170 ( .INP(n1378), .ZN(n1361) );
  INVX0 U171 ( .INP(n1378), .ZN(n1360) );
  INVX0 U172 ( .INP(n1378), .ZN(n1359) );
  INVX0 U173 ( .INP(n1378), .ZN(n1358) );
  INVX0 U174 ( .INP(n1561), .ZN(n1514) );
  INVX0 U175 ( .INP(n1561), .ZN(n1515) );
  INVX0 U176 ( .INP(n1561), .ZN(n1516) );
  INVX0 U177 ( .INP(n1561), .ZN(n1517) );
  INVX0 U178 ( .INP(n1562), .ZN(n1498) );
  INVX0 U179 ( .INP(n1562), .ZN(n1499) );
  INVX0 U180 ( .INP(n1562), .ZN(n1500) );
  INVX0 U181 ( .INP(n1562), .ZN(n1501) );
  INVX0 U182 ( .INP(n1562), .ZN(n1502) );
  INVX0 U183 ( .INP(n1562), .ZN(n1503) );
  INVX0 U184 ( .INP(n1562), .ZN(n1504) );
  INVX0 U185 ( .INP(n1562), .ZN(n1505) );
  INVX0 U186 ( .INP(n1562), .ZN(n1506) );
  INVX0 U187 ( .INP(n1563), .ZN(n1497) );
  INVX0 U188 ( .INP(n1563), .ZN(n1494) );
  INVX0 U189 ( .INP(n1563), .ZN(n1495) );
  INVX0 U190 ( .INP(n1563), .ZN(n1496) );
  INVX0 U191 ( .INP(n1564), .ZN(n1482) );
  INVX0 U192 ( .INP(n1564), .ZN(n1483) );
  INVX0 U193 ( .INP(n1564), .ZN(n1484) );
  INVX0 U194 ( .INP(n1564), .ZN(n1485) );
  INVX0 U195 ( .INP(n1558), .ZN(n1546) );
  INVX0 U196 ( .INP(n1558), .ZN(n1547) );
  INVX0 U197 ( .INP(n1563), .ZN(n1488) );
  INVX0 U198 ( .INP(n1563), .ZN(n1489) );
  INVX0 U199 ( .INP(n1563), .ZN(n1490) );
  INVX0 U200 ( .INP(n1563), .ZN(n1491) );
  INVX0 U201 ( .INP(n1563), .ZN(n1492) );
  INVX0 U202 ( .INP(n1563), .ZN(n1493) );
  INVX0 U203 ( .INP(n1558), .ZN(n1554) );
  INVX0 U204 ( .INP(n1558), .ZN(n1553) );
  INVX0 U205 ( .INP(n1563), .ZN(n1486) );
  INVX0 U206 ( .INP(n1564), .ZN(n1480) );
  INVX0 U207 ( .INP(n1563), .ZN(n1487) );
  INVX0 U208 ( .INP(n1561), .ZN(n1513) );
  INVX0 U209 ( .INP(n1562), .ZN(n1507) );
  INVX0 U210 ( .INP(n1562), .ZN(n1508) );
  INVX0 U211 ( .INP(n1562), .ZN(n1509) );
  INVX0 U212 ( .INP(n1561), .ZN(n1511) );
  INVX0 U213 ( .INP(n1561), .ZN(n1512) );
  INVX0 U214 ( .INP(n1561), .ZN(n1510) );
  INVX0 U215 ( .INP(n1559), .ZN(n1544) );
  INVX0 U216 ( .INP(n1559), .ZN(n1542) );
  INVX0 U217 ( .INP(n1559), .ZN(n1545) );
  INVX0 U218 ( .INP(n1558), .ZN(n1556) );
  INVX0 U219 ( .INP(n1559), .ZN(n1543) );
  INVX0 U220 ( .INP(n1559), .ZN(n1539) );
  INVX0 U221 ( .INP(n1559), .ZN(n1540) );
  INVX0 U222 ( .INP(n1559), .ZN(n1541) );
  INVX0 U223 ( .INP(n1560), .ZN(n1527) );
  INVX0 U224 ( .INP(n1558), .ZN(n1552) );
  INVX0 U225 ( .INP(n1558), .ZN(n1548) );
  INVX0 U226 ( .INP(n1558), .ZN(n1549) );
  INVX0 U227 ( .INP(n1558), .ZN(n1550) );
  INVX0 U228 ( .INP(n1558), .ZN(n1551) );
  INVX0 U229 ( .INP(n1559), .ZN(n1534) );
  INVX0 U230 ( .INP(n1564), .ZN(n1481) );
  INVX0 U231 ( .INP(n1558), .ZN(n1555) );
  INVX0 U232 ( .INP(n1560), .ZN(n1533) );
  INVX0 U233 ( .INP(n1559), .ZN(n1535) );
  INVX0 U234 ( .INP(n1560), .ZN(n1532) );
  INVX0 U235 ( .INP(n1561), .ZN(n1519) );
  INVX0 U236 ( .INP(n1561), .ZN(n1518) );
  INVX0 U237 ( .INP(n1559), .ZN(n1538) );
  INVX0 U238 ( .INP(n1559), .ZN(n1537) );
  INVX0 U239 ( .INP(n1561), .ZN(n1520) );
  INVX0 U240 ( .INP(n1561), .ZN(n1521) );
  INVX0 U241 ( .INP(n1560), .ZN(n1522) );
  INVX0 U242 ( .INP(n1560), .ZN(n1523) );
  INVX0 U243 ( .INP(n1560), .ZN(n1524) );
  INVX0 U244 ( .INP(n1560), .ZN(n1525) );
  INVX0 U245 ( .INP(n1560), .ZN(n1526) );
  INVX0 U246 ( .INP(n1560), .ZN(n1531) );
  INVX0 U247 ( .INP(n1559), .ZN(n1536) );
  INVX0 U248 ( .INP(n1560), .ZN(n1530) );
  INVX0 U249 ( .INP(n1560), .ZN(n1528) );
  INVX0 U250 ( .INP(n1560), .ZN(n1529) );
  INVX0 U251 ( .INP(n1564), .ZN(n1479) );
  INVX0 U252 ( .INP(n1564), .ZN(n1474) );
  INVX0 U253 ( .INP(n1564), .ZN(n1475) );
  INVX0 U254 ( .INP(n1564), .ZN(n1477) );
  INVX0 U255 ( .INP(n1564), .ZN(n1478) );
  INVX0 U256 ( .INP(n1564), .ZN(n1476) );
  INVX0 U257 ( .INP(n1377), .ZN(n1376) );
  INVX0 U258 ( .INP(n1586), .ZN(n1578) );
  INVX0 U259 ( .INP(n1586), .ZN(n1579) );
  INVX0 U260 ( .INP(n1586), .ZN(n1580) );
  INVX0 U261 ( .INP(n1586), .ZN(n1581) );
  INVX0 U262 ( .INP(n1586), .ZN(n1582) );
  INVX0 U263 ( .INP(n1586), .ZN(n1583) );
  INVX0 U264 ( .INP(n1586), .ZN(n1584) );
  INVX0 U265 ( .INP(n1586), .ZN(n1577) );
  INVX0 U266 ( .INP(n1586), .ZN(n1574) );
  INVX0 U267 ( .INP(n1586), .ZN(n1576) );
  INVX0 U268 ( .INP(n1586), .ZN(n1575) );
  INVX0 U269 ( .INP(n1587), .ZN(n1569) );
  INVX0 U270 ( .INP(n1587), .ZN(n1570) );
  INVX0 U271 ( .INP(n1587), .ZN(n1568) );
  INVX0 U272 ( .INP(n1587), .ZN(n1571) );
  INVX0 U273 ( .INP(n1587), .ZN(n1573) );
  INVX0 U274 ( .INP(n1587), .ZN(n1572) );
  INVX0 U275 ( .INP(n1587), .ZN(n1567) );
  INVX0 U276 ( .INP(n1587), .ZN(n1565) );
  INVX0 U277 ( .INP(n1587), .ZN(n1566) );
  INVX0 U278 ( .INP(n1558), .ZN(n1557) );
  INVX0 U279 ( .INP(n1586), .ZN(n1585) );
  INVX0 U280 ( .INP(n1588), .ZN(n1357) );
  INVX0 U281 ( .INP(\fpu_add_exp_dp/n448 ), .ZN(n1586) );
  INVX0 U282 ( .INP(\fpu_add_exp_dp/n448 ), .ZN(n1587) );
  NBUFFX2 U283 ( .INP(n1342), .Z(n1563) );
  NBUFFX2 U284 ( .INP(n1342), .Z(n1562) );
  NBUFFX2 U285 ( .INP(n1342), .Z(n1564) );
  NBUFFX2 U286 ( .INP(n1342), .Z(n1558) );
  NBUFFX2 U287 ( .INP(n1342), .Z(n1561) );
  NBUFFX2 U288 ( .INP(n1342), .Z(n1559) );
  NBUFFX2 U289 ( .INP(n1342), .Z(n1560) );
  NBUFFX2 U290 ( .INP(n1341), .Z(n1377) );
  NBUFFX2 U291 ( .INP(n1341), .Z(n1378) );
  OR2X1 U292 ( .IN1(n1343), .IN2(se_add_frac), .Q(n1341) );
  OR2X1 U293 ( .IN1(\fpu_add_frac_dp/n998 ), .IN2(\fpu_add_frac_dp/n2189 ), 
        .Q(n1342) );
  AO22X1 U294 ( .IN1(n1343), .IN2(n612), .IN3(inq_in1[0]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4285 ) );
  AO22X1 U295 ( .IN1(n1349), .IN2(n93), .IN3(inq_in1[1]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4284 ) );
  AO22X1 U296 ( .IN1(n1349), .IN2(n182), .IN3(inq_in1[2]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4283 ) );
  AO22X1 U297 ( .IN1(n1349), .IN2(n599), .IN3(inq_in1[3]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4282 ) );
  AO22X1 U298 ( .IN1(n1349), .IN2(n183), .IN3(inq_in1[4]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4281 ) );
  AO22X1 U299 ( .IN1(n1349), .IN2(n600), .IN3(inq_in1[5]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4280 ) );
  AO22X1 U300 ( .IN1(n1349), .IN2(n184), .IN3(inq_in1[6]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4279 ) );
  AO22X1 U301 ( .IN1(n1349), .IN2(n601), .IN3(inq_in1[7]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4278 ) );
  AO22X1 U302 ( .IN1(n1349), .IN2(n185), .IN3(inq_in1[8]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4277 ) );
  AO22X1 U303 ( .IN1(n1349), .IN2(n602), .IN3(inq_in1[9]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4276 ) );
  AO22X1 U304 ( .IN1(n1349), .IN2(n186), .IN3(inq_in1[10]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4275 ) );
  AO22X1 U305 ( .IN1(n1349), .IN2(n603), .IN3(inq_in1[11]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4274 ) );
  AO22X1 U306 ( .IN1(n1349), .IN2(n187), .IN3(inq_in1[12]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4273 ) );
  AO22X1 U307 ( .IN1(n1348), .IN2(n604), .IN3(inq_in1[13]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4272 ) );
  AO22X1 U308 ( .IN1(n1348), .IN2(n188), .IN3(inq_in1[14]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4271 ) );
  AO22X1 U309 ( .IN1(n1348), .IN2(n605), .IN3(inq_in1[15]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4270 ) );
  AO22X1 U310 ( .IN1(n1348), .IN2(n189), .IN3(inq_in1[16]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4269 ) );
  AO22X1 U311 ( .IN1(n1348), .IN2(n606), .IN3(inq_in1[17]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4268 ) );
  AO22X1 U312 ( .IN1(n1348), .IN2(n190), .IN3(inq_in1[18]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4267 ) );
  AO22X1 U313 ( .IN1(n1348), .IN2(n607), .IN3(inq_in1[19]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4266 ) );
  AO22X1 U314 ( .IN1(n1348), .IN2(n191), .IN3(inq_in1[20]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4265 ) );
  AO22X1 U315 ( .IN1(n1348), .IN2(n608), .IN3(inq_in1[21]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4264 ) );
  AO22X1 U316 ( .IN1(n1348), .IN2(n192), .IN3(inq_in1[22]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4263 ) );
  AO22X1 U317 ( .IN1(n1348), .IN2(n609), .IN3(inq_in1[23]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4262 ) );
  AO22X1 U318 ( .IN1(n1348), .IN2(n193), .IN3(inq_in1[24]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4261 ) );
  AO22X1 U319 ( .IN1(n1348), .IN2(n610), .IN3(inq_in1[25]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4260 ) );
  AO22X1 U320 ( .IN1(n1348), .IN2(n194), .IN3(inq_in1[26]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4259 ) );
  AO22X1 U321 ( .IN1(n1348), .IN2(n611), .IN3(inq_in1[27]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4258 ) );
  AO22X1 U322 ( .IN1(n1348), .IN2(n207), .IN3(inq_in1[28]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4257 ) );
  AO22X1 U323 ( .IN1(n1348), .IN2(n644), .IN3(inq_in1[29]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4256 ) );
  AO22X1 U324 ( .IN1(n1347), .IN2(n698), .IN3(inq_in1[30]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4255 ) );
  AO22X1 U325 ( .IN1(n1347), .IN2(n699), .IN3(inq_in1[31]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4254 ) );
  AO22X1 U326 ( .IN1(n1347), .IN2(n176), .IN3(inq_in1[32]), .IN4(n1374), .Q(
        \fpu_add_frac_dp/n4253 ) );
  AO22X1 U327 ( .IN1(n1347), .IN2(n208), .IN3(inq_in1[33]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4252 ) );
  AO22X1 U328 ( .IN1(n1347), .IN2(n99), .IN3(inq_in1[34]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4251 ) );
  AO22X1 U329 ( .IN1(n1347), .IN2(n614), .IN3(inq_in1[35]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4250 ) );
  AO22X1 U330 ( .IN1(n1347), .IN2(n615), .IN3(inq_in1[36]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4249 ) );
  AO22X1 U331 ( .IN1(n1347), .IN2(n209), .IN3(inq_in1[37]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4248 ) );
  AO22X1 U332 ( .IN1(n1347), .IN2(n210), .IN3(inq_in1[38]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4247 ) );
  AO22X1 U333 ( .IN1(n1347), .IN2(n211), .IN3(inq_in1[39]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4246 ) );
  AO22X1 U334 ( .IN1(n1347), .IN2(n616), .IN3(inq_in1[40]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4245 ) );
  AO22X1 U335 ( .IN1(n1347), .IN2(n617), .IN3(inq_in1[41]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4244 ) );
  AO22X1 U336 ( .IN1(n1347), .IN2(n618), .IN3(inq_in1[42]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4243 ) );
  AO22X1 U337 ( .IN1(n1347), .IN2(n212), .IN3(inq_in1[43]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4242 ) );
  AO22X1 U338 ( .IN1(n1347), .IN2(n213), .IN3(inq_in1[44]), .IN4(n1373), .Q(
        \fpu_add_frac_dp/n4241 ) );
  AO22X1 U339 ( .IN1(n1347), .IN2(n214), .IN3(inq_in1[45]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4240 ) );
  AO22X1 U340 ( .IN1(n1347), .IN2(n619), .IN3(inq_in1[46]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4239 ) );
  AO22X1 U341 ( .IN1(n1346), .IN2(n620), .IN3(inq_in1[47]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4238 ) );
  AO22X1 U342 ( .IN1(n1346), .IN2(n621), .IN3(inq_in1[48]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4237 ) );
  AO22X1 U343 ( .IN1(n1346), .IN2(n215), .IN3(inq_in1[49]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4236 ) );
  AO22X1 U344 ( .IN1(n1346), .IN2(n216), .IN3(inq_in1[50]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4235 ) );
  AO22X1 U345 ( .IN1(n1346), .IN2(n206), .IN3(inq_in1[51]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4234 ) );
  AO22X1 U346 ( .IN1(n1346), .IN2(n688), .IN3(inq_in1[52]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4233 ) );
  AO22X1 U347 ( .IN1(n1346), .IN2(n689), .IN3(inq_in1[53]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4232 ) );
  AO22X1 U348 ( .IN1(n1346), .IN2(n705), .IN3(inq_in1[54]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4231 ) );
  AO22X1 U349 ( .IN1(n1346), .IN2(n1188), .IN3(inq_in1[55]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4230 ) );
  AO22X1 U350 ( .IN1(n1346), .IN2(n1189), .IN3(inq_in1[56]), .IN4(n1372), .Q(
        \fpu_add_frac_dp/n4229 ) );
  AO22X1 U351 ( .IN1(n1346), .IN2(n714), .IN3(inq_in1[57]), .IN4(n1371), .Q(
        \fpu_add_frac_dp/n4228 ) );
  AO22X1 U352 ( .IN1(n1346), .IN2(n1190), .IN3(inq_in1[58]), .IN4(n1371), .Q(
        \fpu_add_frac_dp/n4227 ) );
  AO22X1 U353 ( .IN1(n1346), .IN2(n713), .IN3(inq_in1[59]), .IN4(n1371), .Q(
        \fpu_add_frac_dp/n4226 ) );
  AO22X1 U354 ( .IN1(n1346), .IN2(n712), .IN3(inq_in1[60]), .IN4(n1371), .Q(
        \fpu_add_frac_dp/n4225 ) );
  AO22X1 U355 ( .IN1(n1346), .IN2(n1191), .IN3(inq_in1[61]), .IN4(n1371), .Q(
        \fpu_add_frac_dp/n4224 ) );
  AO22X1 U356 ( .IN1(n1346), .IN2(n715), .IN3(inq_in1[62]), .IN4(n1371), .Q(
        \fpu_add_frac_dp/n4223 ) );
  AO22X1 U357 ( .IN1(\fpu_add_frac_dp/n2493 ), .IN2(n1356), .IN3(inq_in1[0]), 
        .IN4(n1371), .Q(\fpu_add_frac_dp/n4222 ) );
  AO22X1 U358 ( .IN1(n1345), .IN2(n1185), .IN3(inq_in1[1]), .IN4(n1371), .Q(
        \fpu_add_frac_dp/n4221 ) );
  AO22X1 U359 ( .IN1(n1345), .IN2(n745), .IN3(inq_in1[2]), .IN4(n1371), .Q(
        \fpu_add_frac_dp/n4220 ) );
  AO22X1 U360 ( .IN1(\fpu_add_frac_dp/n2296 ), .IN2(n1356), .IN3(inq_in1[3]), 
        .IN4(n1371), .Q(\fpu_add_frac_dp/n4219 ) );
  AO22X1 U361 ( .IN1(n1345), .IN2(n695), .IN3(inq_in1[4]), .IN4(n1371), .Q(
        \fpu_add_frac_dp/n4218 ) );
  AO22X1 U362 ( .IN1(n1345), .IN2(n1128), .IN3(inq_in1[5]), .IN4(n1371), .Q(
        \fpu_add_frac_dp/n4217 ) );
  AO22X1 U363 ( .IN1(n1345), .IN2(n1133), .IN3(inq_in1[6]), .IN4(n1370), .Q(
        \fpu_add_frac_dp/n4216 ) );
  AO22X1 U364 ( .IN1(n1345), .IN2(n1195), .IN3(inq_in1[7]), .IN4(n1370), .Q(
        \fpu_add_frac_dp/n4215 ) );
  AO22X1 U365 ( .IN1(n1345), .IN2(n1146), .IN3(inq_in1[8]), .IN4(n1370), .Q(
        \fpu_add_frac_dp/n4214 ) );
  AO22X1 U366 ( .IN1(n1345), .IN2(n577), .IN3(inq_in1[9]), .IN4(n1370), .Q(
        \fpu_add_frac_dp/n4213 ) );
  AO22X1 U367 ( .IN1(n1345), .IN2(n145), .IN3(inq_in1[10]), .IN4(n1370), .Q(
        \fpu_add_frac_dp/n4212 ) );
  AO22X1 U368 ( .IN1(n1345), .IN2(n854), .IN3(inq_in1[11]), .IN4(n1370), .Q(
        \fpu_add_frac_dp/n4211 ) );
  AO22X1 U369 ( .IN1(\fpu_add_frac_dp/n2484 ), .IN2(n1356), .IN3(inq_in1[12]), 
        .IN4(n1370), .Q(\fpu_add_frac_dp/n4210 ) );
  AO22X1 U370 ( .IN1(n1345), .IN2(n1184), .IN3(inq_in1[13]), .IN4(n1370), .Q(
        \fpu_add_frac_dp/n4209 ) );
  AO22X1 U371 ( .IN1(n1345), .IN2(n988), .IN3(inq_in1[14]), .IN4(n1370), .Q(
        \fpu_add_frac_dp/n4208 ) );
  AO22X1 U372 ( .IN1(\fpu_add_frac_dp/n2453 ), .IN2(n1356), .IN3(inq_in1[15]), 
        .IN4(n1370), .Q(\fpu_add_frac_dp/n4207 ) );
  AO22X1 U373 ( .IN1(n1345), .IN2(n703), .IN3(inq_in1[16]), .IN4(n1370), .Q(
        \fpu_add_frac_dp/n4206 ) );
  AO22X1 U374 ( .IN1(n1345), .IN2(n853), .IN3(inq_in1[17]), .IN4(n1370), .Q(
        \fpu_add_frac_dp/n4205 ) );
  AO22X1 U375 ( .IN1(n1345), .IN2(n1153), .IN3(inq_in1[18]), .IN4(n1369), .Q(
        \fpu_add_frac_dp/n4204 ) );
  AO22X1 U376 ( .IN1(n1345), .IN2(n1197), .IN3(inq_in1[19]), .IN4(n1369), .Q(
        \fpu_add_frac_dp/n4203 ) );
  AO22X1 U377 ( .IN1(n1345), .IN2(n1143), .IN3(inq_in1[20]), .IN4(n1369), .Q(
        \fpu_add_frac_dp/n4202 ) );
  AO22X1 U378 ( .IN1(\fpu_add_frac_dp/n2444 ), .IN2(n1356), .IN3(inq_in1[21]), 
        .IN4(n1369), .Q(\fpu_add_frac_dp/n4201 ) );
  AO22X1 U379 ( .IN1(n1344), .IN2(n1204), .IN3(inq_in1[22]), .IN4(n1369), .Q(
        \fpu_add_frac_dp/n4200 ) );
  AO22X1 U380 ( .IN1(n1344), .IN2(n1206), .IN3(inq_in1[23]), .IN4(n1369), .Q(
        \fpu_add_frac_dp/n4199 ) );
  AO22X1 U381 ( .IN1(\fpu_add_frac_dp/n2488 ), .IN2(n1356), .IN3(inq_in1[24]), 
        .IN4(n1369), .Q(\fpu_add_frac_dp/n4198 ) );
  AO22X1 U382 ( .IN1(n1344), .IN2(n1209), .IN3(inq_in1[25]), .IN4(n1369), .Q(
        \fpu_add_frac_dp/n4197 ) );
  AO22X1 U383 ( .IN1(n1344), .IN2(n550), .IN3(inq_in1[26]), .IN4(n1369), .Q(
        \fpu_add_frac_dp/n4196 ) );
  AO22X1 U384 ( .IN1(n1344), .IN2(n647), .IN3(inq_in1[27]), .IN4(n1369), .Q(
        \fpu_add_frac_dp/n4195 ) );
  AO22X1 U385 ( .IN1(n1344), .IN2(n54), .IN3(inq_in1[28]), .IN4(n1369), .Q(
        \fpu_add_frac_dp/n4194 ) );
  AO22X1 U386 ( .IN1(n1344), .IN2(n856), .IN3(inq_in1[29]), .IN4(n1369), .Q(
        \fpu_add_frac_dp/n4193 ) );
  AO22X1 U387 ( .IN1(\fpu_add_frac_dp/n2445 ), .IN2(n1356), .IN3(inq_in1[30]), 
        .IN4(n1368), .Q(\fpu_add_frac_dp/n4192 ) );
  AO22X1 U388 ( .IN1(n1344), .IN2(n704), .IN3(inq_in1[31]), .IN4(n1368), .Q(
        \fpu_add_frac_dp/n4191 ) );
  AO22X1 U389 ( .IN1(n1344), .IN2(n855), .IN3(inq_in1[32]), .IN4(n1368), .Q(
        \fpu_add_frac_dp/n4190 ) );
  AO22X1 U390 ( .IN1(\fpu_add_frac_dp/n2295 ), .IN2(n1356), .IN3(inq_in1[33]), 
        .IN4(n1368), .Q(\fpu_add_frac_dp/n4189 ) );
  AO22X1 U391 ( .IN1(n1344), .IN2(n857), .IN3(inq_in1[34]), .IN4(n1368), .Q(
        \fpu_add_frac_dp/n4188 ) );
  AO22X1 U392 ( .IN1(n1344), .IN2(n1215), .IN3(inq_in1[35]), .IN4(n1368), .Q(
        \fpu_add_frac_dp/n4187 ) );
  AO22X1 U393 ( .IN1(n1344), .IN2(n292), .IN3(inq_in1[36]), .IN4(n1368), .Q(
        \fpu_add_frac_dp/n4186 ) );
  AO22X1 U394 ( .IN1(n1344), .IN2(n125), .IN3(inq_in1[37]), .IN4(n1368), .Q(
        \fpu_add_frac_dp/n4185 ) );
  AO22X1 U395 ( .IN1(n1344), .IN2(n46), .IN3(inq_in1[38]), .IN4(n1368), .Q(
        \fpu_add_frac_dp/n4184 ) );
  AO22X1 U396 ( .IN1(\fpu_add_frac_dp/n2452 ), .IN2(n1356), .IN3(inq_in1[39]), 
        .IN4(n1368), .Q(\fpu_add_frac_dp/n4183 ) );
  AO22X1 U397 ( .IN1(n1344), .IN2(n709), .IN3(inq_in1[40]), .IN4(n1368), .Q(
        \fpu_add_frac_dp/n4182 ) );
  AO22X1 U398 ( .IN1(n1344), .IN2(n1129), .IN3(inq_in1[41]), .IN4(n1368), .Q(
        \fpu_add_frac_dp/n4181 ) );
  AO22X1 U399 ( .IN1(\fpu_add_frac_dp/n2462 ), .IN2(n1356), .IN3(inq_in1[42]), 
        .IN4(n1367), .Q(\fpu_add_frac_dp/n4180 ) );
  AO22X1 U400 ( .IN1(n1344), .IN2(n848), .IN3(inq_in1[43]), .IN4(n1367), .Q(
        \fpu_add_frac_dp/n4179 ) );
  AO22X1 U401 ( .IN1(n1343), .IN2(n57), .IN3(inq_in1[44]), .IN4(n1367), .Q(
        \fpu_add_frac_dp/n4178 ) );
  AO22X1 U402 ( .IN1(n1343), .IN2(n677), .IN3(inq_in1[45]), .IN4(n1367), .Q(
        \fpu_add_frac_dp/n4177 ) );
  AO22X1 U403 ( .IN1(n1343), .IN2(n1198), .IN3(inq_in1[46]), .IN4(n1367), .Q(
        \fpu_add_frac_dp/n4176 ) );
  AO22X1 U404 ( .IN1(n1343), .IN2(n1202), .IN3(inq_in1[47]), .IN4(n1367), .Q(
        \fpu_add_frac_dp/n4175 ) );
  AO22X1 U405 ( .IN1(\fpu_add_frac_dp/n2476 ), .IN2(n1588), .IN3(inq_in1[48]), 
        .IN4(n1367), .Q(\fpu_add_frac_dp/n4174 ) );
  AO22X1 U406 ( .IN1(n1343), .IN2(n917), .IN3(inq_in1[49]), .IN4(n1367), .Q(
        \fpu_add_frac_dp/n4173 ) );
  AO22X1 U407 ( .IN1(\fpu_add_frac_dp/n2350 ), .IN2(n1354), .IN3(inq_in1[50]), 
        .IN4(n1367), .Q(\fpu_add_frac_dp/n4172 ) );
  AO22X1 U408 ( .IN1(n1343), .IN2(n340), .IN3(inq_in1[51]), .IN4(n1367), .Q(
        \fpu_add_frac_dp/n4171 ) );
  AO22X1 U409 ( .IN1(n1343), .IN2(n548), .IN3(inq_in1[52]), .IN4(n1367), .Q(
        \fpu_add_frac_dp/n4170 ) );
  AO22X1 U410 ( .IN1(n1343), .IN2(n747), .IN3(inq_in1[53]), .IN4(n1367), .Q(
        \fpu_add_frac_dp/n4169 ) );
  AO22X1 U411 ( .IN1(n1343), .IN2(n283), .IN3(inq_in1[54]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4168 ) );
  AO22X1 U412 ( .IN1(n1343), .IN2(n36), .IN3(inq_in2[0]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4167 ) );
  AO22X1 U413 ( .IN1(n1349), .IN2(n170), .IN3(inq_in2[1]), .IN4(n1376), .Q(
        \fpu_add_frac_dp/n4166 ) );
  AO22X1 U414 ( .IN1(n1343), .IN2(n10), .IN3(inq_in2[2]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4165 ) );
  AO22X1 U415 ( .IN1(n1343), .IN2(n1589), .IN3(inq_in2[3]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4164 ) );
  AO22X1 U416 ( .IN1(n1343), .IN2(n11), .IN3(inq_in2[4]), .IN4(n1363), .Q(
        \fpu_add_frac_dp/n4163 ) );
  AO22X1 U417 ( .IN1(n1346), .IN2(n30), .IN3(inq_in2[5]), .IN4(n1362), .Q(
        \fpu_add_frac_dp/n4162 ) );
  AO22X1 U418 ( .IN1(n1349), .IN2(n79), .IN3(inq_in2[6]), .IN4(n1361), .Q(
        \fpu_add_frac_dp/n4161 ) );
  AO22X1 U419 ( .IN1(n1349), .IN2(n31), .IN3(inq_in2[7]), .IN4(n1360), .Q(
        \fpu_add_frac_dp/n4160 ) );
  AO22X1 U420 ( .IN1(n1349), .IN2(n80), .IN3(inq_in2[8]), .IN4(n1359), .Q(
        \fpu_add_frac_dp/n4159 ) );
  AO22X1 U421 ( .IN1(n1349), .IN2(n32), .IN3(inq_in2[9]), .IN4(n1358), .Q(
        \fpu_add_frac_dp/n4158 ) );
  AO22X1 U422 ( .IN1(n1350), .IN2(n81), .IN3(inq_in2[10]), .IN4(n1375), .Q(
        \fpu_add_frac_dp/n4157 ) );
  AO22X1 U423 ( .IN1(n1350), .IN2(n39), .IN3(inq_in2[11]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4156 ) );
  AO22X1 U424 ( .IN1(n1350), .IN2(n120), .IN3(inq_in2[12]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4155 ) );
  AO22X1 U425 ( .IN1(n1350), .IN2(n52), .IN3(inq_in2[13]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4154 ) );
  AO22X1 U426 ( .IN1(n1350), .IN2(n121), .IN3(inq_in2[14]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4153 ) );
  AO22X1 U427 ( .IN1(n1350), .IN2(n53), .IN3(inq_in2[15]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4152 ) );
  AO22X1 U428 ( .IN1(n1350), .IN2(n122), .IN3(inq_in2[16]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4151 ) );
  AO22X1 U429 ( .IN1(n1350), .IN2(n272), .IN3(inq_in2[17]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4150 ) );
  AO22X1 U430 ( .IN1(n1350), .IN2(n633), .IN3(inq_in2[18]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4149 ) );
  AO22X1 U431 ( .IN1(n1350), .IN2(n273), .IN3(inq_in2[19]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4148 ) );
  AO22X1 U432 ( .IN1(n1350), .IN2(n634), .IN3(inq_in2[20]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4147 ) );
  AO22X1 U433 ( .IN1(n1350), .IN2(n274), .IN3(inq_in2[21]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4146 ) );
  AO22X1 U434 ( .IN1(n1350), .IN2(n635), .IN3(inq_in2[22]), .IN4(n1366), .Q(
        \fpu_add_frac_dp/n4145 ) );
  AO22X1 U435 ( .IN1(n1350), .IN2(n275), .IN3(inq_in2[23]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4144 ) );
  AO22X1 U436 ( .IN1(n1351), .IN2(n636), .IN3(inq_in2[24]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4143 ) );
  AO22X1 U437 ( .IN1(n1351), .IN2(n276), .IN3(inq_in2[25]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4142 ) );
  AO22X1 U438 ( .IN1(n1350), .IN2(n637), .IN3(inq_in2[26]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4141 ) );
  AO22X1 U439 ( .IN1(n1351), .IN2(n277), .IN3(inq_in2[27]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4140 ) );
  AO22X1 U440 ( .IN1(n1351), .IN2(n639), .IN3(inq_in2[28]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4139 ) );
  AO22X1 U441 ( .IN1(n1351), .IN2(n112), .IN3(inq_in2[29]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4138 ) );
  AO22X1 U442 ( .IN1(n1351), .IN2(n113), .IN3(inq_in2[30]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4137 ) );
  AO22X1 U443 ( .IN1(n1351), .IN2(n114), .IN3(inq_in2[31]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4136 ) );
  AO22X1 U444 ( .IN1(n1351), .IN2(n7), .IN3(inq_in2[32]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4135 ) );
  AO22X1 U445 ( .IN1(n1351), .IN2(n8), .IN3(inq_in2[33]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4134 ) );
  AO22X1 U446 ( .IN1(n1351), .IN2(n9), .IN3(inq_in2[34]), .IN4(n1365), .Q(
        \fpu_add_frac_dp/n4133 ) );
  AO22X1 U447 ( .IN1(n1351), .IN2(n24), .IN3(inq_in2[35]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4132 ) );
  AO22X1 U448 ( .IN1(n1351), .IN2(n25), .IN3(inq_in2[36]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4131 ) );
  AO22X1 U449 ( .IN1(n1351), .IN2(n26), .IN3(inq_in2[37]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4130 ) );
  AO22X1 U450 ( .IN1(n1352), .IN2(n76), .IN3(inq_in2[38]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4129 ) );
  AO22X1 U451 ( .IN1(n1352), .IN2(n77), .IN3(inq_in2[39]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4128 ) );
  AO22X1 U452 ( .IN1(n1351), .IN2(n167), .IN3(inq_in2[40]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4127 ) );
  AO22X1 U453 ( .IN1(n1352), .IN2(n27), .IN3(inq_in2[41]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4126 ) );
  AO22X1 U454 ( .IN1(n1352), .IN2(n28), .IN3(inq_in2[42]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4125 ) );
  AO22X1 U455 ( .IN1(n1352), .IN2(n29), .IN3(inq_in2[43]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4124 ) );
  AO22X1 U456 ( .IN1(n1352), .IN2(n163), .IN3(inq_in2[44]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4123 ) );
  AO22X1 U457 ( .IN1(n1352), .IN2(n164), .IN3(inq_in2[45]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4122 ) );
  AO22X1 U458 ( .IN1(n1352), .IN2(n587), .IN3(inq_in2[46]), .IN4(n1364), .Q(
        \fpu_add_frac_dp/n4121 ) );
  AO22X1 U459 ( .IN1(n1352), .IN2(n588), .IN3(inq_in2[47]), .IN4(n1363), .Q(
        \fpu_add_frac_dp/n4120 ) );
  AO22X1 U460 ( .IN1(n1352), .IN2(n589), .IN3(inq_in2[48]), .IN4(n1363), .Q(
        \fpu_add_frac_dp/n4119 ) );
  AO22X1 U461 ( .IN1(n1352), .IN2(n78), .IN3(inq_in2[49]), .IN4(n1363), .Q(
        \fpu_add_frac_dp/n4118 ) );
  AO22X1 U462 ( .IN1(n1352), .IN2(n165), .IN3(inq_in2[50]), .IN4(n1363), .Q(
        \fpu_add_frac_dp/n4117 ) );
  AO22X1 U463 ( .IN1(n1351), .IN2(n169), .IN3(inq_in2[51]), .IN4(n1363), .Q(
        \fpu_add_frac_dp/n4116 ) );
  AO22X1 U464 ( .IN1(n1353), .IN2(n591), .IN3(inq_in2[52]), .IN4(n1363), .Q(
        \fpu_add_frac_dp/n4115 ) );
  AO22X1 U465 ( .IN1(n1353), .IN2(n592), .IN3(inq_in2[53]), .IN4(n1363), .Q(
        \fpu_add_frac_dp/n4114 ) );
  AO22X1 U466 ( .IN1(n1353), .IN2(n593), .IN3(inq_in2[54]), .IN4(n1363), .Q(
        \fpu_add_frac_dp/n4113 ) );
  AO22X1 U467 ( .IN1(\fpu_add_frac_dp/n2446 ), .IN2(n1356), .IN3(inq_in2[55]), 
        .IN4(n1363), .Q(\fpu_add_frac_dp/n4112 ) );
  AO22X1 U468 ( .IN1(\fpu_add_frac_dp/n2473 ), .IN2(n1356), .IN3(inq_in2[56]), 
        .IN4(n1363), .Q(\fpu_add_frac_dp/n4111 ) );
  AO22X1 U469 ( .IN1(\fpu_add_frac_dp/n2466 ), .IN2(n1356), .IN3(inq_in2[57]), 
        .IN4(n1363), .Q(\fpu_add_frac_dp/n4110 ) );
  AO22X1 U470 ( .IN1(\fpu_add_frac_dp/n2474 ), .IN2(n1356), .IN3(inq_in2[58]), 
        .IN4(n1363), .Q(\fpu_add_frac_dp/n4109 ) );
  AO22X1 U471 ( .IN1(\fpu_add_frac_dp/n2467 ), .IN2(n1356), .IN3(inq_in2[59]), 
        .IN4(n1362), .Q(\fpu_add_frac_dp/n4108 ) );
  AO22X1 U472 ( .IN1(\fpu_add_frac_dp/n2475 ), .IN2(n1356), .IN3(inq_in2[60]), 
        .IN4(n1362), .Q(\fpu_add_frac_dp/n4107 ) );
  AO22X1 U473 ( .IN1(\fpu_add_frac_dp/n2468 ), .IN2(n1356), .IN3(inq_in2[61]), 
        .IN4(n1362), .Q(\fpu_add_frac_dp/n4106 ) );
  AO22X1 U474 ( .IN1(\fpu_add_frac_dp/n2469 ), .IN2(n1355), .IN3(inq_in2[62]), 
        .IN4(n1362), .Q(\fpu_add_frac_dp/n4105 ) );
  AO22X1 U475 ( .IN1(n1353), .IN2(n1080), .IN3(inq_in2[63]), .IN4(n1362), .Q(
        \fpu_add_frac_dp/n4104 ) );
  AO22X1 U476 ( .IN1(n1353), .IN2(n702), .IN3(inq_in2[0]), .IN4(n1362), .Q(
        \fpu_add_frac_dp/n4103 ) );
  AO22X1 U477 ( .IN1(\fpu_add_frac_dp/n2455 ), .IN2(n1355), .IN3(inq_in2[1]), 
        .IN4(n1362), .Q(\fpu_add_frac_dp/n4102 ) );
  AO22X1 U478 ( .IN1(n1353), .IN2(n337), .IN3(inq_in2[2]), .IN4(n1362), .Q(
        \fpu_add_frac_dp/n4101 ) );
  AO22X1 U479 ( .IN1(n1353), .IN2(n1205), .IN3(inq_in2[3]), .IN4(n1362), .Q(
        \fpu_add_frac_dp/n4100 ) );
  AO22X1 U480 ( .IN1(n1352), .IN2(n900), .IN3(inq_in2[4]), .IN4(n1362), .Q(
        \fpu_add_frac_dp/n4099 ) );
  AO22X1 U481 ( .IN1(\fpu_add_frac_dp/n2459 ), .IN2(n1355), .IN3(inq_in2[5]), 
        .IN4(n1362), .Q(\fpu_add_frac_dp/n4098 ) );
  AO22X1 U482 ( .IN1(\fpu_add_frac_dp/n2490 ), .IN2(n1355), .IN3(inq_in2[6]), 
        .IN4(n1362), .Q(\fpu_add_frac_dp/n4097 ) );
  AO22X1 U483 ( .IN1(\fpu_add_frac_dp/n2489 ), .IN2(n1355), .IN3(inq_in2[7]), 
        .IN4(n1361), .Q(\fpu_add_frac_dp/n4096 ) );
  AO22X1 U484 ( .IN1(\fpu_add_frac_dp/n2472 ), .IN2(n1355), .IN3(inq_in2[8]), 
        .IN4(n1361), .Q(\fpu_add_frac_dp/n4095 ) );
  AO22X1 U485 ( .IN1(n1354), .IN2(n697), .IN3(inq_in2[9]), .IN4(n1361), .Q(
        \fpu_add_frac_dp/n4094 ) );
  AO22X1 U486 ( .IN1(\fpu_add_frac_dp/n2483 ), .IN2(n1355), .IN3(inq_in2[10]), 
        .IN4(n1361), .Q(\fpu_add_frac_dp/n4093 ) );
  AO22X1 U487 ( .IN1(\fpu_add_frac_dp/n2457 ), .IN2(n1355), .IN3(inq_in2[11]), 
        .IN4(n1361), .Q(\fpu_add_frac_dp/n4092 ) );
  AO22X1 U488 ( .IN1(n1354), .IN2(n670), .IN3(inq_in2[12]), .IN4(n1361), .Q(
        \fpu_add_frac_dp/n4091 ) );
  AO22X1 U489 ( .IN1(n1354), .IN2(n330), .IN3(inq_in2[13]), .IN4(n1361), .Q(
        \fpu_add_frac_dp/n4090 ) );
  AO22X1 U490 ( .IN1(n1353), .IN2(n1007), .IN3(inq_in2[14]), .IN4(n1361), .Q(
        \fpu_add_frac_dp/n4089 ) );
  AO22X1 U491 ( .IN1(n1353), .IN2(n1203), .IN3(inq_in2[15]), .IN4(n1361), .Q(
        \fpu_add_frac_dp/n4088 ) );
  AO22X1 U492 ( .IN1(n1354), .IN2(n1193), .IN3(inq_in2[16]), .IN4(n1361), .Q(
        \fpu_add_frac_dp/n4087 ) );
  AO22X1 U493 ( .IN1(n1353), .IN2(n1131), .IN3(inq_in2[17]), .IN4(n1361), .Q(
        \fpu_add_frac_dp/n4086 ) );
  AO22X1 U494 ( .IN1(n1354), .IN2(n1192), .IN3(inq_in2[18]), .IN4(n1361), .Q(
        \fpu_add_frac_dp/n4085 ) );
  AO22X1 U495 ( .IN1(\fpu_add_frac_dp/n2485 ), .IN2(n1355), .IN3(inq_in2[19]), 
        .IN4(n1360), .Q(\fpu_add_frac_dp/n4084 ) );
  AO22X1 U496 ( .IN1(\fpu_add_frac_dp/n2487 ), .IN2(n1355), .IN3(inq_in2[20]), 
        .IN4(n1360), .Q(\fpu_add_frac_dp/n4083 ) );
  AO22X1 U497 ( .IN1(n1354), .IN2(n335), .IN3(inq_in2[21]), .IN4(n1360), .Q(
        \fpu_add_frac_dp/n4082 ) );
  AO22X1 U498 ( .IN1(\fpu_add_frac_dp/n2492 ), .IN2(n1355), .IN3(inq_in2[22]), 
        .IN4(n1360), .Q(\fpu_add_frac_dp/n4081 ) );
  AO22X1 U499 ( .IN1(\fpu_add_frac_dp/n2458 ), .IN2(n1355), .IN3(inq_in2[23]), 
        .IN4(n1360), .Q(\fpu_add_frac_dp/n4080 ) );
  AO22X1 U500 ( .IN1(n1354), .IN2(n1127), .IN3(inq_in2[24]), .IN4(n1360), .Q(
        \fpu_add_frac_dp/n4079 ) );
  AO22X1 U501 ( .IN1(\fpu_add_frac_dp/n2486 ), .IN2(n1355), .IN3(inq_in2[25]), 
        .IN4(n1360), .Q(\fpu_add_frac_dp/n4078 ) );
  AO22X1 U502 ( .IN1(\fpu_add_frac_dp/n2482 ), .IN2(n1355), .IN3(inq_in2[26]), 
        .IN4(n1360), .Q(\fpu_add_frac_dp/n4077 ) );
  AO22X1 U503 ( .IN1(\fpu_add_frac_dp/n5608 ), .IN2(n1355), .IN3(inq_in2[27]), 
        .IN4(n1360), .Q(\fpu_add_frac_dp/n4076 ) );
  AO22X1 U504 ( .IN1(\fpu_add_frac_dp/n5605 ), .IN2(n1354), .IN3(inq_in2[28]), 
        .IN4(n1360), .Q(\fpu_add_frac_dp/n4075 ) );
  AO22X1 U505 ( .IN1(n1353), .IN2(n1132), .IN3(inq_in2[29]), .IN4(n1360), .Q(
        \fpu_add_frac_dp/n4074 ) );
  AO22X1 U506 ( .IN1(n1353), .IN2(n132), .IN3(inq_in2[30]), .IN4(n1360), .Q(
        \fpu_add_frac_dp/n4073 ) );
  AO22X1 U507 ( .IN1(n1353), .IN2(n1194), .IN3(inq_in2[31]), .IN4(n1359), .Q(
        \fpu_add_frac_dp/n4072 ) );
  AO22X1 U508 ( .IN1(\fpu_add_frac_dp/n5622 ), .IN2(n1354), .IN3(inq_in2[32]), 
        .IN4(n1359), .Q(\fpu_add_frac_dp/n4071 ) );
  AO22X1 U509 ( .IN1(n1353), .IN2(n326), .IN3(inq_in2[33]), .IN4(n1359), .Q(
        \fpu_add_frac_dp/n4070 ) );
  AO22X1 U510 ( .IN1(n1353), .IN2(n916), .IN3(inq_in2[34]), .IN4(n1359), .Q(
        \fpu_add_frac_dp/n4069 ) );
  AO22X1 U511 ( .IN1(\fpu_add_frac_dp/n5623 ), .IN2(n1354), .IN3(inq_in2[35]), 
        .IN4(n1359), .Q(\fpu_add_frac_dp/n4068 ) );
  AO22X1 U512 ( .IN1(n1352), .IN2(n1207), .IN3(inq_in2[36]), .IN4(n1359), .Q(
        \fpu_add_frac_dp/n4067 ) );
  AO22X1 U513 ( .IN1(\fpu_add_frac_dp/n5612 ), .IN2(n1354), .IN3(inq_in2[37]), 
        .IN4(n1359), .Q(\fpu_add_frac_dp/n4066 ) );
  AO22X1 U514 ( .IN1(\fpu_add_frac_dp/n5613 ), .IN2(n1354), .IN3(inq_in2[38]), 
        .IN4(n1359), .Q(\fpu_add_frac_dp/n4065 ) );
  AO22X1 U515 ( .IN1(n1352), .IN2(n141), .IN3(inq_in2[39]), .IN4(n1359), .Q(
        \fpu_add_frac_dp/n4064 ) );
  AO22X1 U516 ( .IN1(n1353), .IN2(n463), .IN3(inq_in2[40]), .IN4(n1359), .Q(
        \fpu_add_frac_dp/n4063 ) );
  AO22X1 U517 ( .IN1(\fpu_add_frac_dp/n5620 ), .IN2(n1355), .IN3(inq_in2[41]), 
        .IN4(n1359), .Q(\fpu_add_frac_dp/n4062 ) );
  AO22X1 U518 ( .IN1(n1352), .IN2(n1199), .IN3(inq_in2[42]), .IN4(n1359), .Q(
        \fpu_add_frac_dp/n4061 ) );
  AO22X1 U519 ( .IN1(n1352), .IN2(n763), .IN3(inq_in2[43]), .IN4(n1358), .Q(
        \fpu_add_frac_dp/n4060 ) );
  AO22X1 U520 ( .IN1(\fpu_add_frac_dp/n5621 ), .IN2(n1354), .IN3(inq_in2[44]), 
        .IN4(n1358), .Q(\fpu_add_frac_dp/n4059 ) );
  AO22X1 U521 ( .IN1(n1351), .IN2(n1208), .IN3(inq_in2[45]), .IN4(n1358), .Q(
        \fpu_add_frac_dp/n4058 ) );
  AO22X1 U522 ( .IN1(\fpu_add_frac_dp/n5611 ), .IN2(n1354), .IN3(inq_in2[46]), 
        .IN4(n1358), .Q(\fpu_add_frac_dp/n4057 ) );
  AO22X1 U523 ( .IN1(\fpu_add_frac_dp/n5624 ), .IN2(n1355), .IN3(inq_in2[47]), 
        .IN4(n1358), .Q(\fpu_add_frac_dp/n4056 ) );
  AO22X1 U524 ( .IN1(n1351), .IN2(n1211), .IN3(inq_in2[48]), .IN4(n1358), .Q(
        \fpu_add_frac_dp/n4055 ) );
  AO22X1 U525 ( .IN1(n1350), .IN2(n1065), .IN3(inq_in2[49]), .IN4(n1358), .Q(
        \fpu_add_frac_dp/n4054 ) );
  AO22X1 U526 ( .IN1(n1350), .IN2(n427), .IN3(inq_in2[50]), .IN4(n1358), .Q(
        \fpu_add_frac_dp/n4053 ) );
  AO22X1 U527 ( .IN1(\fpu_add_frac_dp/n2491 ), .IN2(n1354), .IN3(inq_in2[51]), 
        .IN4(n1358), .Q(\fpu_add_frac_dp/n4052 ) );
  AO22X1 U528 ( .IN1(\fpu_add_frac_dp/n5644 ), .IN2(n1354), .IN3(inq_in2[52]), 
        .IN4(n1358), .Q(\fpu_add_frac_dp/n4051 ) );
  AO22X1 U529 ( .IN1(n1353), .IN2(n650), .IN3(inq_in2[53]), .IN4(n1358), .Q(
        \fpu_add_frac_dp/n4050 ) );
  AO22X1 U530 ( .IN1(n1343), .IN2(n1130), .IN3(inq_in2[54]), .IN4(n1358), .Q(
        \fpu_add_frac_dp/n4049 ) );
  NOR2X0 U531 ( .IN1(a1stg_step), .IN2(se_add_frac), .QN(n1588) );
  AO22X1 U532 ( .IN1(n1426), .IN2(n307), .IN3(n1590), .IN4(n36), .Q(
        \fpu_add_frac_dp/n4048 ) );
  AO22X1 U533 ( .IN1(n1422), .IN2(n625), .IN3(n1590), .IN4(n170), .Q(
        \fpu_add_frac_dp/n4047 ) );
  AO22X1 U534 ( .IN1(n1422), .IN2(n220), .IN3(n1590), .IN4(n10), .Q(
        \fpu_add_frac_dp/n4046 ) );
  AO22X1 U535 ( .IN1(n1422), .IN2(n310), .IN3(n1590), .IN4(n1589), .Q(
        \fpu_add_frac_dp/n4045 ) );
  AO22X1 U536 ( .IN1(n1422), .IN2(n288), .IN3(n1590), .IN4(n11), .Q(
        \fpu_add_frac_dp/n4044 ) );
  AO22X1 U537 ( .IN1(n1422), .IN2(n223), .IN3(n1590), .IN4(n30), .Q(
        \fpu_add_frac_dp/n4043 ) );
  AO22X1 U538 ( .IN1(n1422), .IN2(n225), .IN3(n1590), .IN4(n79), .Q(
        \fpu_add_frac_dp/n4042 ) );
  AO22X1 U539 ( .IN1(n1422), .IN2(n222), .IN3(n1590), .IN4(n31), .Q(
        \fpu_add_frac_dp/n4041 ) );
  AO22X1 U540 ( .IN1(n1422), .IN2(n224), .IN3(n1590), .IN4(n80), .Q(
        \fpu_add_frac_dp/n4040 ) );
  AO22X1 U541 ( .IN1(n1422), .IN2(n261), .IN3(n1590), .IN4(n32), .Q(
        \fpu_add_frac_dp/n4039 ) );
  AO22X1 U542 ( .IN1(n1422), .IN2(n260), .IN3(n1590), .IN4(n81), .Q(
        \fpu_add_frac_dp/n4038 ) );
  AO221X1 U543 ( .IN1(n1591), .IN2(n612), .IN3(n1389), .IN4(n253), .IN5(n1592), 
        .Q(\fpu_add_frac_dp/n4037 ) );
  AO221X1 U544 ( .IN1(n1593), .IN2(n1594), .IN3(n1590), .IN4(n39), .IN5(n1595), 
        .Q(n1592) );
  AND2X1 U545 ( .IN1(n1596), .IN2(n1597), .Q(n1590) );
  NOR2X0 U546 ( .IN1(\fpu_add_frac_dp/n898 ), .IN2(n1598), .QN(n1593) );
  AO221X1 U547 ( .IN1(n1597), .IN2(n1599), .IN3(n1390), .IN4(n252), .IN5(n1600), .Q(\fpu_add_frac_dp/n4036 ) );
  AO221X1 U548 ( .IN1(n1601), .IN2(n612), .IN3(n1591), .IN4(n93), .IN5(n1595), 
        .Q(n1600) );
  AO221X1 U549 ( .IN1(n1597), .IN2(n1602), .IN3(n1392), .IN4(n327), .IN5(n1603), .Q(\fpu_add_frac_dp/n4035 ) );
  AO221X1 U550 ( .IN1(n1601), .IN2(n93), .IN3(n1591), .IN4(n182), .IN5(n1595), 
        .Q(n1603) );
  AO221X1 U551 ( .IN1(n1597), .IN2(n1604), .IN3(n1392), .IN4(n180), .IN5(n1605), .Q(\fpu_add_frac_dp/n4034 ) );
  AO221X1 U552 ( .IN1(n1601), .IN2(n182), .IN3(n1591), .IN4(n599), .IN5(n1595), 
        .Q(n1605) );
  AO221X1 U553 ( .IN1(n1597), .IN2(n1606), .IN3(n1392), .IN4(n268), .IN5(n1607), .Q(\fpu_add_frac_dp/n4033 ) );
  AO221X1 U554 ( .IN1(n1601), .IN2(n599), .IN3(n1591), .IN4(n183), .IN5(n1595), 
        .Q(n1607) );
  AO221X1 U555 ( .IN1(n1597), .IN2(n1608), .IN3(n1393), .IN4(n179), .IN5(n1609), .Q(\fpu_add_frac_dp/n4032 ) );
  AO221X1 U556 ( .IN1(n1601), .IN2(n183), .IN3(n1591), .IN4(n600), .IN5(n1595), 
        .Q(n1609) );
  AO221X1 U557 ( .IN1(n1597), .IN2(n1610), .IN3(n1393), .IN4(n251), .IN5(n1611), .Q(\fpu_add_frac_dp/n4031 ) );
  AO221X1 U558 ( .IN1(n1601), .IN2(n600), .IN3(n1591), .IN4(n184), .IN5(n1595), 
        .Q(n1611) );
  AO221X1 U559 ( .IN1(n1597), .IN2(n1612), .IN3(n1393), .IN4(n250), .IN5(n1613), .Q(\fpu_add_frac_dp/n4030 ) );
  AO221X1 U560 ( .IN1(n1601), .IN2(n184), .IN3(n1591), .IN4(n601), .IN5(n1595), 
        .Q(n1613) );
  AO221X1 U561 ( .IN1(n1597), .IN2(n1614), .IN3(n1393), .IN4(n249), .IN5(n1615), .Q(\fpu_add_frac_dp/n4029 ) );
  AO221X1 U562 ( .IN1(n1601), .IN2(n601), .IN3(n1591), .IN4(n185), .IN5(n1595), 
        .Q(n1615) );
  AO221X1 U563 ( .IN1(n1597), .IN2(n1616), .IN3(n1393), .IN4(n263), .IN5(n1617), .Q(\fpu_add_frac_dp/n4028 ) );
  AO221X1 U564 ( .IN1(n1601), .IN2(n185), .IN3(n1591), .IN4(n602), .IN5(n1595), 
        .Q(n1617) );
  AO221X1 U565 ( .IN1(n1597), .IN2(n1618), .IN3(n1393), .IN4(n267), .IN5(n1619), .Q(\fpu_add_frac_dp/n4027 ) );
  AO221X1 U566 ( .IN1(n1601), .IN2(n602), .IN3(n1591), .IN4(n186), .IN5(n1595), 
        .Q(n1619) );
  AO221X1 U567 ( .IN1(n1597), .IN2(n1620), .IN3(n1393), .IN4(n279), .IN5(n1621), .Q(\fpu_add_frac_dp/n4026 ) );
  AO221X1 U568 ( .IN1(n1601), .IN2(n186), .IN3(n1591), .IN4(n603), .IN5(n1595), 
        .Q(n1621) );
  AO221X1 U569 ( .IN1(n1597), .IN2(n1622), .IN3(n1393), .IN4(n318), .IN5(n1623), .Q(\fpu_add_frac_dp/n4025 ) );
  AO221X1 U570 ( .IN1(n1601), .IN2(n603), .IN3(n1591), .IN4(n187), .IN5(n1595), 
        .Q(n1623) );
  AO221X1 U571 ( .IN1(n1597), .IN2(n1624), .IN3(n1393), .IN4(n248), .IN5(n1625), .Q(\fpu_add_frac_dp/n4024 ) );
  AO221X1 U572 ( .IN1(n1601), .IN2(n187), .IN3(n1591), .IN4(n604), .IN5(n1595), 
        .Q(n1625) );
  AO221X1 U573 ( .IN1(n1597), .IN2(n1626), .IN3(n1394), .IN4(n247), .IN5(n1627), .Q(\fpu_add_frac_dp/n4023 ) );
  AO221X1 U574 ( .IN1(n1601), .IN2(n604), .IN3(n1591), .IN4(n188), .IN5(n1595), 
        .Q(n1627) );
  AO221X1 U575 ( .IN1(n1597), .IN2(n1628), .IN3(n1395), .IN4(n246), .IN5(n1629), .Q(\fpu_add_frac_dp/n4022 ) );
  AO221X1 U576 ( .IN1(n1601), .IN2(n188), .IN3(n1591), .IN4(n605), .IN5(n1595), 
        .Q(n1629) );
  AO221X1 U577 ( .IN1(n1597), .IN2(n1630), .IN3(n1389), .IN4(n204), .IN5(n1631), .Q(\fpu_add_frac_dp/n4021 ) );
  AO221X1 U578 ( .IN1(n1601), .IN2(n605), .IN3(n1591), .IN4(n189), .IN5(n1595), 
        .Q(n1631) );
  AO221X1 U579 ( .IN1(n1597), .IN2(n1632), .IN3(n1394), .IN4(n245), .IN5(n1633), .Q(\fpu_add_frac_dp/n4020 ) );
  AO221X1 U580 ( .IN1(n1601), .IN2(n189), .IN3(n1591), .IN4(n606), .IN5(n1595), 
        .Q(n1633) );
  AO221X1 U581 ( .IN1(n1597), .IN2(n1634), .IN3(n1394), .IN4(n244), .IN5(n1635), .Q(\fpu_add_frac_dp/n4019 ) );
  AO221X1 U582 ( .IN1(n1601), .IN2(n606), .IN3(n1591), .IN4(n190), .IN5(n1595), 
        .Q(n1635) );
  AO221X1 U583 ( .IN1(n1597), .IN2(n1636), .IN3(n1394), .IN4(n203), .IN5(n1637), .Q(\fpu_add_frac_dp/n4018 ) );
  AO221X1 U584 ( .IN1(n1601), .IN2(n190), .IN3(n1591), .IN4(n607), .IN5(n1595), 
        .Q(n1637) );
  AO221X1 U585 ( .IN1(n1597), .IN2(n1638), .IN3(n1394), .IN4(n243), .IN5(n1639), .Q(\fpu_add_frac_dp/n4017 ) );
  AO221X1 U586 ( .IN1(n1601), .IN2(n607), .IN3(n1591), .IN4(n191), .IN5(n1595), 
        .Q(n1639) );
  AO221X1 U587 ( .IN1(n1597), .IN2(n1640), .IN3(n1394), .IN4(n242), .IN5(n1641), .Q(\fpu_add_frac_dp/n4016 ) );
  AO221X1 U588 ( .IN1(n1601), .IN2(n191), .IN3(n1591), .IN4(n608), .IN5(n1595), 
        .Q(n1641) );
  AO221X1 U589 ( .IN1(n1597), .IN2(n1642), .IN3(n1394), .IN4(n241), .IN5(n1643), .Q(\fpu_add_frac_dp/n4015 ) );
  AO221X1 U590 ( .IN1(n1601), .IN2(n608), .IN3(n1591), .IN4(n192), .IN5(n1595), 
        .Q(n1643) );
  AO221X1 U591 ( .IN1(n1597), .IN2(n1644), .IN3(n1394), .IN4(n240), .IN5(n1645), .Q(\fpu_add_frac_dp/n4014 ) );
  AO221X1 U592 ( .IN1(n1601), .IN2(n192), .IN3(n1591), .IN4(n609), .IN5(n1595), 
        .Q(n1645) );
  AO221X1 U593 ( .IN1(n1597), .IN2(n1646), .IN3(n1394), .IN4(n202), .IN5(n1647), .Q(\fpu_add_frac_dp/n4013 ) );
  AO221X1 U594 ( .IN1(n1601), .IN2(n609), .IN3(n1591), .IN4(n193), .IN5(n1595), 
        .Q(n1647) );
  AO221X1 U595 ( .IN1(n1597), .IN2(n1648), .IN3(n1395), .IN4(n239), .IN5(n1649), .Q(\fpu_add_frac_dp/n4012 ) );
  AO221X1 U596 ( .IN1(n1601), .IN2(n193), .IN3(n1591), .IN4(n610), .IN5(n1595), 
        .Q(n1649) );
  AO221X1 U597 ( .IN1(n1597), .IN2(n1650), .IN3(n1395), .IN4(n201), .IN5(n1651), .Q(\fpu_add_frac_dp/n4011 ) );
  AO221X1 U598 ( .IN1(n1601), .IN2(n610), .IN3(n1591), .IN4(n194), .IN5(n1595), 
        .Q(n1651) );
  AO221X1 U599 ( .IN1(n1597), .IN2(n1652), .IN3(n1395), .IN4(n238), .IN5(n1653), .Q(\fpu_add_frac_dp/n4010 ) );
  AO221X1 U600 ( .IN1(n1601), .IN2(n194), .IN3(n1591), .IN4(n611), .IN5(n1595), 
        .Q(n1653) );
  AO221X1 U601 ( .IN1(n1597), .IN2(n1654), .IN3(n1395), .IN4(n200), .IN5(n1655), .Q(\fpu_add_frac_dp/n4009 ) );
  AO221X1 U602 ( .IN1(n1601), .IN2(n611), .IN3(n1591), .IN4(n207), .IN5(n1595), 
        .Q(n1655) );
  AND4X1 U603 ( .IN1(n1656), .IN2(n1657), .IN3(n1658), .IN4(n1659), .Q(n1595)
         );
  NAND4X0 U604 ( .IN1(n1660), .IN2(n1661), .IN3(n1662), .IN4(n1663), .QN(
        \fpu_add_frac_dp/n4008 ) );
  AOI222X1 U605 ( .IN1(n259), .IN2(n1422), .IN3(n644), .IN4(n1591), .IN5(n1664), .IN6(n1597), .QN(n1663) );
  NOR2X0 U606 ( .IN1(n1665), .IN2(n1666), .QN(n1591) );
  NAND2X0 U607 ( .IN1(n1601), .IN2(n207), .QN(n1662) );
  AND2X1 U608 ( .IN1(n1667), .IN2(n1668), .Q(n1601) );
  NAND3X0 U609 ( .IN1(n1668), .IN2(n176), .IN3(n1669), .QN(n1660) );
  AO221X1 U610 ( .IN1(n1597), .IN2(n1670), .IN3(n1395), .IN4(n237), .IN5(n1671), .Q(\fpu_add_frac_dp/n4007 ) );
  AO21X1 U611 ( .IN1(n1668), .IN2(n1672), .IN3(n1673), .Q(n1671) );
  AO221X1 U612 ( .IN1(n1597), .IN2(n1674), .IN3(n1394), .IN4(n199), .IN5(n1675), .Q(\fpu_add_frac_dp/n4006 ) );
  AO21X1 U613 ( .IN1(n1668), .IN2(n1676), .IN3(n1673), .Q(n1675) );
  AO221X1 U614 ( .IN1(n1597), .IN2(n1677), .IN3(n1395), .IN4(n236), .IN5(n1678), .Q(\fpu_add_frac_dp/n4005 ) );
  AO21X1 U615 ( .IN1(n1668), .IN2(n1679), .IN3(n1673), .Q(n1678) );
  AO221X1 U616 ( .IN1(n1597), .IN2(n1680), .IN3(n1395), .IN4(n235), .IN5(n1681), .Q(\fpu_add_frac_dp/n4004 ) );
  AO21X1 U617 ( .IN1(n1668), .IN2(n1682), .IN3(n1673), .Q(n1681) );
  AO221X1 U618 ( .IN1(n1597), .IN2(n1683), .IN3(n1395), .IN4(n234), .IN5(n1684), .Q(\fpu_add_frac_dp/n4003 ) );
  AO21X1 U619 ( .IN1(n1668), .IN2(n1685), .IN3(n1673), .Q(n1684) );
  AO221X1 U620 ( .IN1(n1597), .IN2(n1686), .IN3(n1395), .IN4(n198), .IN5(n1687), .Q(\fpu_add_frac_dp/n4002 ) );
  AO21X1 U621 ( .IN1(n1668), .IN2(n1688), .IN3(n1673), .Q(n1687) );
  AO221X1 U622 ( .IN1(n1597), .IN2(n1689), .IN3(n1396), .IN4(n197), .IN5(n1690), .Q(\fpu_add_frac_dp/n4001 ) );
  AO21X1 U623 ( .IN1(n1668), .IN2(n1691), .IN3(n1673), .Q(n1690) );
  AO221X1 U624 ( .IN1(n1597), .IN2(n1692), .IN3(n1396), .IN4(n233), .IN5(n1693), .Q(\fpu_add_frac_dp/n4000 ) );
  AO21X1 U625 ( .IN1(n1668), .IN2(n1694), .IN3(n1673), .Q(n1693) );
  AO221X1 U626 ( .IN1(n1597), .IN2(n1695), .IN3(n1395), .IN4(n232), .IN5(n1696), .Q(\fpu_add_frac_dp/n3999 ) );
  AO21X1 U627 ( .IN1(n1668), .IN2(n1697), .IN3(n1673), .Q(n1696) );
  AO221X1 U628 ( .IN1(n1597), .IN2(n1698), .IN3(n1396), .IN4(n231), .IN5(n1699), .Q(\fpu_add_frac_dp/n3998 ) );
  AO21X1 U629 ( .IN1(n1668), .IN2(n1700), .IN3(n1673), .Q(n1699) );
  AO221X1 U630 ( .IN1(n1597), .IN2(n1701), .IN3(n1394), .IN4(n230), .IN5(n1702), .Q(\fpu_add_frac_dp/n3997 ) );
  AO21X1 U631 ( .IN1(n1668), .IN2(n1703), .IN3(n1673), .Q(n1702) );
  AO221X1 U632 ( .IN1(n1597), .IN2(n1704), .IN3(n1396), .IN4(n229), .IN5(n1705), .Q(\fpu_add_frac_dp/n3996 ) );
  AO21X1 U633 ( .IN1(n1668), .IN2(n1706), .IN3(n1673), .Q(n1705) );
  AO221X1 U634 ( .IN1(n1597), .IN2(n1707), .IN3(n1394), .IN4(n228), .IN5(n1708), .Q(\fpu_add_frac_dp/n3995 ) );
  AO21X1 U635 ( .IN1(n1668), .IN2(n1709), .IN3(n1673), .Q(n1708) );
  AO221X1 U636 ( .IN1(n1597), .IN2(n1710), .IN3(n1396), .IN4(n227), .IN5(n1711), .Q(\fpu_add_frac_dp/n3994 ) );
  AO21X1 U637 ( .IN1(n1668), .IN2(n1712), .IN3(n1673), .Q(n1711) );
  AO221X1 U638 ( .IN1(n1597), .IN2(n1713), .IN3(n1394), .IN4(n196), .IN5(n1714), .Q(\fpu_add_frac_dp/n3993 ) );
  AO21X1 U639 ( .IN1(n1668), .IN2(n1715), .IN3(n1673), .Q(n1714) );
  AO221X1 U640 ( .IN1(n1597), .IN2(n1716), .IN3(n1396), .IN4(n294), .IN5(n1717), .Q(\fpu_add_frac_dp/n3992 ) );
  AO21X1 U641 ( .IN1(n1668), .IN2(n1718), .IN3(n1673), .Q(n1717) );
  AO221X1 U642 ( .IN1(n1597), .IN2(n1719), .IN3(n1395), .IN4(n332), .IN5(n1720), .Q(\fpu_add_frac_dp/n3991 ) );
  AO21X1 U643 ( .IN1(n1668), .IN2(n1721), .IN3(n1673), .Q(n1720) );
  AO221X1 U644 ( .IN1(n1597), .IN2(n1722), .IN3(n1396), .IN4(n334), .IN5(n1723), .Q(\fpu_add_frac_dp/n3990 ) );
  AO21X1 U645 ( .IN1(n1668), .IN2(n1724), .IN3(n1673), .Q(n1723) );
  AO221X1 U646 ( .IN1(n1597), .IN2(n1725), .IN3(n1395), .IN4(n293), .IN5(n1726), .Q(\fpu_add_frac_dp/n3989 ) );
  AO21X1 U647 ( .IN1(n1668), .IN2(n1727), .IN3(n1673), .Q(n1726) );
  AO221X1 U648 ( .IN1(n1597), .IN2(n1728), .IN3(n1396), .IN4(n317), .IN5(n1729), .Q(\fpu_add_frac_dp/n3988 ) );
  AO21X1 U649 ( .IN1(n1668), .IN2(n1730), .IN3(n1673), .Q(n1729) );
  AO221X1 U650 ( .IN1(n1597), .IN2(n1731), .IN3(n1395), .IN4(n195), .IN5(n1732), .Q(\fpu_add_frac_dp/n3987 ) );
  AO21X1 U651 ( .IN1(n1668), .IN2(n1733), .IN3(n1673), .Q(n1732) );
  AO221X1 U652 ( .IN1(n1597), .IN2(n1734), .IN3(n1396), .IN4(n226), .IN5(n1735), .Q(\fpu_add_frac_dp/n3986 ) );
  AO221X1 U653 ( .IN1(n1736), .IN2(n1737), .IN3(n1668), .IN4(n1738), .IN5(
        n1673), .Q(n1735) );
  INVX0 U654 ( .INP(n1661), .ZN(n1673) );
  NAND2X0 U655 ( .IN1(n1739), .IN2(n1659), .QN(n1661) );
  INVX0 U656 ( .INP(n1740), .ZN(n1739) );
  AND2X1 U657 ( .IN1(n1741), .IN2(n1659), .Q(n1736) );
  NAND2X0 U658 ( .IN1(n1598), .IN2(n1666), .QN(n1659) );
  AO222X1 U659 ( .IN1(n1597), .IN2(n1742), .IN3(n1668), .IN4(n1743), .IN5(
        n1384), .IN6(n850), .Q(\fpu_add_frac_dp/n3985 ) );
  INVX0 U660 ( .INP(n1666), .ZN(n1668) );
  AO21X1 U661 ( .IN1(n1737), .IN2(n1744), .IN3(n1745), .Q(n1666) );
  NAND3X0 U662 ( .IN1(n1435), .IN2(n1744), .IN3(n1737), .QN(n1598) );
  AO221X1 U663 ( .IN1(n1747), .IN2(n1748), .IN3(n1749), .IN4(n1750), .IN5(
        n1751), .Q(n1744) );
  OR2X1 U664 ( .IN1(n1752), .IN2(n1753), .Q(n1747) );
  AO22X1 U665 ( .IN1(n1419), .IN2(n1196), .IN3(n1754), .IN4(n36), .Q(
        \fpu_add_frac_dp/n3984 ) );
  AO22X1 U666 ( .IN1(n1419), .IN2(n1134), .IN3(n1754), .IN4(n170), .Q(
        \fpu_add_frac_dp/n3983 ) );
  AO22X1 U667 ( .IN1(n1419), .IN2(n1135), .IN3(n1754), .IN4(n10), .Q(
        \fpu_add_frac_dp/n3982 ) );
  AO22X1 U668 ( .IN1(n1419), .IN2(n1136), .IN3(n1754), .IN4(n1589), .Q(
        \fpu_add_frac_dp/n3981 ) );
  AO22X1 U669 ( .IN1(n1419), .IN2(n1137), .IN3(n1754), .IN4(n11), .Q(
        \fpu_add_frac_dp/n3980 ) );
  AO22X1 U670 ( .IN1(n1419), .IN2(n1149), .IN3(n1754), .IN4(n30), .Q(
        \fpu_add_frac_dp/n3979 ) );
  AO22X1 U671 ( .IN1(n1419), .IN2(n1138), .IN3(n1754), .IN4(n79), .Q(
        \fpu_add_frac_dp/n3978 ) );
  AO22X1 U672 ( .IN1(n1419), .IN2(n1139), .IN3(n1754), .IN4(n31), .Q(
        \fpu_add_frac_dp/n3977 ) );
  AO22X1 U673 ( .IN1(n1418), .IN2(n1140), .IN3(n1754), .IN4(n80), .Q(
        \fpu_add_frac_dp/n3976 ) );
  AO22X1 U674 ( .IN1(n1418), .IN2(n1141), .IN3(n1754), .IN4(n32), .Q(
        \fpu_add_frac_dp/n3975 ) );
  AO22X1 U675 ( .IN1(n1418), .IN2(n1142), .IN3(n1754), .IN4(n81), .Q(
        \fpu_add_frac_dp/n3974 ) );
  AO21X1 U676 ( .IN1(n1397), .IN2(n1111), .IN3(n1755), .Q(
        \fpu_add_frac_dp/n3973 ) );
  AO21X1 U677 ( .IN1(\fpu_add_frac_dp/n2389 ), .IN2(n1415), .IN3(n1756), .Q(
        \fpu_add_frac_dp/n3972 ) );
  AO21X1 U678 ( .IN1(n1398), .IN2(n1091), .IN3(n1757), .Q(
        \fpu_add_frac_dp/n3971 ) );
  AO21X1 U679 ( .IN1(n1398), .IN2(n1122), .IN3(n1758), .Q(
        \fpu_add_frac_dp/n3970 ) );
  AO21X1 U680 ( .IN1(n1398), .IN2(n1125), .IN3(n1759), .Q(
        \fpu_add_frac_dp/n3969 ) );
  AO21X1 U681 ( .IN1(n1398), .IN2(n1123), .IN3(n1760), .Q(
        \fpu_add_frac_dp/n3968 ) );
  AO21X1 U682 ( .IN1(n1398), .IN2(n722), .IN3(n1761), .Q(
        \fpu_add_frac_dp/n3967 ) );
  AO21X1 U683 ( .IN1(n1398), .IN2(n423), .IN3(n1762), .Q(
        \fpu_add_frac_dp/n3966 ) );
  AO21X1 U684 ( .IN1(n1398), .IN2(n1104), .IN3(n1763), .Q(
        \fpu_add_frac_dp/n3965 ) );
  AO21X1 U685 ( .IN1(n1398), .IN2(n1092), .IN3(n1764), .Q(
        \fpu_add_frac_dp/n3964 ) );
  AO21X1 U686 ( .IN1(n1398), .IN2(n1112), .IN3(n1765), .Q(
        \fpu_add_frac_dp/n3963 ) );
  AO21X1 U687 ( .IN1(n1398), .IN2(n724), .IN3(n1766), .Q(
        \fpu_add_frac_dp/n3962 ) );
  AO21X1 U688 ( .IN1(n1398), .IN2(n426), .IN3(n1767), .Q(
        \fpu_add_frac_dp/n3961 ) );
  AO21X1 U689 ( .IN1(n1398), .IN2(n1105), .IN3(n1768), .Q(
        \fpu_add_frac_dp/n3960 ) );
  AO21X1 U690 ( .IN1(n1398), .IN2(n1093), .IN3(n1769), .Q(
        \fpu_add_frac_dp/n3959 ) );
  AO21X1 U691 ( .IN1(n1398), .IN2(n1113), .IN3(n1770), .Q(
        \fpu_add_frac_dp/n3958 ) );
  AO21X1 U692 ( .IN1(n1399), .IN2(n723), .IN3(n1771), .Q(
        \fpu_add_frac_dp/n3957 ) );
  AO21X1 U693 ( .IN1(n1399), .IN2(n424), .IN3(n1772), .Q(
        \fpu_add_frac_dp/n3956 ) );
  AO21X1 U694 ( .IN1(n1399), .IN2(n1106), .IN3(n1773), .Q(
        \fpu_add_frac_dp/n3955 ) );
  AO21X1 U695 ( .IN1(n1399), .IN2(n1094), .IN3(n1774), .Q(
        \fpu_add_frac_dp/n3954 ) );
  AO21X1 U696 ( .IN1(n1399), .IN2(n1114), .IN3(n1775), .Q(
        \fpu_add_frac_dp/n3953 ) );
  AO21X1 U697 ( .IN1(n1399), .IN2(n1107), .IN3(n1776), .Q(
        \fpu_add_frac_dp/n3952 ) );
  AO21X1 U698 ( .IN1(n1399), .IN2(n1095), .IN3(n1777), .Q(
        \fpu_add_frac_dp/n3951 ) );
  AO21X1 U699 ( .IN1(n1399), .IN2(n1096), .IN3(n1778), .Q(
        \fpu_add_frac_dp/n3950 ) );
  AO21X1 U700 ( .IN1(n1399), .IN2(n1115), .IN3(n1779), .Q(
        \fpu_add_frac_dp/n3949 ) );
  AO21X1 U701 ( .IN1(n1399), .IN2(n1108), .IN3(n1780), .Q(
        \fpu_add_frac_dp/n3948 ) );
  AO21X1 U702 ( .IN1(n1399), .IN2(n1097), .IN3(n1781), .Q(
        \fpu_add_frac_dp/n3947 ) );
  AO21X1 U703 ( .IN1(n1399), .IN2(n1098), .IN3(n1782), .Q(
        \fpu_add_frac_dp/n3946 ) );
  AO21X1 U704 ( .IN1(n1399), .IN2(n1116), .IN3(n1783), .Q(
        \fpu_add_frac_dp/n3945 ) );
  AO21X1 U705 ( .IN1(n1400), .IN2(n1109), .IN3(n1784), .Q(
        \fpu_add_frac_dp/n3944 ) );
  AO21X1 U706 ( .IN1(n1400), .IN2(n1099), .IN3(n1785), .Q(
        \fpu_add_frac_dp/n3943 ) );
  AO21X1 U707 ( .IN1(n1400), .IN2(n1102), .IN3(n1786), .Q(
        \fpu_add_frac_dp/n3942 ) );
  AO21X1 U708 ( .IN1(n1400), .IN2(n1117), .IN3(n1787), .Q(
        \fpu_add_frac_dp/n3941 ) );
  AO21X1 U709 ( .IN1(n1400), .IN2(n58), .IN3(n1788), .Q(
        \fpu_add_frac_dp/n3940 ) );
  AO21X1 U710 ( .IN1(n1400), .IN2(n143), .IN3(n1789), .Q(
        \fpu_add_frac_dp/n3939 ) );
  AO21X1 U711 ( .IN1(n1400), .IN2(n344), .IN3(n1790), .Q(
        \fpu_add_frac_dp/n3938 ) );
  AO21X1 U712 ( .IN1(n1396), .IN2(n707), .IN3(n1791), .Q(
        \fpu_add_frac_dp/n3937 ) );
  AO21X1 U713 ( .IN1(n1404), .IN2(n59), .IN3(n1792), .Q(
        \fpu_add_frac_dp/n3936 ) );
  AO21X1 U714 ( .IN1(n1404), .IN2(n144), .IN3(n1793), .Q(
        \fpu_add_frac_dp/n3935 ) );
  AO21X1 U715 ( .IN1(n1404), .IN2(n345), .IN3(n1794), .Q(
        \fpu_add_frac_dp/n3934 ) );
  AO21X1 U716 ( .IN1(n1404), .IN2(n708), .IN3(n1795), .Q(
        \fpu_add_frac_dp/n3933 ) );
  AO21X1 U717 ( .IN1(n1404), .IN2(n1110), .IN3(n1796), .Q(
        \fpu_add_frac_dp/n3932 ) );
  AO21X1 U718 ( .IN1(n1403), .IN2(n1100), .IN3(n1797), .Q(
        \fpu_add_frac_dp/n3931 ) );
  AO21X1 U719 ( .IN1(n1403), .IN2(n1103), .IN3(n1798), .Q(
        \fpu_add_frac_dp/n3930 ) );
  AO21X1 U720 ( .IN1(n1403), .IN2(n1118), .IN3(n1799), .Q(
        \fpu_add_frac_dp/n3929 ) );
  AO21X1 U721 ( .IN1(n1403), .IN2(n343), .IN3(n1800), .Q(
        \fpu_add_frac_dp/n3928 ) );
  AO21X1 U722 ( .IN1(\fpu_add_frac_dp/n2392 ), .IN2(n1415), .IN3(n1801), .Q(
        \fpu_add_frac_dp/n3927 ) );
  AO21X1 U723 ( .IN1(\fpu_add_frac_dp/n2390 ), .IN2(n1415), .IN3(n1802), .Q(
        \fpu_add_frac_dp/n3926 ) );
  AO21X1 U724 ( .IN1(\fpu_add_frac_dp/n2391 ), .IN2(n1415), .IN3(n1803), .Q(
        \fpu_add_frac_dp/n3925 ) );
  AO21X1 U725 ( .IN1(\fpu_add_frac_dp/n2384 ), .IN2(n1415), .IN3(n1804), .Q(
        \fpu_add_frac_dp/n3924 ) );
  AO21X1 U726 ( .IN1(n1403), .IN2(n706), .IN3(n1805), .Q(
        \fpu_add_frac_dp/n3923 ) );
  AO21X1 U727 ( .IN1(n1403), .IN2(n142), .IN3(n1806), .Q(
        \fpu_add_frac_dp/n3922 ) );
  AO21X1 U728 ( .IN1(n1403), .IN2(n1101), .IN3(n1807), .Q(
        \fpu_add_frac_dp/n3921 ) );
  AO22X1 U729 ( .IN1(n1428), .IN2(n896), .IN3(n1754), .IN4(n36), .Q(
        \fpu_add_frac_dp/n3920 ) );
  AO22X1 U730 ( .IN1(n1430), .IN2(n902), .IN3(n1754), .IN4(n170), .Q(
        \fpu_add_frac_dp/n3919 ) );
  AO22X1 U731 ( .IN1(n1429), .IN2(n690), .IN3(n1754), .IN4(n10), .Q(
        \fpu_add_frac_dp/n3918 ) );
  AO22X1 U732 ( .IN1(n1430), .IN2(n899), .IN3(n1754), .IN4(n1589), .Q(
        \fpu_add_frac_dp/n3917 ) );
  AO22X1 U733 ( .IN1(n1429), .IN2(n660), .IN3(n1754), .IN4(n11), .Q(
        \fpu_add_frac_dp/n3916 ) );
  AO22X1 U734 ( .IN1(n1429), .IN2(n898), .IN3(n1754), .IN4(n30), .Q(
        \fpu_add_frac_dp/n3915 ) );
  AO22X1 U735 ( .IN1(n1428), .IN2(n655), .IN3(n1754), .IN4(n79), .Q(
        \fpu_add_frac_dp/n3914 ) );
  AO22X1 U736 ( .IN1(n1429), .IN2(n901), .IN3(n1754), .IN4(n31), .Q(
        \fpu_add_frac_dp/n3913 ) );
  AO22X1 U737 ( .IN1(n1429), .IN2(n659), .IN3(n1754), .IN4(n80), .Q(
        \fpu_add_frac_dp/n3912 ) );
  AO22X1 U738 ( .IN1(n1429), .IN2(n75), .IN3(n1754), .IN4(n32), .Q(
        \fpu_add_frac_dp/n3911 ) );
  AO22X1 U739 ( .IN1(n1429), .IN2(n161), .IN3(n1754), .IN4(n81), .Q(
        \fpu_add_frac_dp/n3910 ) );
  AO21X1 U740 ( .IN1(n1403), .IN2(n627), .IN3(n1755), .Q(
        \fpu_add_frac_dp/n3909 ) );
  AO222X1 U741 ( .IN1(n1754), .IN2(n39), .IN3(n1808), .IN4(n1809), .IN5(n1810), 
        .IN6(n612), .Q(n1755) );
  NOR2X0 U742 ( .IN1(\fpu_add_frac_dp/n898 ), .IN2(n1811), .QN(n1808) );
  AND2X1 U743 ( .IN1(n1809), .IN2(n1596), .Q(n1754) );
  AO21X1 U744 ( .IN1(n1403), .IN2(n150), .IN3(n1756), .Q(
        \fpu_add_frac_dp/n3908 ) );
  AO222X1 U745 ( .IN1(n1810), .IN2(n93), .IN3(n1809), .IN4(n1599), .IN5(n1812), 
        .IN6(n612), .Q(n1756) );
  AO222X1 U746 ( .IN1(n1813), .IN2(n36), .IN3(n1596), .IN4(n120), .IN5(n1594), 
        .IN6(n170), .Q(n1599) );
  AO21X1 U747 ( .IN1(n1403), .IN2(n721), .IN3(n1757), .Q(
        \fpu_add_frac_dp/n3907 ) );
  AO222X1 U748 ( .IN1(n1810), .IN2(n182), .IN3(n1809), .IN4(n1602), .IN5(n1812), .IN6(n93), .Q(n1757) );
  AO222X1 U749 ( .IN1(n1813), .IN2(n170), .IN3(n1596), .IN4(n52), .IN5(n1594), 
        .IN6(n10), .Q(n1602) );
  AO21X1 U750 ( .IN1(n1403), .IN2(n425), .IN3(n1758), .Q(
        \fpu_add_frac_dp/n3906 ) );
  AO222X1 U751 ( .IN1(n1810), .IN2(n599), .IN3(n1809), .IN4(n1604), .IN5(n1812), .IN6(n182), .Q(n1758) );
  AO222X1 U752 ( .IN1(n1813), .IN2(n10), .IN3(n1596), .IN4(n121), .IN5(n1594), 
        .IN6(n1589), .Q(n1604) );
  AO21X1 U753 ( .IN1(n1403), .IN2(n935), .IN3(n1759), .Q(
        \fpu_add_frac_dp/n3905 ) );
  AO222X1 U754 ( .IN1(n1810), .IN2(n183), .IN3(n1809), .IN4(n1606), .IN5(n1812), .IN6(n599), .Q(n1759) );
  AO222X1 U755 ( .IN1(n1813), .IN2(n1589), .IN3(n1596), .IN4(n53), .IN5(n1594), 
        .IN6(n11), .Q(n1606) );
  INVX0 U756 ( .INP(\fpu_add_frac_dp/n895 ), .ZN(n1589) );
  AO21X1 U757 ( .IN1(n1403), .IN2(n930), .IN3(n1760), .Q(
        \fpu_add_frac_dp/n3904 ) );
  AO222X1 U758 ( .IN1(n1810), .IN2(n600), .IN3(n1809), .IN4(n1608), .IN5(n1812), .IN6(n183), .Q(n1760) );
  AO222X1 U759 ( .IN1(n1813), .IN2(n11), .IN3(n1596), .IN4(n122), .IN5(n1594), 
        .IN6(n30), .Q(n1608) );
  AO21X1 U760 ( .IN1(n1403), .IN2(n1151), .IN3(n1761), .Q(
        \fpu_add_frac_dp/n3903 ) );
  AO222X1 U761 ( .IN1(n1810), .IN2(n184), .IN3(n1809), .IN4(n1610), .IN5(n1812), .IN6(n600), .Q(n1761) );
  AO222X1 U762 ( .IN1(n1813), .IN2(n30), .IN3(n1596), .IN4(n272), .IN5(n1594), 
        .IN6(n79), .Q(n1610) );
  AO21X1 U763 ( .IN1(n1402), .IN2(n1152), .IN3(n1762), .Q(
        \fpu_add_frac_dp/n3902 ) );
  AO222X1 U764 ( .IN1(n1810), .IN2(n601), .IN3(n1809), .IN4(n1612), .IN5(n1812), .IN6(n184), .Q(n1762) );
  AO222X1 U765 ( .IN1(n1813), .IN2(n79), .IN3(n1596), .IN4(n633), .IN5(n1594), 
        .IN6(n31), .Q(n1612) );
  AO21X1 U766 ( .IN1(n1402), .IN2(n717), .IN3(n1763), .Q(
        \fpu_add_frac_dp/n3901 ) );
  AO222X1 U767 ( .IN1(n1810), .IN2(n185), .IN3(n1809), .IN4(n1614), .IN5(n1812), .IN6(n601), .Q(n1763) );
  AO222X1 U768 ( .IN1(n1813), .IN2(n31), .IN3(n1596), .IN4(n273), .IN5(n1594), 
        .IN6(n80), .Q(n1614) );
  AO21X1 U769 ( .IN1(n1402), .IN2(n314), .IN3(n1764), .Q(
        \fpu_add_frac_dp/n3900 ) );
  AO222X1 U770 ( .IN1(n1810), .IN2(n602), .IN3(n1809), .IN4(n1616), .IN5(n1812), .IN6(n185), .Q(n1764) );
  AO222X1 U771 ( .IN1(n1813), .IN2(n80), .IN3(n1596), .IN4(n634), .IN5(n1594), 
        .IN6(n32), .Q(n1616) );
  AO21X1 U772 ( .IN1(n1402), .IN2(n131), .IN3(n1765), .Q(
        \fpu_add_frac_dp/n3899 ) );
  AO222X1 U773 ( .IN1(n1810), .IN2(n186), .IN3(n1809), .IN4(n1618), .IN5(n1812), .IN6(n602), .Q(n1765) );
  AO222X1 U774 ( .IN1(n1813), .IN2(n32), .IN3(n1596), .IN4(n274), .IN5(n1594), 
        .IN6(n81), .Q(n1618) );
  AO21X1 U775 ( .IN1(n1402), .IN2(n934), .IN3(n1766), .Q(
        \fpu_add_frac_dp/n3898 ) );
  AO222X1 U776 ( .IN1(n1810), .IN2(n603), .IN3(n1809), .IN4(n1620), .IN5(n1812), .IN6(n186), .Q(n1766) );
  AO222X1 U777 ( .IN1(n1813), .IN2(n81), .IN3(n1596), .IN4(n635), .IN5(n1594), 
        .IN6(n39), .Q(n1620) );
  AO21X1 U778 ( .IN1(n1402), .IN2(n931), .IN3(n1767), .Q(
        \fpu_add_frac_dp/n3897 ) );
  AO222X1 U779 ( .IN1(n1810), .IN2(n187), .IN3(n1809), .IN4(n1622), .IN5(n1812), .IN6(n603), .Q(n1767) );
  AO222X1 U780 ( .IN1(n1813), .IN2(n39), .IN3(n1596), .IN4(n275), .IN5(n1594), 
        .IN6(n120), .Q(n1622) );
  AO21X1 U781 ( .IN1(n1402), .IN2(n929), .IN3(n1768), .Q(
        \fpu_add_frac_dp/n3896 ) );
  AO222X1 U782 ( .IN1(n1810), .IN2(n604), .IN3(n1809), .IN4(n1624), .IN5(n1812), .IN6(n187), .Q(n1768) );
  AO222X1 U783 ( .IN1(n1813), .IN2(n120), .IN3(n1596), .IN4(n636), .IN5(n1594), 
        .IN6(n52), .Q(n1624) );
  AO21X1 U784 ( .IN1(n1402), .IN2(n932), .IN3(n1769), .Q(
        \fpu_add_frac_dp/n3895 ) );
  AO222X1 U785 ( .IN1(n1810), .IN2(n188), .IN3(n1809), .IN4(n1626), .IN5(n1812), .IN6(n604), .Q(n1769) );
  AO222X1 U786 ( .IN1(n1813), .IN2(n52), .IN3(n1596), .IN4(n276), .IN5(n1594), 
        .IN6(n121), .Q(n1626) );
  AO21X1 U787 ( .IN1(n1402), .IN2(n312), .IN3(n1770), .Q(
        \fpu_add_frac_dp/n3894 ) );
  AO222X1 U788 ( .IN1(n1810), .IN2(n605), .IN3(n1809), .IN4(n1628), .IN5(n1812), .IN6(n188), .Q(n1770) );
  AO222X1 U789 ( .IN1(n1813), .IN2(n121), .IN3(n1596), .IN4(n637), .IN5(n1594), 
        .IN6(n53), .Q(n1628) );
  AO21X1 U790 ( .IN1(n1402), .IN2(n720), .IN3(n1771), .Q(
        \fpu_add_frac_dp/n3893 ) );
  AO222X1 U791 ( .IN1(n1810), .IN2(n189), .IN3(n1809), .IN4(n1630), .IN5(n1812), .IN6(n605), .Q(n1771) );
  AO222X1 U792 ( .IN1(n1813), .IN2(n53), .IN3(n1596), .IN4(n277), .IN5(n1594), 
        .IN6(n122), .Q(n1630) );
  AO21X1 U793 ( .IN1(n1402), .IN2(n106), .IN3(n1772), .Q(
        \fpu_add_frac_dp/n3892 ) );
  AO222X1 U794 ( .IN1(n1810), .IN2(n606), .IN3(n1809), .IN4(n1632), .IN5(n1812), .IN6(n189), .Q(n1772) );
  AO222X1 U795 ( .IN1(n1813), .IN2(n122), .IN3(n1596), .IN4(n639), .IN5(n1594), 
        .IN6(n272), .Q(n1632) );
  AO21X1 U796 ( .IN1(n1402), .IN2(n679), .IN3(n1773), .Q(
        \fpu_add_frac_dp/n3891 ) );
  AO222X1 U797 ( .IN1(n1810), .IN2(n190), .IN3(n1809), .IN4(n1634), .IN5(n1812), .IN6(n606), .Q(n1773) );
  AO222X1 U798 ( .IN1(n1813), .IN2(n272), .IN3(n1596), .IN4(n112), .IN5(n1594), 
        .IN6(n633), .Q(n1634) );
  AO21X1 U799 ( .IN1(n1402), .IN2(n678), .IN3(n1774), .Q(
        \fpu_add_frac_dp/n3890 ) );
  AO222X1 U800 ( .IN1(n1810), .IN2(n607), .IN3(n1809), .IN4(n1636), .IN5(n1812), .IN6(n190), .Q(n1774) );
  AO222X1 U801 ( .IN1(n1813), .IN2(n633), .IN3(n1596), .IN4(n113), .IN5(n1594), 
        .IN6(n273), .Q(n1636) );
  AO21X1 U802 ( .IN1(n1402), .IN2(n696), .IN3(n1775), .Q(
        \fpu_add_frac_dp/n3889 ) );
  AO222X1 U803 ( .IN1(n1810), .IN2(n191), .IN3(n1809), .IN4(n1638), .IN5(n1812), .IN6(n607), .Q(n1775) );
  AO222X1 U804 ( .IN1(n1813), .IN2(n273), .IN3(n1596), .IN4(n114), .IN5(n1594), 
        .IN6(n634), .Q(n1638) );
  AO21X1 U805 ( .IN1(n1401), .IN2(n218), .IN3(n1776), .Q(
        \fpu_add_frac_dp/n3888 ) );
  AO222X1 U806 ( .IN1(n1810), .IN2(n608), .IN3(n1809), .IN4(n1640), .IN5(n1812), .IN6(n191), .Q(n1776) );
  AO222X1 U807 ( .IN1(n1813), .IN2(n634), .IN3(n1596), .IN4(n7), .IN5(n1594), 
        .IN6(n274), .Q(n1640) );
  AO21X1 U808 ( .IN1(n1399), .IN2(n278), .IN3(n1777), .Q(
        \fpu_add_frac_dp/n3887 ) );
  AO222X1 U809 ( .IN1(n1810), .IN2(n192), .IN3(n1809), .IN4(n1642), .IN5(n1812), .IN6(n608), .Q(n1777) );
  AO222X1 U810 ( .IN1(n1813), .IN2(n274), .IN3(n1596), .IN4(n8), .IN5(n1594), 
        .IN6(n635), .Q(n1642) );
  AO21X1 U811 ( .IN1(\fpu_add_frac_dp/n2393 ), .IN2(n1415), .IN3(n1778), .Q(
        \fpu_add_frac_dp/n3886 ) );
  AO222X1 U812 ( .IN1(n1810), .IN2(n609), .IN3(n1809), .IN4(n1644), .IN5(n1812), .IN6(n192), .Q(n1778) );
  AO222X1 U813 ( .IN1(n1813), .IN2(n635), .IN3(n1596), .IN4(n9), .IN5(n1594), 
        .IN6(n275), .Q(n1644) );
  AO21X1 U814 ( .IN1(n1401), .IN2(n205), .IN3(n1779), .Q(
        \fpu_add_frac_dp/n3885 ) );
  AO222X1 U815 ( .IN1(n1810), .IN2(n193), .IN3(n1809), .IN4(n1646), .IN5(n1812), .IN6(n609), .Q(n1779) );
  AO222X1 U816 ( .IN1(n1813), .IN2(n275), .IN3(n1596), .IN4(n24), .IN5(n1594), 
        .IN6(n636), .Q(n1646) );
  AO21X1 U817 ( .IN1(n1401), .IN2(n6), .IN3(n1780), .Q(\fpu_add_frac_dp/n3884 ) );
  AO222X1 U818 ( .IN1(n1810), .IN2(n610), .IN3(n1809), .IN4(n1648), .IN5(n1812), .IN6(n193), .Q(n1780) );
  AO222X1 U819 ( .IN1(n1813), .IN2(n636), .IN3(n1596), .IN4(n25), .IN5(n1594), 
        .IN6(n276), .Q(n1648) );
  AO21X1 U820 ( .IN1(n1401), .IN2(n162), .IN3(n1781), .Q(
        \fpu_add_frac_dp/n3883 ) );
  AO222X1 U821 ( .IN1(n1810), .IN2(n194), .IN3(n1809), .IN4(n1650), .IN5(n1812), .IN6(n610), .Q(n1781) );
  AO222X1 U822 ( .IN1(n1813), .IN2(n276), .IN3(n1596), .IN4(n26), .IN5(n1594), 
        .IN6(n637), .Q(n1650) );
  AO21X1 U823 ( .IN1(n1401), .IN2(n23), .IN3(n1782), .Q(
        \fpu_add_frac_dp/n3882 ) );
  AO222X1 U824 ( .IN1(n1810), .IN2(n611), .IN3(n1809), .IN4(n1652), .IN5(n1812), .IN6(n194), .Q(n1782) );
  AO222X1 U825 ( .IN1(n1813), .IN2(n637), .IN3(n1596), .IN4(n76), .IN5(n1594), 
        .IN6(n277), .Q(n1652) );
  AO21X1 U826 ( .IN1(n1401), .IN2(n271), .IN3(n1783), .Q(
        \fpu_add_frac_dp/n3881 ) );
  AO222X1 U827 ( .IN1(n1810), .IN2(n207), .IN3(n1809), .IN4(n1654), .IN5(n1812), .IN6(n611), .Q(n1783) );
  AO222X1 U828 ( .IN1(n1813), .IN2(n277), .IN3(n1596), .IN4(n77), .IN5(n1594), 
        .IN6(n639), .Q(n1654) );
  AO21X1 U829 ( .IN1(n1401), .IN2(n168), .IN3(n1784), .Q(
        \fpu_add_frac_dp/n3880 ) );
  AO221X1 U830 ( .IN1(n1810), .IN2(n644), .IN3(n1812), .IN4(n207), .IN5(n1814), 
        .Q(n1784) );
  AO22X1 U831 ( .IN1(n1809), .IN2(n1664), .IN3(n1815), .IN4(n1816), .Q(n1814)
         );
  NOR2X0 U832 ( .IN1(\fpu_add_frac_dp/n965 ), .IN2(n1817), .QN(n1815) );
  AO221X1 U833 ( .IN1(n1818), .IN2(n7), .IN3(n1594), .IN4(n112), .IN5(n1819), 
        .Q(n1664) );
  AO22X1 U834 ( .IN1(n1813), .IN2(n639), .IN3(n1596), .IN4(n167), .Q(n1819) );
  AND2X1 U835 ( .IN1(n1816), .IN2(n1667), .Q(n1812) );
  AND2X1 U836 ( .IN1(n1816), .IN2(n1820), .Q(n1810) );
  AO21X1 U837 ( .IN1(\fpu_add_frac_dp/n2380 ), .IN2(n1415), .IN3(n1785), .Q(
        \fpu_add_frac_dp/n3879 ) );
  AO22X1 U838 ( .IN1(n1809), .IN2(n1670), .IN3(n1816), .IN4(n1672), .Q(n1785)
         );
  AO221X1 U839 ( .IN1(n1669), .IN2(n208), .IN3(n1820), .IN4(n698), .IN5(n1821), 
        .Q(n1672) );
  AO22X1 U840 ( .IN1(n1667), .IN2(n644), .IN3(n1822), .IN4(n176), .Q(n1821) );
  AO221X1 U841 ( .IN1(n1818), .IN2(n8), .IN3(n1594), .IN4(n113), .IN5(n1823), 
        .Q(n1670) );
  AO222X1 U842 ( .IN1(n1824), .IN2(n7), .IN3(n1596), .IN4(n27), .IN5(n1813), 
        .IN6(n112), .Q(n1823) );
  AO21X1 U843 ( .IN1(n1401), .IN2(n70), .IN3(n1786), .Q(
        \fpu_add_frac_dp/n3878 ) );
  AO22X1 U844 ( .IN1(n1809), .IN2(n1674), .IN3(n1816), .IN4(n1676), .Q(n1786)
         );
  AO221X1 U845 ( .IN1(n1669), .IN2(n99), .IN3(n1820), .IN4(n699), .IN5(n1825), 
        .Q(n1676) );
  AO22X1 U846 ( .IN1(n1667), .IN2(n698), .IN3(n1822), .IN4(n208), .Q(n1825) );
  AO221X1 U847 ( .IN1(n1818), .IN2(n9), .IN3(n1594), .IN4(n114), .IN5(n1826), 
        .Q(n1674) );
  AO222X1 U848 ( .IN1(n1824), .IN2(n8), .IN3(n1596), .IN4(n28), .IN5(n1813), 
        .IN6(n113), .Q(n1826) );
  AO21X1 U849 ( .IN1(n1401), .IN2(n174), .IN3(n1787), .Q(
        \fpu_add_frac_dp/n3877 ) );
  AO22X1 U850 ( .IN1(n1809), .IN2(n1677), .IN3(n1816), .IN4(n1679), .Q(n1787)
         );
  AO221X1 U851 ( .IN1(n1669), .IN2(n614), .IN3(n1820), .IN4(n176), .IN5(n1827), 
        .Q(n1679) );
  AO22X1 U852 ( .IN1(n1667), .IN2(n699), .IN3(n1822), .IN4(n99), .Q(n1827) );
  AO221X1 U853 ( .IN1(n1818), .IN2(n24), .IN3(n1594), .IN4(n7), .IN5(n1828), 
        .Q(n1677) );
  AO222X1 U854 ( .IN1(n1824), .IN2(n9), .IN3(n1596), .IN4(n29), .IN5(n1813), 
        .IN6(n114), .Q(n1828) );
  AO21X1 U855 ( .IN1(n1401), .IN2(n638), .IN3(n1788), .Q(
        \fpu_add_frac_dp/n3876 ) );
  AO22X1 U856 ( .IN1(n1809), .IN2(n1680), .IN3(n1816), .IN4(n1682), .Q(n1788)
         );
  AO221X1 U857 ( .IN1(n1669), .IN2(n615), .IN3(n1820), .IN4(n208), .IN5(n1829), 
        .Q(n1682) );
  AO22X1 U858 ( .IN1(n1667), .IN2(n176), .IN3(n1822), .IN4(n614), .Q(n1829) );
  AO221X1 U859 ( .IN1(n1818), .IN2(n25), .IN3(n1594), .IN4(n8), .IN5(n1830), 
        .Q(n1680) );
  AO222X1 U860 ( .IN1(n1824), .IN2(n24), .IN3(n1596), .IN4(n163), .IN5(n1813), 
        .IN6(n7), .Q(n1830) );
  AO21X1 U861 ( .IN1(n1401), .IN2(n281), .IN3(n1789), .Q(
        \fpu_add_frac_dp/n3875 ) );
  AO22X1 U862 ( .IN1(n1809), .IN2(n1683), .IN3(n1816), .IN4(n1685), .Q(n1789)
         );
  AO221X1 U863 ( .IN1(n1669), .IN2(n209), .IN3(n1820), .IN4(n99), .IN5(n1831), 
        .Q(n1685) );
  AO22X1 U864 ( .IN1(n1667), .IN2(n208), .IN3(n1822), .IN4(n615), .Q(n1831) );
  AO221X1 U865 ( .IN1(n1818), .IN2(n26), .IN3(n1594), .IN4(n9), .IN5(n1832), 
        .Q(n1683) );
  AO222X1 U866 ( .IN1(n1824), .IN2(n25), .IN3(n1596), .IN4(n164), .IN5(n1813), 
        .IN6(n8), .Q(n1832) );
  AO21X1 U867 ( .IN1(n1401), .IN2(n280), .IN3(n1790), .Q(
        \fpu_add_frac_dp/n3874 ) );
  AO22X1 U868 ( .IN1(n1809), .IN2(n1686), .IN3(n1816), .IN4(n1688), .Q(n1790)
         );
  AO221X1 U869 ( .IN1(n1669), .IN2(n210), .IN3(n1820), .IN4(n614), .IN5(n1833), 
        .Q(n1688) );
  AO22X1 U870 ( .IN1(n1667), .IN2(n99), .IN3(n1822), .IN4(n209), .Q(n1833) );
  AO221X1 U871 ( .IN1(n1818), .IN2(n76), .IN3(n1594), .IN4(n24), .IN5(n1834), 
        .Q(n1686) );
  AO222X1 U872 ( .IN1(n1824), .IN2(n26), .IN3(n1596), .IN4(n587), .IN5(n1813), 
        .IN6(n9), .Q(n1834) );
  AO21X1 U873 ( .IN1(n1401), .IN2(n217), .IN3(n1791), .Q(
        \fpu_add_frac_dp/n3873 ) );
  AO22X1 U874 ( .IN1(n1809), .IN2(n1689), .IN3(n1816), .IN4(n1691), .Q(n1791)
         );
  AO221X1 U875 ( .IN1(n1669), .IN2(n211), .IN3(n1820), .IN4(n615), .IN5(n1835), 
        .Q(n1691) );
  AO22X1 U876 ( .IN1(n1667), .IN2(n614), .IN3(n1822), .IN4(n210), .Q(n1835) );
  AO221X1 U877 ( .IN1(n1818), .IN2(n77), .IN3(n1594), .IN4(n25), .IN5(n1836), 
        .Q(n1689) );
  AO222X1 U878 ( .IN1(n1824), .IN2(n76), .IN3(n1596), .IN4(n588), .IN5(n1813), 
        .IN6(n24), .Q(n1836) );
  AO21X1 U879 ( .IN1(n1401), .IN2(n96), .IN3(n1792), .Q(
        \fpu_add_frac_dp/n3872 ) );
  AO22X1 U880 ( .IN1(n1809), .IN2(n1692), .IN3(n1816), .IN4(n1694), .Q(n1792)
         );
  AO221X1 U881 ( .IN1(n1669), .IN2(n616), .IN3(n1820), .IN4(n209), .IN5(n1837), 
        .Q(n1694) );
  AO22X1 U882 ( .IN1(n1667), .IN2(n615), .IN3(n1822), .IN4(n211), .Q(n1837) );
  AO221X1 U883 ( .IN1(n1818), .IN2(n167), .IN3(n1594), .IN4(n26), .IN5(n1838), 
        .Q(n1692) );
  AO222X1 U884 ( .IN1(n1824), .IN2(n77), .IN3(n1596), .IN4(n589), .IN5(n1813), 
        .IN6(n25), .Q(n1838) );
  AO21X1 U885 ( .IN1(n1400), .IN2(n631), .IN3(n1793), .Q(
        \fpu_add_frac_dp/n3871 ) );
  AO22X1 U886 ( .IN1(n1809), .IN2(n1695), .IN3(n1816), .IN4(n1697), .Q(n1793)
         );
  AO221X1 U887 ( .IN1(n1669), .IN2(n617), .IN3(n1820), .IN4(n210), .IN5(n1839), 
        .Q(n1697) );
  AO22X1 U888 ( .IN1(n1667), .IN2(n209), .IN3(n1822), .IN4(n616), .Q(n1839) );
  AO221X1 U889 ( .IN1(n1818), .IN2(n27), .IN3(n1594), .IN4(n76), .IN5(n1840), 
        .Q(n1695) );
  AO222X1 U890 ( .IN1(n1824), .IN2(n167), .IN3(n1596), .IN4(n78), .IN5(n1813), 
        .IN6(n26), .Q(n1840) );
  AO21X1 U891 ( .IN1(n1400), .IN2(n630), .IN3(n1794), .Q(
        \fpu_add_frac_dp/n3870 ) );
  AO22X1 U892 ( .IN1(n1809), .IN2(n1698), .IN3(n1816), .IN4(n1700), .Q(n1794)
         );
  AO221X1 U893 ( .IN1(n1669), .IN2(n618), .IN3(n1820), .IN4(n211), .IN5(n1841), 
        .Q(n1700) );
  AO22X1 U894 ( .IN1(n1667), .IN2(n210), .IN3(n1822), .IN4(n617), .Q(n1841) );
  AO221X1 U895 ( .IN1(n1818), .IN2(n28), .IN3(n1594), .IN4(n77), .IN5(n1842), 
        .Q(n1698) );
  AO222X1 U896 ( .IN1(n1824), .IN2(n27), .IN3(n1596), .IN4(n165), .IN5(n1813), 
        .IN6(n76), .Q(n1842) );
  AO21X1 U897 ( .IN1(n1400), .IN2(n632), .IN3(n1795), .Q(
        \fpu_add_frac_dp/n3869 ) );
  AO22X1 U898 ( .IN1(n1809), .IN2(n1701), .IN3(n1816), .IN4(n1703), .Q(n1795)
         );
  AO221X1 U899 ( .IN1(n1669), .IN2(n212), .IN3(n1820), .IN4(n616), .IN5(n1843), 
        .Q(n1703) );
  AO22X1 U900 ( .IN1(n1667), .IN2(n211), .IN3(n1822), .IN4(n618), .Q(n1843) );
  AO221X1 U901 ( .IN1(n1818), .IN2(n29), .IN3(n1594), .IN4(n167), .IN5(n1844), 
        .Q(n1701) );
  AO222X1 U902 ( .IN1(n1824), .IN2(n28), .IN3(n1596), .IN4(n169), .IN5(n1813), 
        .IN6(n77), .Q(n1844) );
  AO21X1 U903 ( .IN1(n1400), .IN2(n95), .IN3(n1796), .Q(
        \fpu_add_frac_dp/n3868 ) );
  AO22X1 U904 ( .IN1(n1809), .IN2(n1704), .IN3(n1816), .IN4(n1706), .Q(n1796)
         );
  AO221X1 U905 ( .IN1(n1669), .IN2(n213), .IN3(n1820), .IN4(n617), .IN5(n1845), 
        .Q(n1706) );
  AO22X1 U906 ( .IN1(n1667), .IN2(n616), .IN3(n1822), .IN4(n212), .Q(n1845) );
  AO221X1 U907 ( .IN1(n1818), .IN2(n163), .IN3(n1594), .IN4(n27), .IN5(n1846), 
        .Q(n1704) );
  AO222X1 U908 ( .IN1(n1824), .IN2(n29), .IN3(n1596), .IN4(n591), .IN5(n1813), 
        .IN6(n167), .Q(n1846) );
  AO21X1 U909 ( .IN1(n1400), .IN2(n613), .IN3(n1797), .Q(
        \fpu_add_frac_dp/n3867 ) );
  AO22X1 U910 ( .IN1(n1809), .IN2(n1707), .IN3(n1816), .IN4(n1709), .Q(n1797)
         );
  AO221X1 U911 ( .IN1(n1669), .IN2(n214), .IN3(n1820), .IN4(n618), .IN5(n1847), 
        .Q(n1709) );
  AO22X1 U912 ( .IN1(n1667), .IN2(n617), .IN3(n1822), .IN4(n213), .Q(n1847) );
  AO221X1 U913 ( .IN1(n1818), .IN2(n164), .IN3(n1594), .IN4(n28), .IN5(n1848), 
        .Q(n1707) );
  AO222X1 U914 ( .IN1(n1824), .IN2(n163), .IN3(n1596), .IN4(n592), .IN5(n1813), 
        .IN6(n27), .Q(n1848) );
  AO21X1 U915 ( .IN1(n1404), .IN2(n97), .IN3(n1798), .Q(
        \fpu_add_frac_dp/n3866 ) );
  AO22X1 U916 ( .IN1(n1809), .IN2(n1710), .IN3(n1816), .IN4(n1712), .Q(n1798)
         );
  AO221X1 U917 ( .IN1(n1669), .IN2(n619), .IN3(n1820), .IN4(n212), .IN5(n1849), 
        .Q(n1712) );
  AO22X1 U918 ( .IN1(n1667), .IN2(n618), .IN3(n1822), .IN4(n214), .Q(n1849) );
  AO221X1 U919 ( .IN1(n1818), .IN2(n587), .IN3(n1594), .IN4(n29), .IN5(n1850), 
        .Q(n1710) );
  AO222X1 U920 ( .IN1(n1824), .IN2(n164), .IN3(n1596), .IN4(n593), .IN5(n1813), 
        .IN6(n28), .Q(n1850) );
  AO21X1 U921 ( .IN1(n1400), .IN2(n98), .IN3(n1799), .Q(
        \fpu_add_frac_dp/n3865 ) );
  AO22X1 U922 ( .IN1(n1809), .IN2(n1713), .IN3(n1816), .IN4(n1715), .Q(n1799)
         );
  AO221X1 U923 ( .IN1(n1669), .IN2(n620), .IN3(n1820), .IN4(n213), .IN5(n1851), 
        .Q(n1715) );
  AO22X1 U924 ( .IN1(n1667), .IN2(n212), .IN3(n1822), .IN4(n619), .Q(n1851) );
  AO221X1 U925 ( .IN1(n1818), .IN2(n588), .IN3(n1594), .IN4(n163), .IN5(n1852), 
        .Q(n1713) );
  AO222X1 U926 ( .IN1(n1824), .IN2(n587), .IN3(n1596), .IN4(
        \fpu_add_frac_dp/n2446 ), .IN5(n1813), .IN6(n29), .Q(n1852) );
  AO21X1 U927 ( .IN1(n1400), .IN2(n4), .IN3(n1800), .Q(\fpu_add_frac_dp/n3864 ) );
  AO22X1 U928 ( .IN1(n1809), .IN2(n1716), .IN3(n1816), .IN4(n1718), .Q(n1800)
         );
  AO221X1 U929 ( .IN1(n1669), .IN2(n621), .IN3(n1820), .IN4(n214), .IN5(n1853), 
        .Q(n1718) );
  AO22X1 U930 ( .IN1(n1667), .IN2(n213), .IN3(n1822), .IN4(n620), .Q(n1853) );
  AO221X1 U931 ( .IN1(n1818), .IN2(n589), .IN3(n1594), .IN4(n164), .IN5(n1854), 
        .Q(n1716) );
  AO222X1 U932 ( .IN1(n1824), .IN2(n588), .IN3(n1596), .IN4(
        \fpu_add_frac_dp/n2473 ), .IN5(n1813), .IN6(n163), .Q(n1854) );
  AO21X1 U933 ( .IN1(n1397), .IN2(n157), .IN3(n1801), .Q(
        \fpu_add_frac_dp/n3863 ) );
  AO22X1 U934 ( .IN1(n1809), .IN2(n1719), .IN3(n1816), .IN4(n1721), .Q(n1801)
         );
  AO221X1 U935 ( .IN1(n1669), .IN2(n215), .IN3(n1820), .IN4(n619), .IN5(n1855), 
        .Q(n1721) );
  AO22X1 U936 ( .IN1(n1667), .IN2(n214), .IN3(n1822), .IN4(n621), .Q(n1855) );
  AO221X1 U937 ( .IN1(n1818), .IN2(n78), .IN3(n1594), .IN4(n587), .IN5(n1856), 
        .Q(n1719) );
  AO222X1 U938 ( .IN1(n1824), .IN2(n589), .IN3(n1596), .IN4(
        \fpu_add_frac_dp/n2466 ), .IN5(n1813), .IN6(n164), .Q(n1856) );
  AO21X1 U939 ( .IN1(n1397), .IN2(n1857), .IN3(n1802), .Q(
        \fpu_add_frac_dp/n3862 ) );
  AO22X1 U940 ( .IN1(n1809), .IN2(n1722), .IN3(n1816), .IN4(n1724), .Q(n1802)
         );
  AO221X1 U941 ( .IN1(n1669), .IN2(n216), .IN3(n1820), .IN4(n620), .IN5(n1858), 
        .Q(n1724) );
  AO22X1 U942 ( .IN1(n1667), .IN2(n619), .IN3(n1822), .IN4(n215), .Q(n1858) );
  AO221X1 U943 ( .IN1(n1818), .IN2(n165), .IN3(n1594), .IN4(n588), .IN5(n1859), 
        .Q(n1722) );
  AO222X1 U944 ( .IN1(n1824), .IN2(n78), .IN3(n1596), .IN4(
        \fpu_add_frac_dp/n2474 ), .IN5(n1813), .IN6(n587), .Q(n1859) );
  AO21X1 U945 ( .IN1(n1397), .IN2(n68), .IN3(n1803), .Q(
        \fpu_add_frac_dp/n3861 ) );
  AO22X1 U946 ( .IN1(n1809), .IN2(n1725), .IN3(n1816), .IN4(n1727), .Q(n1803)
         );
  AO221X1 U947 ( .IN1(n1669), .IN2(n206), .IN3(n1820), .IN4(n621), .IN5(n1860), 
        .Q(n1727) );
  AO22X1 U948 ( .IN1(n1667), .IN2(n620), .IN3(n1822), .IN4(n216), .Q(n1860) );
  AO221X1 U949 ( .IN1(n1818), .IN2(n169), .IN3(n1594), .IN4(n589), .IN5(n1861), 
        .Q(n1725) );
  AO222X1 U950 ( .IN1(n1824), .IN2(n165), .IN3(n1596), .IN4(
        \fpu_add_frac_dp/n2467 ), .IN5(n1813), .IN6(n588), .Q(n1861) );
  AO21X1 U951 ( .IN1(n1397), .IN2(n156), .IN3(n1804), .Q(
        \fpu_add_frac_dp/n3860 ) );
  AO22X1 U952 ( .IN1(n1809), .IN2(n1728), .IN3(n1816), .IN4(n1730), .Q(n1804)
         );
  AO221X1 U953 ( .IN1(n1669), .IN2(n688), .IN3(n1820), .IN4(n215), .IN5(n1862), 
        .Q(n1730) );
  AO22X1 U954 ( .IN1(n1667), .IN2(n621), .IN3(n1822), .IN4(n206), .Q(n1862) );
  AO221X1 U955 ( .IN1(n1818), .IN2(n591), .IN3(n1594), .IN4(n78), .IN5(n1863), 
        .Q(n1728) );
  AO222X1 U956 ( .IN1(n1824), .IN2(n169), .IN3(n1596), .IN4(
        \fpu_add_frac_dp/n2475 ), .IN5(n1813), .IN6(n589), .Q(n1863) );
  AO21X1 U957 ( .IN1(n1397), .IN2(n3), .IN3(n1805), .Q(\fpu_add_frac_dp/n3859 ) );
  AO22X1 U958 ( .IN1(n1809), .IN2(n1731), .IN3(n1816), .IN4(n1733), .Q(n1805)
         );
  AO221X1 U959 ( .IN1(n1669), .IN2(n689), .IN3(n1820), .IN4(n216), .IN5(n1864), 
        .Q(n1733) );
  AO22X1 U960 ( .IN1(n1667), .IN2(n215), .IN3(n1822), .IN4(n688), .Q(n1864) );
  AO221X1 U961 ( .IN1(n1818), .IN2(n592), .IN3(n1594), .IN4(n165), .IN5(n1865), 
        .Q(n1731) );
  AO222X1 U962 ( .IN1(n1824), .IN2(n591), .IN3(n1596), .IN4(
        \fpu_add_frac_dp/n2468 ), .IN5(n1813), .IN6(n78), .Q(n1865) );
  AO21X1 U963 ( .IN1(n1397), .IN2(n16), .IN3(n1806), .Q(
        \fpu_add_frac_dp/n3858 ) );
  AO22X1 U964 ( .IN1(n1816), .IN2(n1738), .IN3(n1809), .IN4(n1866), .Q(n1806)
         );
  AO21X1 U965 ( .IN1(n1751), .IN2(n1867), .IN3(n1734), .Q(n1866) );
  AO221X1 U966 ( .IN1(n1818), .IN2(n593), .IN3(n1594), .IN4(n169), .IN5(n1868), 
        .Q(n1734) );
  AO222X1 U967 ( .IN1(n1824), .IN2(n592), .IN3(n1596), .IN4(
        \fpu_add_frac_dp/n2469 ), .IN5(n1813), .IN6(n165), .Q(n1868) );
  INVX0 U968 ( .INP(n1869), .ZN(n1818) );
  AO221X1 U969 ( .IN1(n1669), .IN2(n705), .IN3(n1820), .IN4(n206), .IN5(n1870), 
        .Q(n1738) );
  AO22X1 U970 ( .IN1(n1667), .IN2(n216), .IN3(n1822), .IN4(n689), .Q(n1870) );
  INVX0 U971 ( .INP(n1665), .ZN(n1820) );
  INVX0 U972 ( .INP(n1817), .ZN(n1669) );
  AO21X1 U973 ( .IN1(n1397), .IN2(n15), .IN3(n1807), .Q(
        \fpu_add_frac_dp/n3857 ) );
  AO22X1 U974 ( .IN1(n1816), .IN2(n1743), .IN3(n1809), .IN4(n1742), .Q(n1807)
         );
  NAND4X0 U975 ( .IN1(n1869), .IN2(n1811), .IN3(n1871), .IN4(n1872), .QN(n1742) );
  AOI22X1 U976 ( .IN1(n593), .IN2(n1824), .IN3(n169), .IN4(n1813), .QN(n1872)
         );
  NOR2X0 U977 ( .IN1(\fpu_add_ctl/n117 ), .IN2(\fpu_add_ctl/n327 ), .QN(n1813)
         );
  NOR2X0 U978 ( .IN1(\fpu_add_ctl/n117 ), .IN2(\fpu_add_ctl/n328 ), .QN(n1824)
         );
  NAND2X0 U979 ( .IN1(n1596), .IN2(n1080), .QN(n1871) );
  NAND2X0 U980 ( .IN1(\fpu_add_ctl/n117 ), .IN2(n700), .QN(n1811) );
  NAND2X0 U981 ( .IN1(\fpu_add_ctl/n117 ), .IN2(n701), .QN(n1869) );
  AOI21X1 U982 ( .IN1(n1737), .IN2(n1873), .IN3(n1745), .QN(n1809) );
  NAND2X0 U983 ( .IN1(n1874), .IN2(n1875), .QN(n1873) );
  INVX0 U984 ( .INP(n1748), .ZN(n1875) );
  NAND3X0 U985 ( .IN1(n1817), .IN2(n1665), .IN3(n1876), .QN(n1743) );
  AOI22X1 U986 ( .IN1(n705), .IN2(n1822), .IN3(n206), .IN4(n1667), .QN(n1876)
         );
  NOR2X0 U987 ( .IN1(\fpu_add_ctl/n122 ), .IN2(\fpu_add_ctl/n327 ), .QN(n1667)
         );
  NOR2X0 U988 ( .IN1(\fpu_add_ctl/n122 ), .IN2(\fpu_add_ctl/n328 ), .QN(n1822)
         );
  NAND2X0 U989 ( .IN1(\fpu_add_ctl/n122 ), .IN2(n700), .QN(n1665) );
  NAND2X0 U990 ( .IN1(\fpu_add_ctl/n122 ), .IN2(n701), .QN(n1817) );
  AND3X1 U991 ( .IN1(n1449), .IN2(n1748), .IN3(n1874), .Q(n1816) );
  NOR2X0 U992 ( .IN1(n1867), .IN2(n1877), .QN(n1874) );
  AO222X1 U993 ( .IN1(\fpu_add_exp_dp/n45 ), .IN2(n1878), .IN3(
        \fpu_add_exp_dp/n47 ), .IN4(n1879), .IN5(n1880), .IN6(n1881), .Q(n1748) );
  NAND2X0 U994 ( .IN1(n961), .IN2(n1882), .QN(n1879) );
  INVX0 U995 ( .INP(n1882), .ZN(n1878) );
  AO22X1 U996 ( .IN1(n1883), .IN2(n445), .IN3(n1884), .IN4(n1000), .Q(n1882)
         );
  OR2X1 U997 ( .IN1(n445), .IN2(n1883), .Q(n1884) );
  AO22X1 U998 ( .IN1(n1885), .IN2(n446), .IN3(n1886), .IN4(n999), .Q(n1883) );
  OR2X1 U999 ( .IN1(n446), .IN2(n1885), .Q(n1886) );
  AO22X1 U1000 ( .IN1(n1887), .IN2(n323), .IN3(n1888), .IN4(n998), .Q(n1885)
         );
  OR2X1 U1001 ( .IN1(n323), .IN2(n1887), .Q(n1888) );
  AO22X1 U1002 ( .IN1(n1889), .IN2(n322), .IN3(n1890), .IN4(n997), .Q(n1887)
         );
  OR2X1 U1003 ( .IN1(n322), .IN2(n1889), .Q(n1890) );
  AO22X1 U1004 ( .IN1(n1891), .IN2(n321), .IN3(n1892), .IN4(n996), .Q(n1889)
         );
  OR2X1 U1005 ( .IN1(n321), .IN2(n1891), .Q(n1892) );
  AO22X1 U1006 ( .IN1(n1893), .IN2(n320), .IN3(n1894), .IN4(n995), .Q(n1891)
         );
  OR2X1 U1007 ( .IN1(n320), .IN2(n1893), .Q(n1894) );
  AO22X1 U1008 ( .IN1(n1895), .IN2(n319), .IN3(n1896), .IN4(n994), .Q(n1893)
         );
  OR2X1 U1009 ( .IN1(n319), .IN2(n1895), .Q(n1896) );
  AO22X1 U1010 ( .IN1(n1897), .IN2(n309), .IN3(n1898), .IN4(n993), .Q(n1895)
         );
  OR2X1 U1011 ( .IN1(n309), .IN2(n1897), .Q(n1898) );
  AO21X1 U1012 ( .IN1(n56), .IN2(n138), .IN3(n1899), .Q(n1897) );
  OA22X1 U1013 ( .IN1(n56), .IN2(n138), .IN3(n491), .IN4(n992), .Q(n1899) );
  AO22X1 U1014 ( .IN1(n1443), .IN2(n625), .IN3(n1409), .IN4(n465), .Q(
        \fpu_add_frac_dp/n3856 ) );
  AO22X1 U1015 ( .IN1(n1443), .IN2(n220), .IN3(n1409), .IN4(n828), .Q(
        \fpu_add_frac_dp/n3855 ) );
  AO22X1 U1016 ( .IN1(n1443), .IN2(n310), .IN3(n1410), .IN4(n827), .Q(
        \fpu_add_frac_dp/n3854 ) );
  AO22X1 U1017 ( .IN1(n1443), .IN2(n288), .IN3(n1409), .IN4(n826), .Q(
        \fpu_add_frac_dp/n3853 ) );
  AO22X1 U1018 ( .IN1(n1443), .IN2(n223), .IN3(n1409), .IN4(n825), .Q(
        \fpu_add_frac_dp/n3852 ) );
  AO22X1 U1019 ( .IN1(n1443), .IN2(n225), .IN3(n1409), .IN4(n824), .Q(
        \fpu_add_frac_dp/n3851 ) );
  AO22X1 U1020 ( .IN1(n1443), .IN2(n222), .IN3(n1409), .IN4(n823), .Q(
        \fpu_add_frac_dp/n3850 ) );
  AO22X1 U1021 ( .IN1(n1443), .IN2(n224), .IN3(n1409), .IN4(n822), .Q(
        \fpu_add_frac_dp/n3849 ) );
  AO22X1 U1022 ( .IN1(n1443), .IN2(n261), .IN3(n1409), .IN4(n821), .Q(
        \fpu_add_frac_dp/n3848 ) );
  AO22X1 U1023 ( .IN1(n1443), .IN2(n260), .IN3(n1409), .IN4(n820), .Q(
        \fpu_add_frac_dp/n3847 ) );
  AO22X1 U1024 ( .IN1(n1443), .IN2(n253), .IN3(n1409), .IN4(n819), .Q(
        \fpu_add_frac_dp/n3846 ) );
  AO22X1 U1025 ( .IN1(n1443), .IN2(n252), .IN3(n1409), .IN4(n818), .Q(
        \fpu_add_frac_dp/n3845 ) );
  AO22X1 U1026 ( .IN1(n1443), .IN2(n327), .IN3(n1408), .IN4(n817), .Q(
        \fpu_add_frac_dp/n3844 ) );
  AO22X1 U1027 ( .IN1(n1443), .IN2(n180), .IN3(n1408), .IN4(n816), .Q(
        \fpu_add_frac_dp/n3843 ) );
  AO22X1 U1028 ( .IN1(n1443), .IN2(n268), .IN3(n1409), .IN4(n815), .Q(
        \fpu_add_frac_dp/n3842 ) );
  AO22X1 U1029 ( .IN1(n1444), .IN2(n179), .IN3(n1408), .IN4(n814), .Q(
        \fpu_add_frac_dp/n3841 ) );
  AO22X1 U1030 ( .IN1(n1443), .IN2(n251), .IN3(n1408), .IN4(n813), .Q(
        \fpu_add_frac_dp/n3840 ) );
  AO22X1 U1031 ( .IN1(n1444), .IN2(n250), .IN3(n1409), .IN4(n812), .Q(
        \fpu_add_frac_dp/n3839 ) );
  AO22X1 U1032 ( .IN1(n1444), .IN2(n249), .IN3(n1409), .IN4(n811), .Q(
        \fpu_add_frac_dp/n3838 ) );
  AO22X1 U1033 ( .IN1(n1444), .IN2(n263), .IN3(n1408), .IN4(n810), .Q(
        \fpu_add_frac_dp/n3837 ) );
  AO22X1 U1034 ( .IN1(n1444), .IN2(n267), .IN3(n1408), .IN4(n809), .Q(
        \fpu_add_frac_dp/n3836 ) );
  AO22X1 U1035 ( .IN1(n1444), .IN2(n279), .IN3(n1408), .IN4(n808), .Q(
        \fpu_add_frac_dp/n3835 ) );
  AO22X1 U1036 ( .IN1(n1444), .IN2(n318), .IN3(n1408), .IN4(n807), .Q(
        \fpu_add_frac_dp/n3834 ) );
  AO22X1 U1037 ( .IN1(n1444), .IN2(n248), .IN3(n1408), .IN4(n806), .Q(
        \fpu_add_frac_dp/n3833 ) );
  AO22X1 U1038 ( .IN1(n1444), .IN2(n247), .IN3(n1408), .IN4(n805), .Q(
        \fpu_add_frac_dp/n3832 ) );
  AO22X1 U1039 ( .IN1(n1444), .IN2(n246), .IN3(n1408), .IN4(n804), .Q(
        \fpu_add_frac_dp/n3831 ) );
  AO22X1 U1040 ( .IN1(n1444), .IN2(n204), .IN3(n1410), .IN4(n803), .Q(
        \fpu_add_frac_dp/n3830 ) );
  AO22X1 U1041 ( .IN1(n1444), .IN2(n245), .IN3(n1407), .IN4(n802), .Q(
        \fpu_add_frac_dp/n3829 ) );
  AO22X1 U1042 ( .IN1(n1444), .IN2(n244), .IN3(n1407), .IN4(n801), .Q(
        \fpu_add_frac_dp/n3828 ) );
  AO22X1 U1043 ( .IN1(n1446), .IN2(n203), .IN3(n1408), .IN4(n800), .Q(
        \fpu_add_frac_dp/n3827 ) );
  AO22X1 U1044 ( .IN1(n1444), .IN2(n243), .IN3(n1407), .IN4(n799), .Q(
        \fpu_add_frac_dp/n3826 ) );
  AO22X1 U1045 ( .IN1(n1444), .IN2(n242), .IN3(n1407), .IN4(n798), .Q(
        \fpu_add_frac_dp/n3825 ) );
  AO22X1 U1046 ( .IN1(n1444), .IN2(n241), .IN3(n1407), .IN4(n797), .Q(
        \fpu_add_frac_dp/n3824 ) );
  AO22X1 U1047 ( .IN1(n1444), .IN2(n240), .IN3(n1407), .IN4(n796), .Q(
        \fpu_add_frac_dp/n3823 ) );
  AO22X1 U1048 ( .IN1(n1446), .IN2(n202), .IN3(n1407), .IN4(n795), .Q(
        \fpu_add_frac_dp/n3822 ) );
  AO22X1 U1049 ( .IN1(n1444), .IN2(n239), .IN3(n1408), .IN4(n794), .Q(
        \fpu_add_frac_dp/n3821 ) );
  AO22X1 U1050 ( .IN1(n1445), .IN2(n201), .IN3(n1407), .IN4(n793), .Q(
        \fpu_add_frac_dp/n3820 ) );
  AO22X1 U1051 ( .IN1(n1445), .IN2(n238), .IN3(n1407), .IN4(n792), .Q(
        \fpu_add_frac_dp/n3819 ) );
  AO22X1 U1052 ( .IN1(n1445), .IN2(n200), .IN3(n1407), .IN4(n791), .Q(
        \fpu_add_frac_dp/n3818 ) );
  AO22X1 U1053 ( .IN1(n1445), .IN2(n259), .IN3(n1408), .IN4(n790), .Q(
        \fpu_add_frac_dp/n3817 ) );
  AO22X1 U1054 ( .IN1(n1445), .IN2(n237), .IN3(n1406), .IN4(n789), .Q(
        \fpu_add_frac_dp/n3816 ) );
  AO22X1 U1055 ( .IN1(n1445), .IN2(n199), .IN3(n1407), .IN4(n788), .Q(
        \fpu_add_frac_dp/n3815 ) );
  AO22X1 U1056 ( .IN1(n1445), .IN2(n236), .IN3(n1406), .IN4(n787), .Q(
        \fpu_add_frac_dp/n3814 ) );
  AO22X1 U1057 ( .IN1(n1445), .IN2(n235), .IN3(n1406), .IN4(n786), .Q(
        \fpu_add_frac_dp/n3813 ) );
  AO22X1 U1058 ( .IN1(n1445), .IN2(n234), .IN3(n1407), .IN4(n785), .Q(
        \fpu_add_frac_dp/n3812 ) );
  AO22X1 U1059 ( .IN1(n1445), .IN2(n198), .IN3(n1406), .IN4(n784), .Q(
        \fpu_add_frac_dp/n3811 ) );
  AO22X1 U1060 ( .IN1(n1445), .IN2(n197), .IN3(n1406), .IN4(n783), .Q(
        \fpu_add_frac_dp/n3810 ) );
  AO22X1 U1061 ( .IN1(n1445), .IN2(n233), .IN3(n1407), .IN4(n782), .Q(
        \fpu_add_frac_dp/n3809 ) );
  AO22X1 U1062 ( .IN1(n1445), .IN2(n232), .IN3(n1406), .IN4(n781), .Q(
        \fpu_add_frac_dp/n3808 ) );
  AO22X1 U1063 ( .IN1(n1445), .IN2(n231), .IN3(n1406), .IN4(n780), .Q(
        \fpu_add_frac_dp/n3807 ) );
  AO22X1 U1064 ( .IN1(n1445), .IN2(n230), .IN3(n1407), .IN4(n779), .Q(
        \fpu_add_frac_dp/n3806 ) );
  AO22X1 U1065 ( .IN1(n1445), .IN2(n229), .IN3(n1406), .IN4(n778), .Q(
        \fpu_add_frac_dp/n3805 ) );
  AO22X1 U1066 ( .IN1(n1445), .IN2(n228), .IN3(n1406), .IN4(n777), .Q(
        \fpu_add_frac_dp/n3804 ) );
  AO22X1 U1067 ( .IN1(n1445), .IN2(n227), .IN3(n1406), .IN4(n776), .Q(
        \fpu_add_frac_dp/n3803 ) );
  AO22X1 U1068 ( .IN1(n1446), .IN2(n196), .IN3(n1414), .IN4(n775), .Q(
        \fpu_add_frac_dp/n3802 ) );
  AO22X1 U1069 ( .IN1(n1446), .IN2(n294), .IN3(n1406), .IN4(n774), .Q(
        \fpu_add_frac_dp/n3801 ) );
  AO22X1 U1070 ( .IN1(n1446), .IN2(n332), .IN3(n1410), .IN4(n773), .Q(
        \fpu_add_frac_dp/n3800 ) );
  AO22X1 U1071 ( .IN1(n1446), .IN2(n334), .IN3(n1414), .IN4(n772), .Q(
        \fpu_add_frac_dp/n3799 ) );
  AO22X1 U1072 ( .IN1(n1446), .IN2(n293), .IN3(n1414), .IN4(n771), .Q(
        \fpu_add_frac_dp/n3798 ) );
  AO22X1 U1073 ( .IN1(n1446), .IN2(n317), .IN3(n1414), .IN4(n770), .Q(
        \fpu_add_frac_dp/n3797 ) );
  AO22X1 U1074 ( .IN1(n1446), .IN2(n195), .IN3(n1415), .IN4(n769), .Q(
        \fpu_add_frac_dp/n3796 ) );
  AO22X1 U1075 ( .IN1(n1446), .IN2(n226), .IN3(n1415), .IN4(n768), .Q(
        \fpu_add_frac_dp/n3795 ) );
  AO22X1 U1076 ( .IN1(n1446), .IN2(n850), .IN3(n1415), .IN4(n453), .Q(
        \fpu_add_frac_dp/n3794 ) );
  AO22X1 U1077 ( .IN1(n1416), .IN2(n1274), .IN3(n1900), .IN4(n1901), .Q(
        \fpu_add_frac_dp/n3792 ) );
  AO22X1 U1078 ( .IN1(n1426), .IN2(n1081), .IN3(n1902), .IN4(n1900), .Q(
        \fpu_add_frac_dp/n3791 ) );
  AO22X1 U1079 ( .IN1(n1422), .IN2(n1250), .IN3(n1903), .IN4(n1904), .Q(
        \fpu_add_frac_dp/n3790 ) );
  AO22X1 U1080 ( .IN1(n1422), .IN2(n1275), .IN3(n1903), .IN4(n1905), .Q(
        \fpu_add_frac_dp/n3789 ) );
  NOR2X0 U1081 ( .IN1(\fpu_add_exp_dp/n146 ), .IN2(n1906), .QN(n1903) );
  AO22X1 U1082 ( .IN1(n1423), .IN2(n1276), .IN3(n1904), .IN4(n1900), .Q(
        \fpu_add_frac_dp/n3788 ) );
  AO22X1 U1083 ( .IN1(n1423), .IN2(n1273), .IN3(n1905), .IN4(n1900), .Q(
        \fpu_add_frac_dp/n3787 ) );
  NOR2X0 U1084 ( .IN1(n73), .IN2(n1906), .QN(n1900) );
  NAND2X0 U1085 ( .IN1(n1907), .IN2(n1908), .QN(n1906) );
  AO22X1 U1086 ( .IN1(n1423), .IN2(n1251), .IN3(n1909), .IN4(n1910), .Q(
        \fpu_add_frac_dp/n3786 ) );
  AO22X1 U1087 ( .IN1(n1423), .IN2(n1277), .IN3(n1911), .IN4(n1910), .Q(
        \fpu_add_frac_dp/n3785 ) );
  AO22X1 U1088 ( .IN1(n1423), .IN2(n1266), .IN3(n1912), .IN4(n1910), .Q(
        \fpu_add_frac_dp/n3784 ) );
  AO22X1 U1089 ( .IN1(n1423), .IN2(n1247), .IN3(n1913), .IN4(n1910), .Q(
        \fpu_add_frac_dp/n3783 ) );
  AO22X1 U1090 ( .IN1(n1423), .IN2(n1278), .IN3(n1914), .IN4(n1910), .Q(
        \fpu_add_frac_dp/n3782 ) );
  AO22X1 U1091 ( .IN1(n1423), .IN2(n1279), .IN3(n1915), .IN4(n1910), .Q(
        \fpu_add_frac_dp/n3781 ) );
  AO22X1 U1092 ( .IN1(n1423), .IN2(n1280), .IN3(n1916), .IN4(n1910), .Q(
        \fpu_add_frac_dp/n3780 ) );
  AO22X1 U1093 ( .IN1(n1423), .IN2(n1281), .IN3(n1917), .IN4(n1910), .Q(
        \fpu_add_frac_dp/n3779 ) );
  AO22X1 U1094 ( .IN1(n1423), .IN2(n1252), .IN3(n1909), .IN4(n1908), .Q(
        \fpu_add_frac_dp/n3778 ) );
  AO22X1 U1095 ( .IN1(n1423), .IN2(n1282), .IN3(n1911), .IN4(n1908), .Q(
        \fpu_add_frac_dp/n3777 ) );
  AO22X1 U1096 ( .IN1(n1423), .IN2(n1283), .IN3(n1912), .IN4(n1908), .Q(
        \fpu_add_frac_dp/n3776 ) );
  AO22X1 U1097 ( .IN1(n1423), .IN2(n1267), .IN3(n1913), .IN4(n1908), .Q(
        \fpu_add_frac_dp/n3775 ) );
  AO22X1 U1098 ( .IN1(n1423), .IN2(n1253), .IN3(n1914), .IN4(n1908), .Q(
        \fpu_add_frac_dp/n3774 ) );
  AO22X1 U1099 ( .IN1(n1424), .IN2(n1284), .IN3(n1915), .IN4(n1908), .Q(
        \fpu_add_frac_dp/n3773 ) );
  AO22X1 U1100 ( .IN1(n1424), .IN2(n1268), .IN3(n1916), .IN4(n1908), .Q(
        \fpu_add_frac_dp/n3772 ) );
  AO22X1 U1101 ( .IN1(n1424), .IN2(n1269), .IN3(n1917), .IN4(n1908), .Q(
        \fpu_add_frac_dp/n3771 ) );
  NOR2X0 U1102 ( .IN1(n290), .IN2(\fpu_add_exp_dp/n142 ), .QN(n1908) );
  AO22X1 U1103 ( .IN1(n1424), .IN2(n1254), .IN3(n1918), .IN4(n1901), .Q(
        \fpu_add_frac_dp/n3770 ) );
  AO22X1 U1104 ( .IN1(n1424), .IN2(n1285), .IN3(n1918), .IN4(n1902), .Q(
        \fpu_add_frac_dp/n3769 ) );
  AO22X1 U1105 ( .IN1(n1424), .IN2(n1243), .IN3(n1919), .IN4(n1901), .Q(
        \fpu_add_frac_dp/n3768 ) );
  AO22X1 U1106 ( .IN1(n1424), .IN2(n1255), .IN3(n1919), .IN4(n1902), .Q(
        \fpu_add_frac_dp/n3767 ) );
  AO22X1 U1107 ( .IN1(n1424), .IN2(n1286), .IN3(n1918), .IN4(n1904), .Q(
        \fpu_add_frac_dp/n3766 ) );
  AO22X1 U1108 ( .IN1(n1424), .IN2(n1256), .IN3(n1918), .IN4(n1905), .Q(
        \fpu_add_frac_dp/n3765 ) );
  AND3X1 U1109 ( .IN1(n1907), .IN2(n73), .IN3(n1920), .Q(n1918) );
  AO22X1 U1110 ( .IN1(n1424), .IN2(n1287), .IN3(n1919), .IN4(n1904), .Q(
        \fpu_add_frac_dp/n3764 ) );
  AO22X1 U1111 ( .IN1(n1424), .IN2(n1288), .IN3(n1919), .IN4(n1905), .Q(
        \fpu_add_frac_dp/n3763 ) );
  AND3X1 U1112 ( .IN1(\fpu_add_exp_dp/n146 ), .IN2(n1907), .IN3(n1920), .Q(
        n1919) );
  AO22X1 U1113 ( .IN1(n1424), .IN2(n1257), .IN3(n1921), .IN4(n1901), .Q(
        \fpu_add_frac_dp/n3762 ) );
  AO22X1 U1114 ( .IN1(n1424), .IN2(n1289), .IN3(n1921), .IN4(n1902), .Q(
        \fpu_add_frac_dp/n3761 ) );
  AO22X1 U1115 ( .IN1(n1424), .IN2(n1290), .IN3(n1922), .IN4(n1901), .Q(
        \fpu_add_frac_dp/n3760 ) );
  AO22X1 U1116 ( .IN1(n1424), .IN2(n1291), .IN3(n1922), .IN4(n1902), .Q(
        \fpu_add_frac_dp/n3759 ) );
  AO22X1 U1117 ( .IN1(n1425), .IN2(n1258), .IN3(n1921), .IN4(n1904), .Q(
        \fpu_add_frac_dp/n3758 ) );
  AO22X1 U1118 ( .IN1(n1425), .IN2(n1292), .IN3(n1921), .IN4(n1905), .Q(
        \fpu_add_frac_dp/n3757 ) );
  AND2X1 U1119 ( .IN1(n1923), .IN2(n73), .Q(n1921) );
  AO22X1 U1120 ( .IN1(n1425), .IN2(n1259), .IN3(n1922), .IN4(n1904), .Q(
        \fpu_add_frac_dp/n3756 ) );
  AO22X1 U1121 ( .IN1(n1425), .IN2(n1293), .IN3(n1922), .IN4(n1905), .Q(
        \fpu_add_frac_dp/n3755 ) );
  AND2X1 U1122 ( .IN1(n1923), .IN2(\fpu_add_exp_dp/n146 ), .Q(n1922) );
  AND2X1 U1123 ( .IN1(n1924), .IN2(n1907), .Q(n1923) );
  AND2X1 U1124 ( .IN1(n1925), .IN2(n648), .Q(n1907) );
  AO22X1 U1125 ( .IN1(n1425), .IN2(n1260), .IN3(n1920), .IN4(n1909), .Q(
        \fpu_add_frac_dp/n3754 ) );
  AO22X1 U1126 ( .IN1(n1425), .IN2(n1294), .IN3(n1920), .IN4(n1911), .Q(
        \fpu_add_frac_dp/n3753 ) );
  AO22X1 U1127 ( .IN1(n1425), .IN2(n1295), .IN3(n1920), .IN4(n1912), .Q(
        \fpu_add_frac_dp/n3752 ) );
  AO22X1 U1128 ( .IN1(n1425), .IN2(n1224), .IN3(n1920), .IN4(n1913), .Q(
        \fpu_add_frac_dp/n3751 ) );
  AO22X1 U1129 ( .IN1(n1425), .IN2(n1261), .IN3(n1920), .IN4(n1914), .Q(
        \fpu_add_frac_dp/n3750 ) );
  AO22X1 U1130 ( .IN1(n1425), .IN2(n1296), .IN3(n1920), .IN4(n1915), .Q(
        \fpu_add_frac_dp/n3749 ) );
  AO22X1 U1131 ( .IN1(n1425), .IN2(n1297), .IN3(n1920), .IN4(n1916), .Q(
        \fpu_add_frac_dp/n3748 ) );
  AO22X1 U1132 ( .IN1(n1425), .IN2(n1244), .IN3(n1920), .IN4(n1917), .Q(
        \fpu_add_frac_dp/n3747 ) );
  AO22X1 U1133 ( .IN1(n1425), .IN2(n1262), .IN3(n1924), .IN4(n1909), .Q(
        \fpu_add_frac_dp/n3746 ) );
  AND2X1 U1134 ( .IN1(n1926), .IN2(n1901), .Q(n1909) );
  AO22X1 U1135 ( .IN1(n1425), .IN2(n1298), .IN3(n1924), .IN4(n1911), .Q(
        \fpu_add_frac_dp/n3745 ) );
  AND2X1 U1136 ( .IN1(n1926), .IN2(n1902), .Q(n1911) );
  AO22X1 U1137 ( .IN1(n1425), .IN2(n1299), .IN3(n1924), .IN4(n1912), .Q(
        \fpu_add_frac_dp/n3744 ) );
  AND2X1 U1138 ( .IN1(n1927), .IN2(n1901), .Q(n1912) );
  AO22X1 U1139 ( .IN1(n1426), .IN2(n1270), .IN3(n1924), .IN4(n1913), .Q(
        \fpu_add_frac_dp/n3743 ) );
  AND2X1 U1140 ( .IN1(n1927), .IN2(n1902), .Q(n1913) );
  NOR2X0 U1141 ( .IN1(n645), .IN2(\fpu_add_exp_dp/n145 ), .QN(n1902) );
  AO22X1 U1142 ( .IN1(n1426), .IN2(n1263), .IN3(n1924), .IN4(n1914), .Q(
        \fpu_add_frac_dp/n3742 ) );
  AND2X1 U1143 ( .IN1(n1926), .IN2(n1904), .Q(n1914) );
  AO22X1 U1144 ( .IN1(n1426), .IN2(n1300), .IN3(n1924), .IN4(n1915), .Q(
        \fpu_add_frac_dp/n3741 ) );
  AND2X1 U1145 ( .IN1(n1926), .IN2(n1905), .Q(n1915) );
  AND2X1 U1146 ( .IN1(n1928), .IN2(n73), .Q(n1926) );
  AO22X1 U1147 ( .IN1(n1426), .IN2(n1301), .IN3(n1924), .IN4(n1916), .Q(
        \fpu_add_frac_dp/n3740 ) );
  AND2X1 U1148 ( .IN1(n1927), .IN2(n1904), .Q(n1916) );
  NOR2X0 U1149 ( .IN1(n287), .IN2(\fpu_add_exp_dp/n147 ), .QN(n1904) );
  AO22X1 U1150 ( .IN1(n1426), .IN2(n1235), .IN3(n1924), .IN4(n1917), .Q(
        \fpu_add_frac_dp/n3739 ) );
  AND2X1 U1151 ( .IN1(n1927), .IN2(n1905), .Q(n1917) );
  NOR2X0 U1152 ( .IN1(n287), .IN2(n645), .QN(n1905) );
  AND2X1 U1153 ( .IN1(n1928), .IN2(\fpu_add_exp_dp/n146 ), .Q(n1927) );
  AND2X1 U1154 ( .IN1(\fpu_add_exp_dp/n143 ), .IN2(n1925), .Q(n1928) );
  AND4X1 U1155 ( .IN1(\fpu_add_exp_dp/n137 ), .IN2(n1929), .IN3(n1449), .IN4(
        n640), .Q(n1925) );
  AO21X1 U1156 ( .IN1(n1396), .IN2(n1219), .IN3(n1930), .Q(
        \fpu_add_frac_dp/n3738 ) );
  AO22X1 U1157 ( .IN1(n1426), .IN2(n852), .IN3(n1931), .IN4(\fpu_add_ctl/n37 ), 
        .Q(\fpu_add_frac_dp/n3737 ) );
  NOR2X0 U1158 ( .IN1(n1932), .IN2(n1933), .QN(n1931) );
  NAND3X0 U1159 ( .IN1(n1934), .IN2(n1935), .IN3(n1936), .QN(
        \fpu_add_frac_dp/n3736 ) );
  NAND2X0 U1160 ( .IN1(n1430), .IN2(n926), .QN(n1936) );
  AO22X1 U1161 ( .IN1(n1426), .IN2(n1264), .IN3(n1442), .IN4(n1937), .Q(
        \fpu_add_frac_dp/n3735 ) );
  NAND4X0 U1162 ( .IN1(n1938), .IN2(n1939), .IN3(n1940), .IN4(n1941), .QN(
        n1937) );
  NOR4X0 U1163 ( .IN1(n1942), .IN2(n1943), .IN3(n1944), .IN4(n1945), .QN(n1941) );
  AO222X1 U1164 ( .IN1(\fpu_add_frac_dp/n2399 ), .IN2(n1946), .IN3(n1947), 
        .IN4(n746), .IN5(n1948), .IN6(n166), .Q(n1943) );
  OR4X1 U1165 ( .IN1(n1949), .IN2(n1950), .IN3(n1951), .IN4(n1952), .Q(n1947)
         );
  NAND4X0 U1166 ( .IN1(n1953), .IN2(n1954), .IN3(n1955), .IN4(n1956), .QN(
        n1942) );
  NOR2X0 U1167 ( .IN1(n1957), .IN2(n1958), .QN(n1956) );
  INVX0 U1168 ( .INP(n1959), .ZN(n1955) );
  INVX0 U1169 ( .INP(n1960), .ZN(n1953) );
  NOR4X0 U1170 ( .IN1(n1961), .IN2(n1962), .IN3(n1963), .IN4(n1964), .QN(n1940) );
  OR3X1 U1171 ( .IN1(n1965), .IN2(n1966), .IN3(n1967), .Q(n1962) );
  OR4X1 U1172 ( .IN1(n1968), .IN2(n1969), .IN3(n1970), .IN4(n1971), .Q(n1961)
         );
  OR2X1 U1173 ( .IN1(n1972), .IN2(n1973), .Q(n1970) );
  NOR4X0 U1174 ( .IN1(n1974), .IN2(n1975), .IN3(n1976), .IN4(n1977), .QN(n1939) );
  OR3X1 U1175 ( .IN1(n1978), .IN2(n1979), .IN3(n1980), .Q(n1975) );
  OR4X1 U1176 ( .IN1(n1981), .IN2(n1982), .IN3(n1983), .IN4(n1984), .Q(n1974)
         );
  OR2X1 U1177 ( .IN1(n1985), .IN2(n1986), .Q(n1984) );
  NOR4X0 U1178 ( .IN1(n1987), .IN2(n1988), .IN3(n1989), .IN4(n1990), .QN(n1938) );
  OR3X1 U1179 ( .IN1(n1991), .IN2(n1992), .IN3(n1993), .Q(n1988) );
  OR4X1 U1180 ( .IN1(n1994), .IN2(n1995), .IN3(n1996), .IN4(n1997), .Q(n1987)
         );
  INVX0 U1181 ( .INP(n1998), .ZN(n1994) );
  AO22X1 U1182 ( .IN1(n1416), .IN2(n1302), .IN3(n1442), .IN4(n1999), .Q(
        \fpu_add_frac_dp/n3734 ) );
  NAND4X0 U1183 ( .IN1(n2000), .IN2(n2001), .IN3(n2002), .IN4(n2003), .QN(
        n1999) );
  OA222X1 U1184 ( .IN1(\fpu_add_frac_dp/n2308 ), .IN2(n2004), .IN3(n2005), 
        .IN4(n2006), .IN5(\fpu_add_frac_dp/n579 ), .IN6(n2007), .Q(n2003) );
  INVX0 U1185 ( .INP(n2008), .ZN(n2007) );
  OA22X1 U1186 ( .IN1(\fpu_add_frac_dp/n2377 ), .IN2(n2009), .IN3(
        \fpu_add_frac_dp/n580 ), .IN4(n2010), .Q(n2002) );
  NOR4X0 U1187 ( .IN1(n2011), .IN2(n2012), .IN3(n2013), .IN4(n2014), .QN(n2010) );
  NOR2X0 U1188 ( .IN1(n2015), .IN2(n2016), .QN(n2013) );
  AO222X1 U1189 ( .IN1(n2017), .IN2(n693), .IN3(n2018), .IN4(n2019), .IN5(
        n2020), .IN6(n2021), .Q(n2011) );
  NOR2X0 U1190 ( .IN1(\fpu_add_frac_dp/n2308 ), .IN2(n2022), .QN(n2018) );
  NAND3X0 U1191 ( .IN1(n2023), .IN2(n2024), .IN3(n2025), .QN(n2017) );
  AOI222X1 U1192 ( .IN1(n255), .IN2(n2026), .IN3(n2027), .IN4(n2021), .IN5(
        n1989), .IN6(n2028), .QN(n2025) );
  INVX0 U1193 ( .INP(n2029), .ZN(n2023) );
  OA221X1 U1194 ( .IN1(n2030), .IN2(n2016), .IN3(\fpu_add_frac_dp/n2308 ), 
        .IN4(n2031), .IN5(n2032), .Q(n2009) );
  AOI21X1 U1195 ( .IN1(n2021), .IN2(n2029), .IN3(n2033), .QN(n2032) );
  NAND2X0 U1196 ( .IN1(\fpu_add_frac_dp/n2306 ), .IN2(n2034), .QN(n2001) );
  NAND4X0 U1197 ( .IN1(n2035), .IN2(n2036), .IN3(n2037), .IN4(n2038), .QN(
        n2034) );
  OA22X1 U1198 ( .IN1(n2039), .IN2(n2016), .IN3(\fpu_add_frac_dp/n2308 ), 
        .IN4(n2040), .Q(n2037) );
  INVX0 U1199 ( .INP(n2041), .ZN(n2036) );
  INVX0 U1200 ( .INP(n2042), .ZN(n2035) );
  NAND2X0 U1201 ( .IN1(n2028), .IN2(n2043), .QN(n2000) );
  AO21X1 U1202 ( .IN1(n1397), .IN2(n1121), .IN3(n1319), .Q(
        \fpu_add_frac_dp/n3733 ) );
  AO22X1 U1203 ( .IN1(\fpu_add_frac_dp/n2369 ), .IN2(n1430), .IN3(n2044), 
        .IN4(n2045), .Q(\fpu_add_frac_dp/n3732 ) );
  INVX0 U1204 ( .INP(n1934), .ZN(n2044) );
  OAI221X1 U1205 ( .IN1(n1934), .IN2(n2045), .IN3(n2046), .IN4(
        \fpu_add_frac_dp/n5614 ), .IN5(n1935), .QN(\fpu_add_frac_dp/n3731 ) );
  NAND3X0 U1206 ( .IN1(n1435), .IN2(n649), .IN3(n2047), .QN(n1935) );
  MUX21X1 U1207 ( .IN1(n2048), .IN2(n2049), .S(n2050), .Q(n2045) );
  NAND3X0 U1208 ( .IN1(n2051), .IN2(n2052), .IN3(n2053), .QN(n2049) );
  INVX0 U1209 ( .INP(n2054), .ZN(n2053) );
  NAND2X0 U1210 ( .IN1(n2055), .IN2(n2056), .QN(n2048) );
  XOR2X1 U1211 ( .IN1(n2057), .IN2(n2058), .Q(n2056) );
  INVX0 U1212 ( .INP(n2059), .ZN(n2055) );
  NAND3X0 U1213 ( .IN1(n1737), .IN2(n1435), .IN3(n1656), .QN(n1934) );
  AO22X1 U1214 ( .IN1(n1417), .IN2(n652), .IN3(n2060), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3730 ) );
  XOR3X1 U1215 ( .IN1(\fpu_add_frac_dp/n2478 ), .IN2(\fpu_add_frac_dp/n2477 ), 
        .IN3(n2061), .Q(n2060) );
  AO22X1 U1216 ( .IN1(n1417), .IN2(n103), .IN3(n2062), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3729 ) );
  XOR3X1 U1217 ( .IN1(n625), .IN2(n2063), .IN3(n2064), .Q(n2062) );
  AO22X1 U1218 ( .IN1(n1417), .IN2(n282), .IN3(n2065), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3728 ) );
  XOR2X1 U1219 ( .IN1(n220), .IN2(n2066), .Q(n2065) );
  NOR2X0 U1220 ( .IN1(n2067), .IN2(n2068), .QN(n2066) );
  AO22X1 U1221 ( .IN1(n1417), .IN2(n671), .IN3(n1441), .IN4(n2069), .Q(
        \fpu_add_frac_dp/n3727 ) );
  XOR3X1 U1222 ( .IN1(n310), .IN2(n2070), .IN3(n2071), .Q(n2069) );
  AO22X1 U1223 ( .IN1(n1417), .IN2(n90), .IN3(n1442), .IN4(n2072), .Q(
        \fpu_add_frac_dp/n3726 ) );
  XOR3X1 U1224 ( .IN1(n2073), .IN2(n288), .IN3(n2074), .Q(n2072) );
  AO22X1 U1225 ( .IN1(n1417), .IN2(n626), .IN3(n2075), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3725 ) );
  XOR3X1 U1226 ( .IN1(n2076), .IN2(n223), .IN3(n2077), .Q(n2075) );
  AO22X1 U1227 ( .IN1(n1417), .IN2(n173), .IN3(n1442), .IN4(n2078), .Q(
        \fpu_add_frac_dp/n3724 ) );
  XOR3X1 U1228 ( .IN1(n2079), .IN2(n225), .IN3(n2080), .Q(n2078) );
  AO22X1 U1229 ( .IN1(n1417), .IN2(n33), .IN3(n2081), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3723 ) );
  XOR3X1 U1230 ( .IN1(n2082), .IN2(n222), .IN3(n2083), .Q(n2081) );
  AO22X1 U1231 ( .IN1(n1418), .IN2(n623), .IN3(n1441), .IN4(n2084), .Q(
        \fpu_add_frac_dp/n3722 ) );
  XOR3X1 U1232 ( .IN1(n2085), .IN2(n224), .IN3(n2086), .Q(n2084) );
  AO22X1 U1233 ( .IN1(n1418), .IN2(n34), .IN3(n2087), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3721 ) );
  XOR3X1 U1234 ( .IN1(n261), .IN2(n2088), .IN3(n2089), .Q(n2087) );
  AO22X1 U1235 ( .IN1(n1417), .IN2(n12), .IN3(n2090), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3720 ) );
  XOR3X1 U1236 ( .IN1(n260), .IN2(n2091), .IN3(n2092), .Q(n2090) );
  AO22X1 U1237 ( .IN1(n1417), .IN2(n691), .IN3(n2093), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3719 ) );
  XOR3X1 U1238 ( .IN1(n253), .IN2(n2094), .IN3(n2095), .Q(n2093) );
  AO22X1 U1239 ( .IN1(n1417), .IN2(n37), .IN3(n2096), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3718 ) );
  XOR3X1 U1240 ( .IN1(n252), .IN2(n2097), .IN3(n2098), .Q(n2096) );
  AO22X1 U1241 ( .IN1(n1417), .IN2(n597), .IN3(n1441), .IN4(n2099), .Q(
        \fpu_add_frac_dp/n3717 ) );
  AO22X1 U1242 ( .IN1(n2100), .IN2(n2101), .IN3(n2102), .IN4(n327), .Q(n2099)
         );
  NAND2X0 U1243 ( .IN1(n2103), .IN2(n2101), .QN(n2102) );
  INVX0 U1244 ( .INP(n2104), .ZN(n2100) );
  AO22X1 U1245 ( .IN1(\fpu_add_frac_dp/n2330 ), .IN2(n1430), .IN3(n2105), 
        .IN4(n1440), .Q(\fpu_add_frac_dp/n3716 ) );
  XOR2X1 U1246 ( .IN1(n180), .IN2(n2106), .Q(n2105) );
  AND2X1 U1247 ( .IN1(n2107), .IN2(n2108), .Q(n2106) );
  AO22X1 U1248 ( .IN1(\fpu_add_frac_dp/n2400 ), .IN2(n1419), .IN3(n2109), 
        .IN4(n1440), .Q(\fpu_add_frac_dp/n3715 ) );
  XOR2X1 U1249 ( .IN1(n268), .IN2(n2110), .Q(n2109) );
  NOR2X0 U1250 ( .IN1(n2111), .IN2(n2112), .QN(n2110) );
  INVX0 U1251 ( .INP(n2113), .ZN(n2111) );
  AO22X1 U1252 ( .IN1(n1417), .IN2(n328), .IN3(n2114), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3714 ) );
  XOR2X1 U1253 ( .IN1(n179), .IN2(n2115), .Q(n2114) );
  OA21X1 U1254 ( .IN1(n2116), .IN2(n2117), .IN3(n2118), .Q(n2115) );
  AO22X1 U1255 ( .IN1(n1418), .IN2(n43), .IN3(n1441), .IN4(n2119), .Q(
        \fpu_add_frac_dp/n3713 ) );
  XOR3X1 U1256 ( .IN1(n251), .IN2(n2120), .IN3(n2121), .Q(n2119) );
  AO22X1 U1257 ( .IN1(n1418), .IN2(n111), .IN3(n2122), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3712 ) );
  XOR3X1 U1258 ( .IN1(n250), .IN2(n2123), .IN3(n2124), .Q(n2122) );
  AO22X1 U1259 ( .IN1(n1418), .IN2(n664), .IN3(n2125), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3711 ) );
  XOR3X1 U1260 ( .IN1(n249), .IN2(n2126), .IN3(n2127), .Q(n2125) );
  AO22X1 U1261 ( .IN1(\fpu_add_frac_dp/n2339 ), .IN2(n1430), .IN3(n2128), 
        .IN4(n1440), .Q(\fpu_add_frac_dp/n3710 ) );
  XOR2X1 U1262 ( .IN1(n263), .IN2(n2129), .Q(n2128) );
  AND2X1 U1263 ( .IN1(n2130), .IN2(n2131), .Q(n2129) );
  AO22X1 U1264 ( .IN1(\fpu_add_frac_dp/n2405 ), .IN2(n1430), .IN3(n2132), 
        .IN4(n1440), .Q(\fpu_add_frac_dp/n3709 ) );
  XOR2X1 U1265 ( .IN1(n267), .IN2(n2133), .Q(n2132) );
  NOR2X0 U1266 ( .IN1(n2134), .IN2(n2135), .QN(n2133) );
  INVX0 U1267 ( .INP(n2136), .ZN(n2134) );
  AO22X1 U1268 ( .IN1(n1418), .IN2(n594), .IN3(n1441), .IN4(n2137), .Q(
        \fpu_add_frac_dp/n3708 ) );
  XOR3X1 U1269 ( .IN1(n2138), .IN2(n279), .IN3(n2139), .Q(n2137) );
  AO22X1 U1270 ( .IN1(n1418), .IN2(n74), .IN3(n2140), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3707 ) );
  XOR3X1 U1271 ( .IN1(\fpu_add_frac_dp/n814 ), .IN2(n2141), .IN3(n2142), .Q(
        n2140) );
  AO22X1 U1272 ( .IN1(n1418), .IN2(n331), .IN3(n2143), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3706 ) );
  XOR3X1 U1273 ( .IN1(n248), .IN2(n2144), .IN3(n2145), .Q(n2143) );
  AO22X1 U1274 ( .IN1(n1418), .IN2(n116), .IN3(n2146), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3705 ) );
  XOR3X1 U1275 ( .IN1(n247), .IN2(n2147), .IN3(n2148), .Q(n2146) );
  AO22X1 U1276 ( .IN1(\fpu_add_frac_dp/n2402 ), .IN2(n1430), .IN3(n2149), 
        .IN4(n1439), .Q(\fpu_add_frac_dp/n3704 ) );
  XOR3X1 U1277 ( .IN1(n246), .IN2(n2150), .IN3(n2151), .Q(n2149) );
  AO22X1 U1278 ( .IN1(\fpu_add_frac_dp/n2313 ), .IN2(n1430), .IN3(n2152), 
        .IN4(n1440), .Q(\fpu_add_frac_dp/n3703 ) );
  XOR2X1 U1279 ( .IN1(n204), .IN2(n2153), .Q(n2152) );
  NOR2X0 U1280 ( .IN1(n2154), .IN2(n2155), .QN(n2153) );
  AO22X1 U1281 ( .IN1(n1418), .IN2(n329), .IN3(n1441), .IN4(n2156), .Q(
        \fpu_add_frac_dp/n3702 ) );
  XOR3X1 U1282 ( .IN1(n245), .IN2(n2157), .IN3(n2158), .Q(n2156) );
  AO22X1 U1283 ( .IN1(n1418), .IN2(n101), .IN3(n2159), .IN4(n1440), .Q(
        \fpu_add_frac_dp/n3701 ) );
  XOR3X1 U1284 ( .IN1(n244), .IN2(n2160), .IN3(n2161), .Q(n2159) );
  AO22X1 U1285 ( .IN1(n1418), .IN2(n262), .IN3(n2162), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3700 ) );
  XOR2X1 U1286 ( .IN1(n203), .IN2(n2163), .Q(n2162) );
  NOR2X0 U1287 ( .IN1(n2164), .IN2(n2165), .QN(n2163) );
  AO22X1 U1288 ( .IN1(\fpu_add_frac_dp/n2335 ), .IN2(n1430), .IN3(n1441), 
        .IN4(n2166), .Q(\fpu_add_frac_dp/n3699 ) );
  XOR3X1 U1289 ( .IN1(n243), .IN2(n2167), .IN3(n2168), .Q(n2166) );
  AO22X1 U1290 ( .IN1(\fpu_add_frac_dp/n2403 ), .IN2(n1430), .IN3(n2169), 
        .IN4(n1439), .Q(\fpu_add_frac_dp/n3698 ) );
  XOR3X1 U1291 ( .IN1(n242), .IN2(n2170), .IN3(n2171), .Q(n2169) );
  AO22X1 U1292 ( .IN1(\fpu_add_frac_dp/n2342 ), .IN2(n1418), .IN3(n2172), 
        .IN4(n1438), .Q(\fpu_add_frac_dp/n3697 ) );
  XOR3X1 U1293 ( .IN1(n241), .IN2(n2173), .IN3(n2174), .Q(n2172) );
  AO22X1 U1294 ( .IN1(\fpu_add_frac_dp/n2289 ), .IN2(n1430), .IN3(n2175), 
        .IN4(n1439), .Q(\fpu_add_frac_dp/n3696 ) );
  XOR3X1 U1295 ( .IN1(n240), .IN2(n2176), .IN3(n2177), .Q(n2175) );
  AO22X1 U1296 ( .IN1(\fpu_add_frac_dp/n2406 ), .IN2(n1417), .IN3(n2178), 
        .IN4(n1439), .Q(\fpu_add_frac_dp/n3695 ) );
  XOR2X1 U1297 ( .IN1(n202), .IN2(n2179), .Q(n2178) );
  NOR2X0 U1298 ( .IN1(n2180), .IN2(n2181), .QN(n2179) );
  AO22X1 U1299 ( .IN1(\fpu_add_frac_dp/n2332 ), .IN2(n1430), .IN3(n1441), 
        .IN4(n2182), .Q(\fpu_add_frac_dp/n3694 ) );
  XOR3X1 U1300 ( .IN1(n239), .IN2(n2183), .IN3(n2184), .Q(n2182) );
  AO22X1 U1301 ( .IN1(n1419), .IN2(n177), .IN3(n2185), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3693 ) );
  XOR2X1 U1302 ( .IN1(n201), .IN2(n2186), .Q(n2185) );
  NOR2X0 U1303 ( .IN1(n2187), .IN2(n2188), .QN(n2186) );
  AO22X1 U1304 ( .IN1(n1419), .IN2(n86), .IN3(n1441), .IN4(n2189), .Q(
        \fpu_add_frac_dp/n3692 ) );
  XOR3X1 U1305 ( .IN1(n238), .IN2(n2190), .IN3(n2191), .Q(n2189) );
  AO22X1 U1306 ( .IN1(n1419), .IN2(n19), .IN3(n2192), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3691 ) );
  XOR2X1 U1307 ( .IN1(n200), .IN2(n2193), .Q(n2192) );
  NOR2X0 U1308 ( .IN1(n2194), .IN2(n2195), .QN(n2193) );
  AO22X1 U1309 ( .IN1(n1419), .IN2(n673), .IN3(n1441), .IN4(n2196), .Q(
        \fpu_add_frac_dp/n3690 ) );
  XOR3X1 U1310 ( .IN1(n259), .IN2(n2197), .IN3(n2198), .Q(n2196) );
  AO22X1 U1311 ( .IN1(n1419), .IN2(n117), .IN3(n2199), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3689 ) );
  XOR3X1 U1312 ( .IN1(n237), .IN2(n2200), .IN3(n2201), .Q(n2199) );
  AO22X1 U1313 ( .IN1(n1419), .IN2(n38), .IN3(n2202), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3688 ) );
  XOR2X1 U1314 ( .IN1(n199), .IN2(n2203), .Q(n2202) );
  NOR2X0 U1315 ( .IN1(n2204), .IN2(n2205), .QN(n2203) );
  AO22X1 U1316 ( .IN1(n1420), .IN2(n83), .IN3(n1441), .IN4(n2206), .Q(
        \fpu_add_frac_dp/n3687 ) );
  XOR3X1 U1317 ( .IN1(n236), .IN2(n2207), .IN3(n2208), .Q(n2206) );
  AO22X1 U1318 ( .IN1(n1420), .IN2(n665), .IN3(n2209), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3686 ) );
  XOR3X1 U1319 ( .IN1(n235), .IN2(n2210), .IN3(n2211), .Q(n2209) );
  AO22X1 U1320 ( .IN1(n1420), .IN2(n100), .IN3(n2212), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3685 ) );
  XOR3X1 U1321 ( .IN1(n234), .IN2(n2213), .IN3(n2214), .Q(n2212) );
  AO22X1 U1322 ( .IN1(n1420), .IN2(n667), .IN3(n2215), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3684 ) );
  XOR2X1 U1323 ( .IN1(n198), .IN2(n2216), .Q(n2215) );
  NOR2X0 U1324 ( .IN1(n2217), .IN2(n2218), .QN(n2216) );
  AO22X1 U1325 ( .IN1(n1420), .IN2(n40), .IN3(n2219), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3683 ) );
  XOR2X1 U1326 ( .IN1(n197), .IN2(n2220), .Q(n2219) );
  NOR2X0 U1327 ( .IN1(n2221), .IN2(n2222), .QN(n2220) );
  AO22X1 U1328 ( .IN1(n1420), .IN2(n104), .IN3(n1441), .IN4(n2223), .Q(
        \fpu_add_frac_dp/n3682 ) );
  XOR3X1 U1329 ( .IN1(n233), .IN2(n2224), .IN3(n2225), .Q(n2223) );
  AO22X1 U1330 ( .IN1(n1420), .IN2(n175), .IN3(n2226), .IN4(n1439), .Q(
        \fpu_add_frac_dp/n3681 ) );
  XOR3X1 U1331 ( .IN1(n232), .IN2(n2227), .IN3(n2228), .Q(n2226) );
  AO22X1 U1332 ( .IN1(n1420), .IN2(n22), .IN3(n2229), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3680 ) );
  XOR3X1 U1333 ( .IN1(n231), .IN2(n2230), .IN3(n2231), .Q(n2229) );
  AO22X1 U1334 ( .IN1(n1420), .IN2(n85), .IN3(n2232), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3679 ) );
  XOR3X1 U1335 ( .IN1(n230), .IN2(n2233), .IN3(n2234), .Q(n2232) );
  AO22X1 U1336 ( .IN1(n1420), .IN2(n313), .IN3(n2235), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3678 ) );
  XOR3X1 U1337 ( .IN1(n229), .IN2(n2236), .IN3(n2237), .Q(n2235) );
  AO22X1 U1338 ( .IN1(n1420), .IN2(n92), .IN3(n2238), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3677 ) );
  XOR3X1 U1339 ( .IN1(n228), .IN2(n2239), .IN3(n2240), .Q(n2238) );
  AO22X1 U1340 ( .IN1(n1420), .IN2(n265), .IN3(n2241), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3676 ) );
  XOR3X1 U1341 ( .IN1(n227), .IN2(n2242), .IN3(n2243), .Q(n2241) );
  AO22X1 U1342 ( .IN1(\fpu_add_frac_dp/n2338 ), .IN2(n1430), .IN3(n2244), 
        .IN4(n1438), .Q(\fpu_add_frac_dp/n3675 ) );
  XOR2X1 U1343 ( .IN1(n196), .IN2(n2245), .Q(n2244) );
  NOR2X0 U1344 ( .IN1(n2246), .IN2(n2247), .QN(n2245) );
  AO22X1 U1345 ( .IN1(\fpu_add_frac_dp/n2407 ), .IN2(n1430), .IN3(n1441), 
        .IN4(n2248), .Q(\fpu_add_frac_dp/n3674 ) );
  XOR3X1 U1346 ( .IN1(n294), .IN2(n2249), .IN3(n2250), .Q(n2248) );
  AO22X1 U1347 ( .IN1(\fpu_add_frac_dp/n2343 ), .IN2(n1430), .IN3(n2251), 
        .IN4(n1438), .Q(\fpu_add_frac_dp/n3673 ) );
  XOR2X1 U1348 ( .IN1(n2252), .IN2(\fpu_add_frac_dp/n780 ), .Q(n2251) );
  NAND2X0 U1349 ( .IN1(n2253), .IN2(n2254), .QN(n2252) );
  INVX0 U1350 ( .INP(n2255), .ZN(n2253) );
  AO22X1 U1351 ( .IN1(n1420), .IN2(n171), .IN3(n1441), .IN4(n2256), .Q(
        \fpu_add_frac_dp/n3672 ) );
  AO22X1 U1352 ( .IN1(n2257), .IN2(n334), .IN3(n2258), .IN4(n2259), .Q(n2256)
         );
  NAND2X0 U1353 ( .IN1(n2260), .IN2(n2261), .QN(n2259) );
  XNOR2X1 U1354 ( .IN1(n2261), .IN2(n2260), .Q(n2257) );
  AO22X1 U1355 ( .IN1(n1420), .IN2(n82), .IN3(n1441), .IN4(n2262), .Q(
        \fpu_add_frac_dp/n3671 ) );
  XOR3X1 U1356 ( .IN1(n293), .IN2(n2263), .IN3(n2264), .Q(n2262) );
  AO22X1 U1357 ( .IN1(\fpu_add_frac_dp/n2337 ), .IN2(n1420), .IN3(n2265), 
        .IN4(n1438), .Q(\fpu_add_frac_dp/n3670 ) );
  XOR3X1 U1358 ( .IN1(\fpu_add_frac_dp/n777 ), .IN2(n2266), .IN3(n2267), .Q(
        n2265) );
  AO22X1 U1359 ( .IN1(n1420), .IN2(n94), .IN3(n2268), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3669 ) );
  XOR2X1 U1360 ( .IN1(n195), .IN2(n2269), .Q(n2268) );
  NOR2X0 U1361 ( .IN1(n2270), .IN2(n2271), .QN(n2269) );
  AO22X1 U1362 ( .IN1(n1421), .IN2(n266), .IN3(n1441), .IN4(n2272), .Q(
        \fpu_add_frac_dp/n3668 ) );
  XOR3X1 U1363 ( .IN1(n226), .IN2(n2273), .IN3(n2274), .Q(n2272) );
  AO22X1 U1364 ( .IN1(n1422), .IN2(n87), .IN3(n1441), .IN4(n2275), .Q(
        \fpu_add_frac_dp/n3667 ) );
  XOR3X1 U1365 ( .IN1(\fpu_add_frac_dp/n5640 ), .IN2(n2276), .IN3(n2277), .Q(
        n2275) );
  NOR2X0 U1366 ( .IN1(\fpu_add_frac_dp/n2369 ), .IN2(n2278), .QN(n2277) );
  MUX21X1 U1367 ( .IN1(n1324), .IN2(n1328), .S(\fpu_add_frac_dp/n2498 ), .Q(
        n2278) );
  OA22X1 U1368 ( .IN1(n2279), .IN2(n226), .IN3(n2280), .IN4(n2281), .Q(n2276)
         );
  NOR2X0 U1369 ( .IN1(n2273), .IN2(n2274), .QN(n2279) );
  INVX0 U1370 ( .INP(n2280), .ZN(n2274) );
  OA21X1 U1371 ( .IN1(n195), .IN2(n2270), .IN3(n2282), .Q(n2280) );
  INVX0 U1372 ( .INP(n2271), .ZN(n2282) );
  NOR2X0 U1373 ( .IN1(n2283), .IN2(n2284), .QN(n2271) );
  AND2X1 U1374 ( .IN1(n2283), .IN2(n2284), .Q(n2270) );
  AO21X1 U1375 ( .IN1(\fpu_add_frac_dp/n2502 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2285), .Q(n2284) );
  MUX21X1 U1376 ( .IN1(n1323), .IN2(n1327), .S(\fpu_add_frac_dp/n2506 ), .Q(
        n2285) );
  AO22X1 U1377 ( .IN1(n2267), .IN2(n2286), .IN3(n2287), .IN4(n317), .Q(n2283)
         );
  NAND2X0 U1378 ( .IN1(n2288), .IN2(n2266), .QN(n2287) );
  INVX0 U1379 ( .INP(n2286), .ZN(n2266) );
  AO21X1 U1380 ( .IN1(\fpu_add_frac_dp/n2506 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2289), .Q(n2286) );
  MUX21X1 U1381 ( .IN1(n1327), .IN2(n1324), .S(\fpu_add_frac_dp/n2384 ), .Q(
        n2289) );
  INVX0 U1382 ( .INP(n2288), .ZN(n2267) );
  OA22X1 U1383 ( .IN1(n2264), .IN2(n2263), .IN3(n2290), .IN4(
        \fpu_add_frac_dp/n778 ), .Q(n2288) );
  AND2X1 U1384 ( .IN1(n2263), .IN2(n2264), .Q(n2290) );
  AOI21X1 U1385 ( .IN1(\fpu_add_frac_dp/n2369 ), .IN2(n1009), .IN3(n2291), 
        .QN(n2263) );
  MUX21X1 U1386 ( .IN1(n64), .IN2(n1323), .S(\fpu_add_frac_dp/n2391 ), .Q(
        n2291) );
  AO21X1 U1387 ( .IN1(n2260), .IN2(n2261), .IN3(n2258), .Q(n2264) );
  OA21X1 U1388 ( .IN1(n2261), .IN2(n2260), .IN3(\fpu_add_frac_dp/n779 ), .Q(
        n2258) );
  OAI21X1 U1389 ( .IN1(n332), .IN2(n2255), .IN3(n2254), .QN(n2261) );
  NAND2X0 U1390 ( .IN1(n2292), .IN2(n2293), .QN(n2254) );
  NOR2X0 U1391 ( .IN1(n2293), .IN2(n2292), .QN(n2255) );
  AOI21X1 U1392 ( .IN1(\fpu_add_frac_dp/n2369 ), .IN2(n561), .IN3(n2294), .QN(
        n2292) );
  MUX21X1 U1393 ( .IN1(n1328), .IN2(n155), .S(\fpu_add_frac_dp/n2392 ), .Q(
        n2294) );
  AO22X1 U1394 ( .IN1(n2249), .IN2(n2250), .IN3(\fpu_add_frac_dp/n781 ), .IN4(
        n2295), .Q(n2293) );
  NAND2X0 U1395 ( .IN1(n2296), .IN2(n2297), .QN(n2295) );
  INVX0 U1396 ( .INP(n2296), .ZN(n2250) );
  OA21X1 U1397 ( .IN1(n196), .IN2(n2246), .IN3(n2298), .Q(n2296) );
  INVX0 U1398 ( .INP(n2247), .ZN(n2298) );
  NOR2X0 U1399 ( .IN1(n2299), .IN2(n2300), .QN(n2247) );
  AND2X1 U1400 ( .IN1(n2299), .IN2(n2300), .Q(n2246) );
  AO21X1 U1401 ( .IN1(\fpu_add_frac_dp/n2357 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2301), .Q(n2300) );
  MUX21X1 U1402 ( .IN1(n155), .IN2(n64), .S(\fpu_add_frac_dp/n2431 ), .Q(n2301) );
  AO22X1 U1403 ( .IN1(n2243), .IN2(n2242), .IN3(n2302), .IN4(n227), .Q(n2299)
         );
  OR2X1 U1404 ( .IN1(n2243), .IN2(n2242), .Q(n2302) );
  AO21X1 U1405 ( .IN1(\fpu_add_frac_dp/n2431 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2303), .Q(n2242) );
  MUX21X1 U1406 ( .IN1(n1325), .IN2(n1328), .S(\fpu_add_frac_dp/n2418 ), .Q(
        n2303) );
  AO22X1 U1407 ( .IN1(n2240), .IN2(n2239), .IN3(n2304), .IN4(n228), .Q(n2243)
         );
  OR2X1 U1408 ( .IN1(n2240), .IN2(n2239), .Q(n2304) );
  AO21X1 U1409 ( .IN1(\fpu_add_frac_dp/n2418 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2305), .Q(n2239) );
  MUX21X1 U1410 ( .IN1(n1324), .IN2(n1327), .S(\fpu_add_frac_dp/n2351 ), .Q(
        n2305) );
  AO22X1 U1411 ( .IN1(n2237), .IN2(n2236), .IN3(n2306), .IN4(n229), .Q(n2240)
         );
  OR2X1 U1412 ( .IN1(n2237), .IN2(n2236), .Q(n2306) );
  AO21X1 U1413 ( .IN1(\fpu_add_frac_dp/n2351 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2307), .Q(n2236) );
  MUX21X1 U1414 ( .IN1(n1323), .IN2(n64), .S(\fpu_add_frac_dp/n2505 ), .Q(
        n2307) );
  AO22X1 U1415 ( .IN1(n2234), .IN2(n2233), .IN3(n2308), .IN4(n230), .Q(n2237)
         );
  OR2X1 U1416 ( .IN1(n2234), .IN2(n2233), .Q(n2308) );
  AO21X1 U1417 ( .IN1(\fpu_add_frac_dp/n2505 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2309), .Q(n2233) );
  MUX21X1 U1418 ( .IN1(n155), .IN2(n1328), .S(\fpu_add_frac_dp/n2501 ), .Q(
        n2309) );
  AO22X1 U1419 ( .IN1(n2231), .IN2(n2230), .IN3(n2310), .IN4(n231), .Q(n2234)
         );
  OR2X1 U1420 ( .IN1(n2231), .IN2(n2230), .Q(n2310) );
  AO21X1 U1421 ( .IN1(\fpu_add_frac_dp/n2501 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2311), .Q(n2230) );
  MUX21X1 U1422 ( .IN1(n1325), .IN2(n1327), .S(\fpu_add_frac_dp/n2512 ), .Q(
        n2311) );
  AO22X1 U1423 ( .IN1(n2228), .IN2(n2227), .IN3(n2312), .IN4(n232), .Q(n2231)
         );
  OR2X1 U1424 ( .IN1(n2228), .IN2(n2227), .Q(n2312) );
  AO21X1 U1425 ( .IN1(\fpu_add_frac_dp/n2512 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2313), .Q(n2227) );
  MUX21X1 U1426 ( .IN1(n1324), .IN2(n64), .S(\fpu_add_frac_dp/n2509 ), .Q(
        n2313) );
  AO22X1 U1427 ( .IN1(n2314), .IN2(n2315), .IN3(n2316), .IN4(n233), .Q(n2228)
         );
  NAND2X0 U1428 ( .IN1(n2224), .IN2(n2225), .QN(n2316) );
  INVX0 U1429 ( .INP(n2314), .ZN(n2225) );
  INVX0 U1430 ( .INP(n2315), .ZN(n2224) );
  AO21X1 U1431 ( .IN1(\fpu_add_frac_dp/n2509 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2317), .Q(n2315) );
  MUX21X1 U1432 ( .IN1(n1323), .IN2(n1328), .S(\fpu_add_frac_dp/n2500 ), .Q(
        n2317) );
  OA21X1 U1433 ( .IN1(n197), .IN2(n2221), .IN3(n2318), .Q(n2314) );
  INVX0 U1434 ( .INP(n2222), .ZN(n2318) );
  NOR2X0 U1435 ( .IN1(n2319), .IN2(n2320), .QN(n2222) );
  AND2X1 U1436 ( .IN1(n2320), .IN2(n2319), .Q(n2221) );
  AO21X1 U1437 ( .IN1(\fpu_add_frac_dp/n2500 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2321), .Q(n2319) );
  MUX21X1 U1438 ( .IN1(n155), .IN2(n1327), .S(\fpu_add_frac_dp/n2303 ), .Q(
        n2321) );
  OA21X1 U1439 ( .IN1(n198), .IN2(n2217), .IN3(n2322), .Q(n2320) );
  INVX0 U1440 ( .INP(n2218), .ZN(n2322) );
  NOR2X0 U1441 ( .IN1(n2323), .IN2(n2324), .QN(n2218) );
  AND2X1 U1442 ( .IN1(n2323), .IN2(n2324), .Q(n2217) );
  AO21X1 U1443 ( .IN1(\fpu_add_frac_dp/n2303 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2325), .Q(n2324) );
  MUX21X1 U1444 ( .IN1(n1325), .IN2(n64), .S(\fpu_add_frac_dp/n2356 ), .Q(
        n2325) );
  AO22X1 U1445 ( .IN1(n2214), .IN2(n2213), .IN3(n2326), .IN4(n234), .Q(n2323)
         );
  OR2X1 U1446 ( .IN1(n2214), .IN2(n2213), .Q(n2326) );
  AO21X1 U1447 ( .IN1(\fpu_add_frac_dp/n2356 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2327), .Q(n2213) );
  MUX21X1 U1448 ( .IN1(n1324), .IN2(n1328), .S(\fpu_add_frac_dp/n2508 ), .Q(
        n2327) );
  AO22X1 U1449 ( .IN1(n2211), .IN2(n2210), .IN3(n2328), .IN4(n235), .Q(n2214)
         );
  OR2X1 U1450 ( .IN1(n2211), .IN2(n2210), .Q(n2328) );
  AO21X1 U1451 ( .IN1(\fpu_add_frac_dp/n2508 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2329), .Q(n2210) );
  MUX21X1 U1452 ( .IN1(n1323), .IN2(n1327), .S(\fpu_add_frac_dp/n2504 ), .Q(
        n2329) );
  AO22X1 U1453 ( .IN1(n2330), .IN2(n2331), .IN3(n2332), .IN4(n236), .Q(n2211)
         );
  NAND2X0 U1454 ( .IN1(n2207), .IN2(n2208), .QN(n2332) );
  INVX0 U1455 ( .INP(n2330), .ZN(n2208) );
  INVX0 U1456 ( .INP(n2331), .ZN(n2207) );
  AO21X1 U1457 ( .IN1(\fpu_add_frac_dp/n2504 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2333), .Q(n2331) );
  MUX21X1 U1458 ( .IN1(n155), .IN2(n64), .S(\fpu_add_frac_dp/n2276 ), .Q(n2333) );
  OA21X1 U1459 ( .IN1(n199), .IN2(n2204), .IN3(n2334), .Q(n2330) );
  INVX0 U1460 ( .INP(n2205), .ZN(n2334) );
  NOR2X0 U1461 ( .IN1(n2335), .IN2(n2336), .QN(n2205) );
  AND2X1 U1462 ( .IN1(n2335), .IN2(n2336), .Q(n2204) );
  AO21X1 U1463 ( .IN1(\fpu_add_frac_dp/n2276 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2337), .Q(n2336) );
  MUX21X1 U1464 ( .IN1(n1325), .IN2(n1328), .S(\fpu_add_frac_dp/n2302 ), .Q(
        n2337) );
  AO22X1 U1465 ( .IN1(n2201), .IN2(n2200), .IN3(n2338), .IN4(n237), .Q(n2335)
         );
  OR2X1 U1466 ( .IN1(n2201), .IN2(n2200), .Q(n2338) );
  AO21X1 U1467 ( .IN1(\fpu_add_frac_dp/n2302 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2339), .Q(n2200) );
  MUX21X1 U1468 ( .IN1(n1324), .IN2(n1327), .S(\fpu_add_frac_dp/n2422 ), .Q(
        n2339) );
  AO22X1 U1469 ( .IN1(n2340), .IN2(n2341), .IN3(n2342), .IN4(n259), .Q(n2201)
         );
  NAND2X0 U1470 ( .IN1(n2197), .IN2(n2198), .QN(n2342) );
  INVX0 U1471 ( .INP(n2340), .ZN(n2198) );
  INVX0 U1472 ( .INP(n2341), .ZN(n2197) );
  AO21X1 U1473 ( .IN1(\fpu_add_frac_dp/n2422 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2343), .Q(n2341) );
  MUX21X1 U1474 ( .IN1(n1323), .IN2(n64), .S(\fpu_add_frac_dp/n2355 ), .Q(
        n2343) );
  OA21X1 U1475 ( .IN1(n200), .IN2(n2194), .IN3(n2344), .Q(n2340) );
  INVX0 U1476 ( .INP(n2195), .ZN(n2344) );
  NOR2X0 U1477 ( .IN1(n2345), .IN2(n2346), .QN(n2195) );
  AND2X1 U1478 ( .IN1(n2345), .IN2(n2346), .Q(n2194) );
  AO21X1 U1479 ( .IN1(\fpu_add_frac_dp/n2355 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2347), .Q(n2346) );
  MUX21X1 U1480 ( .IN1(n155), .IN2(n1328), .S(\fpu_add_frac_dp/n2275 ), .Q(
        n2347) );
  AO22X1 U1481 ( .IN1(n2348), .IN2(n2349), .IN3(n2350), .IN4(n238), .Q(n2345)
         );
  NAND2X0 U1482 ( .IN1(n2190), .IN2(n2191), .QN(n2350) );
  INVX0 U1483 ( .INP(n2348), .ZN(n2191) );
  INVX0 U1484 ( .INP(n2349), .ZN(n2190) );
  AO21X1 U1485 ( .IN1(\fpu_add_frac_dp/n2275 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2351), .Q(n2349) );
  MUX21X1 U1486 ( .IN1(n1325), .IN2(n1327), .S(\fpu_add_frac_dp/n2301 ), .Q(
        n2351) );
  OA21X1 U1487 ( .IN1(n201), .IN2(n2187), .IN3(n2352), .Q(n2348) );
  INVX0 U1488 ( .INP(n2188), .ZN(n2352) );
  NOR2X0 U1489 ( .IN1(n2353), .IN2(n2354), .QN(n2188) );
  AND2X1 U1490 ( .IN1(n2353), .IN2(n2354), .Q(n2187) );
  AO21X1 U1491 ( .IN1(\fpu_add_frac_dp/n2301 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2355), .Q(n2354) );
  MUX21X1 U1492 ( .IN1(n1324), .IN2(n64), .S(\fpu_add_frac_dp/n2421 ), .Q(
        n2355) );
  AO22X1 U1493 ( .IN1(n2356), .IN2(n2357), .IN3(n2358), .IN4(n239), .Q(n2353)
         );
  NAND2X0 U1494 ( .IN1(n2183), .IN2(n2184), .QN(n2358) );
  INVX0 U1495 ( .INP(n2356), .ZN(n2184) );
  INVX0 U1496 ( .INP(n2357), .ZN(n2183) );
  AO21X1 U1497 ( .IN1(\fpu_add_frac_dp/n2421 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2359), .Q(n2357) );
  MUX21X1 U1498 ( .IN1(n1323), .IN2(n1328), .S(\fpu_add_frac_dp/n2511 ), .Q(
        n2359) );
  OA21X1 U1499 ( .IN1(n202), .IN2(n2180), .IN3(n2360), .Q(n2356) );
  INVX0 U1500 ( .INP(n2181), .ZN(n2360) );
  NOR2X0 U1501 ( .IN1(n2361), .IN2(n2362), .QN(n2181) );
  AND2X1 U1502 ( .IN1(n2361), .IN2(n2362), .Q(n2180) );
  AO21X1 U1503 ( .IN1(\fpu_add_frac_dp/n2511 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2363), .Q(n2362) );
  MUX21X1 U1504 ( .IN1(n155), .IN2(n1327), .S(\fpu_add_frac_dp/n2435 ), .Q(
        n2363) );
  AO22X1 U1505 ( .IN1(n2177), .IN2(n2176), .IN3(n2364), .IN4(n240), .Q(n2361)
         );
  OR2X1 U1506 ( .IN1(n2177), .IN2(n2176), .Q(n2364) );
  AO21X1 U1507 ( .IN1(\fpu_add_frac_dp/n2435 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2365), .Q(n2176) );
  MUX21X1 U1508 ( .IN1(n1325), .IN2(n64), .S(\fpu_add_frac_dp/n2354 ), .Q(
        n2365) );
  AO22X1 U1509 ( .IN1(n2174), .IN2(n2173), .IN3(n2366), .IN4(n241), .Q(n2177)
         );
  OR2X1 U1510 ( .IN1(n2174), .IN2(n2173), .Q(n2366) );
  AO21X1 U1511 ( .IN1(\fpu_add_frac_dp/n2354 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2367), .Q(n2173) );
  MUX21X1 U1512 ( .IN1(n1324), .IN2(n1328), .S(\fpu_add_frac_dp/n2274 ), .Q(
        n2367) );
  AO22X1 U1513 ( .IN1(n2171), .IN2(n2170), .IN3(n2368), .IN4(n242), .Q(n2174)
         );
  OR2X1 U1514 ( .IN1(n2171), .IN2(n2170), .Q(n2368) );
  AO21X1 U1515 ( .IN1(\fpu_add_frac_dp/n2274 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2369), .Q(n2170) );
  MUX21X1 U1516 ( .IN1(n1323), .IN2(n1327), .S(\fpu_add_frac_dp/n2300 ), .Q(
        n2369) );
  AO22X1 U1517 ( .IN1(n2370), .IN2(n2371), .IN3(n2372), .IN4(n243), .Q(n2171)
         );
  NAND2X0 U1518 ( .IN1(n2167), .IN2(n2168), .QN(n2372) );
  INVX0 U1519 ( .INP(n2370), .ZN(n2168) );
  INVX0 U1520 ( .INP(n2371), .ZN(n2167) );
  AO21X1 U1521 ( .IN1(\fpu_add_frac_dp/n2300 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2373), .Q(n2371) );
  MUX21X1 U1522 ( .IN1(n155), .IN2(n64), .S(\fpu_add_frac_dp/n2510 ), .Q(n2373) );
  OA21X1 U1523 ( .IN1(n203), .IN2(n2164), .IN3(n2374), .Q(n2370) );
  INVX0 U1524 ( .INP(n2165), .ZN(n2374) );
  NOR2X0 U1525 ( .IN1(n2375), .IN2(n2376), .QN(n2165) );
  AND2X1 U1526 ( .IN1(n2375), .IN2(n2376), .Q(n2164) );
  AO21X1 U1527 ( .IN1(\fpu_add_frac_dp/n2510 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2377), .Q(n2376) );
  MUX21X1 U1528 ( .IN1(n1325), .IN2(n1328), .S(\fpu_add_frac_dp/n2503 ), .Q(
        n2377) );
  AO22X1 U1529 ( .IN1(n2161), .IN2(n2160), .IN3(n2378), .IN4(n244), .Q(n2375)
         );
  OR2X1 U1530 ( .IN1(n2161), .IN2(n2160), .Q(n2378) );
  AO21X1 U1531 ( .IN1(\fpu_add_frac_dp/n2503 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2379), .Q(n2160) );
  MUX21X1 U1532 ( .IN1(n1324), .IN2(n1327), .S(\fpu_add_frac_dp/n2499 ), .Q(
        n2379) );
  AO22X1 U1533 ( .IN1(n2380), .IN2(n2381), .IN3(n2382), .IN4(n245), .Q(n2161)
         );
  NAND2X0 U1534 ( .IN1(n2157), .IN2(n2158), .QN(n2382) );
  INVX0 U1535 ( .INP(n2380), .ZN(n2158) );
  INVX0 U1536 ( .INP(n2381), .ZN(n2157) );
  AO21X1 U1537 ( .IN1(\fpu_add_frac_dp/n2499 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2383), .Q(n2381) );
  MUX21X1 U1538 ( .IN1(n1323), .IN2(n64), .S(\fpu_add_frac_dp/n2507 ), .Q(
        n2383) );
  OA21X1 U1539 ( .IN1(n204), .IN2(n2154), .IN3(n2384), .Q(n2380) );
  INVX0 U1540 ( .INP(n2155), .ZN(n2384) );
  NOR2X0 U1541 ( .IN1(n2385), .IN2(n2386), .QN(n2155) );
  AND2X1 U1542 ( .IN1(n2385), .IN2(n2386), .Q(n2154) );
  AO21X1 U1543 ( .IN1(\fpu_add_frac_dp/n2507 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2387), .Q(n2386) );
  MUX21X1 U1544 ( .IN1(n155), .IN2(n1328), .S(\fpu_add_frac_dp/n2419 ), .Q(
        n2387) );
  AO22X1 U1545 ( .IN1(n2151), .IN2(n2150), .IN3(n2388), .IN4(n246), .Q(n2385)
         );
  OR2X1 U1546 ( .IN1(n2151), .IN2(n2150), .Q(n2388) );
  AO21X1 U1547 ( .IN1(\fpu_add_frac_dp/n2419 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2389), .Q(n2150) );
  MUX21X1 U1548 ( .IN1(n1325), .IN2(n1327), .S(\fpu_add_frac_dp/n2299 ), .Q(
        n2389) );
  AO22X1 U1549 ( .IN1(n2148), .IN2(n2147), .IN3(n2390), .IN4(n247), .Q(n2151)
         );
  OR2X1 U1550 ( .IN1(n2148), .IN2(n2147), .Q(n2390) );
  AO21X1 U1551 ( .IN1(\fpu_add_frac_dp/n2299 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2391), .Q(n2147) );
  MUX21X1 U1552 ( .IN1(n1324), .IN2(n64), .S(\fpu_add_frac_dp/n2420 ), .Q(
        n2391) );
  AO22X1 U1553 ( .IN1(n2145), .IN2(n2144), .IN3(n2392), .IN4(n248), .Q(n2148)
         );
  OR2X1 U1554 ( .IN1(n2145), .IN2(n2144), .Q(n2392) );
  AO21X1 U1555 ( .IN1(\fpu_add_frac_dp/n2420 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2393), .Q(n2144) );
  MUX21X1 U1556 ( .IN1(n1323), .IN2(n1328), .S(\fpu_add_frac_dp/n2273 ), .Q(
        n2393) );
  AO22X1 U1557 ( .IN1(n2142), .IN2(n2394), .IN3(n2395), .IN4(n318), .Q(n2145)
         );
  NAND2X0 U1558 ( .IN1(n2396), .IN2(n2141), .QN(n2395) );
  INVX0 U1559 ( .INP(n2394), .ZN(n2141) );
  AO21X1 U1560 ( .IN1(\fpu_add_frac_dp/n2273 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2397), .Q(n2394) );
  MUX21X1 U1561 ( .IN1(n155), .IN2(n1327), .S(\fpu_add_frac_dp/n2352 ), .Q(
        n2397) );
  INVX0 U1562 ( .INP(n2396), .ZN(n2142) );
  OA22X1 U1563 ( .IN1(n2139), .IN2(n2138), .IN3(n2398), .IN4(
        \fpu_add_frac_dp/n815 ), .Q(n2396) );
  AND2X1 U1564 ( .IN1(n2138), .IN2(n2139), .Q(n2398) );
  AOI21X1 U1565 ( .IN1(\fpu_add_frac_dp/n2352 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2399), .QN(n2138) );
  MUX21X1 U1566 ( .IN1(n1325), .IN2(n64), .S(\fpu_add_frac_dp/n2353 ), .Q(
        n2399) );
  AO21X1 U1567 ( .IN1(\fpu_add_frac_dp/n816 ), .IN2(n2136), .IN3(n2135), .Q(
        n2139) );
  NOR2X0 U1568 ( .IN1(n2400), .IN2(n2401), .QN(n2135) );
  AOI21X1 U1569 ( .IN1(\fpu_add_frac_dp/n817 ), .IN2(n2130), .IN3(n2402), .QN(
        n2401) );
  NAND3X0 U1570 ( .IN1(n2400), .IN2(n2131), .IN3(n2403), .QN(n2136) );
  NAND2X0 U1571 ( .IN1(\fpu_add_frac_dp/n817 ), .IN2(n2130), .QN(n2403) );
  NAND2X0 U1572 ( .IN1(n2404), .IN2(n2405), .QN(n2130) );
  INVX0 U1573 ( .INP(n2402), .ZN(n2131) );
  NOR2X0 U1574 ( .IN1(n2404), .IN2(n2405), .QN(n2402) );
  AO21X1 U1575 ( .IN1(\fpu_add_frac_dp/n2434 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2406), .Q(n2405) );
  MUX21X1 U1576 ( .IN1(n1324), .IN2(n1328), .S(\fpu_add_frac_dp/n2433 ), .Q(
        n2406) );
  AO22X1 U1577 ( .IN1(n2127), .IN2(n2126), .IN3(n2407), .IN4(n249), .Q(n2404)
         );
  OR2X1 U1578 ( .IN1(n2127), .IN2(n2126), .Q(n2407) );
  AO21X1 U1579 ( .IN1(\fpu_add_frac_dp/n2433 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2408), .Q(n2126) );
  MUX21X1 U1580 ( .IN1(n1323), .IN2(n1327), .S(\fpu_add_frac_dp/n2297 ), .Q(
        n2408) );
  AO22X1 U1581 ( .IN1(n2124), .IN2(n2123), .IN3(n2409), .IN4(n250), .Q(n2127)
         );
  OR2X1 U1582 ( .IN1(n2124), .IN2(n2123), .Q(n2409) );
  AO21X1 U1583 ( .IN1(\fpu_add_frac_dp/n2297 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2410), .Q(n2123) );
  MUX21X1 U1584 ( .IN1(n155), .IN2(n64), .S(\fpu_add_frac_dp/n2272 ), .Q(n2410) );
  AO22X1 U1585 ( .IN1(n2121), .IN2(n2120), .IN3(n2411), .IN4(n251), .Q(n2124)
         );
  OR2X1 U1586 ( .IN1(n2120), .IN2(n2121), .Q(n2411) );
  AO21X1 U1587 ( .IN1(\fpu_add_frac_dp/n2272 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2412), .Q(n2120) );
  MUX21X1 U1588 ( .IN1(n1325), .IN2(n1328), .S(\fpu_add_frac_dp/n2298 ), .Q(
        n2412) );
  OA22X1 U1589 ( .IN1(n179), .IN2(n2413), .IN3(n2117), .IN4(n2116), .Q(n2121)
         );
  INVX0 U1590 ( .INP(n2118), .ZN(n2413) );
  NAND2X0 U1591 ( .IN1(n2116), .IN2(n2117), .QN(n2118) );
  AO21X1 U1592 ( .IN1(\fpu_add_frac_dp/n2298 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2414), .Q(n2117) );
  MUX21X1 U1593 ( .IN1(n1324), .IN2(n1327), .S(\fpu_add_frac_dp/n2359 ), .Q(
        n2414) );
  AOI21X1 U1594 ( .IN1(\fpu_add_frac_dp/n822 ), .IN2(n2113), .IN3(n2112), .QN(
        n2116) );
  NOR2X0 U1595 ( .IN1(n2415), .IN2(n2416), .QN(n2112) );
  OA21X1 U1596 ( .IN1(n180), .IN2(n2417), .IN3(n2108), .Q(n2416) );
  NAND3X0 U1597 ( .IN1(n2415), .IN2(n2108), .IN3(n2418), .QN(n2113) );
  NAND2X0 U1598 ( .IN1(\fpu_add_frac_dp/n823 ), .IN2(n2107), .QN(n2418) );
  INVX0 U1599 ( .INP(n2417), .ZN(n2107) );
  NOR2X0 U1600 ( .IN1(n2419), .IN2(n2420), .QN(n2417) );
  NAND2X0 U1601 ( .IN1(n2420), .IN2(n2419), .QN(n2108) );
  NAND2X0 U1602 ( .IN1(n2101), .IN2(n2104), .QN(n2419) );
  NAND2X0 U1603 ( .IN1(\fpu_add_frac_dp/n824 ), .IN2(n2103), .QN(n2104) );
  NAND2X0 U1604 ( .IN1(n2421), .IN2(n2422), .QN(n2103) );
  OR2X1 U1605 ( .IN1(n2422), .IN2(n2421), .Q(n2101) );
  AO21X1 U1606 ( .IN1(\fpu_add_frac_dp/n2362 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2423), .Q(n2421) );
  MUX21X1 U1607 ( .IN1(n1323), .IN2(n64), .S(\fpu_add_frac_dp/n2304 ), .Q(
        n2423) );
  AO22X1 U1608 ( .IN1(n2098), .IN2(n2097), .IN3(n2424), .IN4(n252), .Q(n2422)
         );
  OR2X1 U1609 ( .IN1(n2098), .IN2(n2097), .Q(n2424) );
  AO21X1 U1610 ( .IN1(\fpu_add_frac_dp/n2304 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2425), .Q(n2097) );
  MUX21X1 U1611 ( .IN1(n1327), .IN2(n1325), .S(\fpu_add_frac_dp/n2389 ), .Q(
        n2425) );
  AO22X1 U1612 ( .IN1(n2095), .IN2(n2094), .IN3(n2426), .IN4(n253), .Q(n2098)
         );
  OR2X1 U1613 ( .IN1(n2095), .IN2(n2094), .Q(n2426) );
  AO21X1 U1614 ( .IN1(\fpu_add_frac_dp/n2369 ), .IN2(n904), .IN3(n2427), .Q(
        n2094) );
  MUX21X1 U1615 ( .IN1(n155), .IN2(n1328), .S(\fpu_add_frac_dp/n2277 ), .Q(
        n2427) );
  AO22X1 U1616 ( .IN1(n2092), .IN2(n2091), .IN3(n2428), .IN4(n260), .Q(n2095)
         );
  OR2X1 U1617 ( .IN1(n2092), .IN2(n2091), .Q(n2428) );
  AO21X1 U1618 ( .IN1(\fpu_add_frac_dp/n2277 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2429), .Q(n2091) );
  MUX21X1 U1619 ( .IN1(n1325), .IN2(n1326), .S(\fpu_add_frac_dp/n2531 ), .Q(
        n2429) );
  AO22X1 U1620 ( .IN1(n2089), .IN2(n2088), .IN3(n2430), .IN4(n261), .Q(n2092)
         );
  OR2X1 U1621 ( .IN1(n2089), .IN2(n2088), .Q(n2430) );
  AO21X1 U1622 ( .IN1(\fpu_add_frac_dp/n2531 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2431), .Q(n2088) );
  MUX21X1 U1623 ( .IN1(n1324), .IN2(n1326), .S(\fpu_add_frac_dp/n2530 ), .Q(
        n2431) );
  AO22X1 U1624 ( .IN1(n2086), .IN2(n2085), .IN3(n2432), .IN4(n224), .Q(n2089)
         );
  OR2X1 U1625 ( .IN1(n2085), .IN2(n2086), .Q(n2432) );
  AO21X1 U1626 ( .IN1(\fpu_add_frac_dp/n2530 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2433), .Q(n2085) );
  MUX21X1 U1627 ( .IN1(n1323), .IN2(n1326), .S(\fpu_add_frac_dp/n2529 ), .Q(
        n2433) );
  OA22X1 U1628 ( .IN1(n2082), .IN2(n2083), .IN3(n222), .IN4(n2434), .Q(n2086)
         );
  AND2X1 U1629 ( .IN1(n2083), .IN2(n2082), .Q(n2434) );
  AO22X1 U1630 ( .IN1(n2080), .IN2(n2079), .IN3(n2435), .IN4(n225), .Q(n2083)
         );
  OR2X1 U1631 ( .IN1(n2079), .IN2(n2080), .Q(n2435) );
  AO21X1 U1632 ( .IN1(\fpu_add_frac_dp/n2528 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2436), .Q(n2079) );
  MUX21X1 U1633 ( .IN1(n155), .IN2(n1326), .S(\fpu_add_frac_dp/n2527 ), .Q(
        n2436) );
  OA22X1 U1634 ( .IN1(n2076), .IN2(n2077), .IN3(n223), .IN4(n2437), .Q(n2080)
         );
  AND2X1 U1635 ( .IN1(n2077), .IN2(n2076), .Q(n2437) );
  OAI22X1 U1636 ( .IN1(n2074), .IN2(n2073), .IN3(n2438), .IN4(
        \fpu_add_frac_dp/n833 ), .QN(n2077) );
  AND2X1 U1637 ( .IN1(n2073), .IN2(n2074), .Q(n2438) );
  AOI21X1 U1638 ( .IN1(\fpu_add_frac_dp/n2526 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2439), .QN(n2073) );
  MUX21X1 U1639 ( .IN1(n1325), .IN2(n1326), .S(\fpu_add_frac_dp/n2525 ), .Q(
        n2439) );
  AO22X1 U1640 ( .IN1(n2070), .IN2(n2071), .IN3(\fpu_add_frac_dp/n834 ), .IN4(
        n2440), .Q(n2074) );
  NAND2X0 U1641 ( .IN1(n2441), .IN2(n2442), .QN(n2440) );
  INVX0 U1642 ( .INP(n2441), .ZN(n2071) );
  OA21X1 U1643 ( .IN1(n220), .IN2(n2067), .IN3(n2443), .Q(n2441) );
  INVX0 U1644 ( .INP(n2068), .ZN(n2443) );
  NOR2X0 U1645 ( .IN1(n2444), .IN2(n2445), .QN(n2068) );
  AND2X1 U1646 ( .IN1(n2444), .IN2(n2445), .Q(n2067) );
  AO21X1 U1647 ( .IN1(\fpu_add_frac_dp/n2524 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2446), .Q(n2445) );
  MUX21X1 U1648 ( .IN1(n1324), .IN2(n1326), .S(\fpu_add_frac_dp/n2523 ), .Q(
        n2446) );
  AO22X1 U1649 ( .IN1(n2064), .IN2(n2063), .IN3(n2447), .IN4(n625), .Q(n2444)
         );
  OR2X1 U1650 ( .IN1(n2064), .IN2(n2063), .Q(n2447) );
  AO21X1 U1651 ( .IN1(\fpu_add_frac_dp/n2523 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2448), .Q(n2063) );
  MUX21X1 U1652 ( .IN1(n1323), .IN2(n1326), .S(\fpu_add_frac_dp/n2522 ), .Q(
        n2448) );
  AO22X1 U1653 ( .IN1(n2061), .IN2(n307), .IN3(n2449), .IN4(n926), .Q(n2064)
         );
  OR2X1 U1654 ( .IN1(n2061), .IN2(n307), .Q(n2449) );
  AO21X1 U1655 ( .IN1(\fpu_add_frac_dp/n2522 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2450), .Q(n2061) );
  MUX21X1 U1656 ( .IN1(n155), .IN2(n1326), .S(\fpu_add_frac_dp/n2539 ), .Q(
        n2450) );
  INVX0 U1657 ( .INP(n2442), .ZN(n2070) );
  AO21X1 U1658 ( .IN1(\fpu_add_frac_dp/n2525 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2451), .Q(n2442) );
  MUX21X1 U1659 ( .IN1(n1325), .IN2(n1326), .S(\fpu_add_frac_dp/n2524 ), .Q(
        n2451) );
  AO21X1 U1660 ( .IN1(\fpu_add_frac_dp/n2527 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2452), .Q(n2076) );
  MUX21X1 U1661 ( .IN1(n1324), .IN2(n1326), .S(\fpu_add_frac_dp/n2526 ), .Q(
        n2452) );
  AO21X1 U1662 ( .IN1(\fpu_add_frac_dp/n2529 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2453), .Q(n2082) );
  MUX21X1 U1663 ( .IN1(n1323), .IN2(n1326), .S(\fpu_add_frac_dp/n2528 ), .Q(
        n2453) );
  AOI21X1 U1664 ( .IN1(\fpu_add_frac_dp/n2432 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2454), .QN(n2420) );
  MUX21X1 U1665 ( .IN1(n155), .IN2(n1326), .S(\fpu_add_frac_dp/n2362 ), .Q(
        n2454) );
  AO21X1 U1666 ( .IN1(\fpu_add_frac_dp/n2359 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2455), .Q(n2415) );
  MUX21X1 U1667 ( .IN1(n1325), .IN2(n1326), .S(\fpu_add_frac_dp/n2432 ), .Q(
        n2455) );
  AO21X1 U1668 ( .IN1(\fpu_add_frac_dp/n2353 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2456), .Q(n2400) );
  MUX21X1 U1669 ( .IN1(n1323), .IN2(n1326), .S(\fpu_add_frac_dp/n2434 ), .Q(
        n2456) );
  INVX0 U1670 ( .INP(n2297), .ZN(n2249) );
  AO21X1 U1671 ( .IN1(\fpu_add_frac_dp/n2369 ), .IN2(n62), .IN3(n2457), .Q(
        n2297) );
  MUX21X1 U1672 ( .IN1(n155), .IN2(n1326), .S(\fpu_add_frac_dp/n2357 ), .Q(
        n2457) );
  AOI21X1 U1673 ( .IN1(\fpu_add_frac_dp/n2369 ), .IN2(n153), .IN3(n2458), .QN(
        n2260) );
  MUX21X1 U1674 ( .IN1(n64), .IN2(n1324), .S(\fpu_add_frac_dp/n2390 ), .Q(
        n2458) );
  INVX0 U1675 ( .INP(n2281), .ZN(n2273) );
  AO21X1 U1676 ( .IN1(\fpu_add_frac_dp/n2498 ), .IN2(\fpu_add_frac_dp/n2369 ), 
        .IN3(n2459), .Q(n2281) );
  MUX21X1 U1677 ( .IN1(n1325), .IN2(n1326), .S(\fpu_add_frac_dp/n2502 ), .Q(
        n2459) );
  AO222X1 U1678 ( .IN1(n2460), .IN2(n583), .IN3(n1322), .IN4(n2461), .IN5(
        n1388), .IN6(n154), .Q(\fpu_add_frac_dp/n3666 ) );
  OAI222X1 U1679 ( .IN1(n2462), .IN2(n2463), .IN3(n2464), .IN4(n2465), .IN5(
        n2466), .IN6(n2467), .QN(n2461) );
  INVX0 U1680 ( .INP(n2468), .ZN(n2467) );
  OA221X1 U1681 ( .IN1(n2469), .IN2(n40), .IN3(n2470), .IN4(n2471), .IN5(n2472), .Q(n2466) );
  OA21X1 U1682 ( .IN1(n2473), .IN2(n2474), .IN3(n2475), .Q(n2472) );
  NAND4X0 U1683 ( .IN1(n2476), .IN2(\fpu_add_frac_dp/n2537 ), .IN3(n2477), 
        .IN4(n2478), .QN(n2475) );
  OA21X1 U1684 ( .IN1(\fpu_add_frac_dp/n2361 ), .IN2(n38), .IN3(n2479), .Q(
        n2477) );
  AO21X1 U1685 ( .IN1(\fpu_add_frac_dp/n2342 ), .IN2(n1271), .IN3(n2480), .Q(
        n2474) );
  AO21X1 U1686 ( .IN1(\fpu_add_frac_dp/n2336 ), .IN2(n177), .IN3(n19), .Q(
        n2471) );
  OA21X1 U1687 ( .IN1(\fpu_add_frac_dp/n5609 ), .IN2(n100), .IN3(
        \fpu_add_frac_dp/n5632 ), .Q(n2469) );
  NAND2X0 U1688 ( .IN1(n2481), .IN2(n2482), .QN(n2465) );
  AO221X1 U1689 ( .IN1(n2483), .IN2(n2484), .IN3(n2485), .IN4(n2486), .IN5(
        n2487), .Q(n2482) );
  NOR4X0 U1690 ( .IN1(\fpu_add_frac_dp/n2313 ), .IN2(n2488), .IN3(n2489), 
        .IN4(n2490), .QN(n2487) );
  OA21X1 U1691 ( .IN1(n2491), .IN2(n74), .IN3(n2492), .Q(n2489) );
  OA21X1 U1692 ( .IN1(\fpu_add_frac_dp/n2405 ), .IN2(n447), .IN3(
        \fpu_add_frac_dp/n662 ), .Q(n2491) );
  NOR2X0 U1693 ( .IN1(\fpu_add_frac_dp/n2402 ), .IN2(\fpu_add_frac_dp/n2470 ), 
        .QN(n2488) );
  NAND2X0 U1694 ( .IN1(\fpu_add_frac_dp/n2344 ), .IN2(n43), .QN(n2486) );
  INVX0 U1695 ( .INP(n2493), .ZN(n2485) );
  NAND2X0 U1696 ( .IN1(\fpu_add_frac_dp/n2363 ), .IN2(n101), .QN(n2484) );
  NOR2X0 U1697 ( .IN1(\fpu_add_frac_dp/n2335 ), .IN2(n2494), .QN(n2483) );
  OA221X1 U1698 ( .IN1(n2495), .IN2(n2496), .IN3(n33), .IN4(n2497), .IN5(n2498), .Q(n2464) );
  OA21X1 U1699 ( .IN1(\fpu_add_frac_dp/n2400 ), .IN2(n2499), .IN3(n2500), .Q(
        n2498) );
  AOI21X1 U1700 ( .IN1(n37), .IN2(\fpu_add_frac_dp/n2437 ), .IN3(
        \fpu_add_frac_dp/n2330 ), .QN(n2499) );
  OAI21X1 U1701 ( .IN1(n2501), .IN2(n173), .IN3(n2502), .QN(n2497) );
  OA21X1 U1702 ( .IN1(n2503), .IN2(n90), .IN3(\fpu_add_frac_dp/n2520 ), .Q(
        n2501) );
  OA21X1 U1703 ( .IN1(\fpu_add_frac_dp/n5642 ), .IN2(n282), .IN3(
        \fpu_add_frac_dp/n670 ), .Q(n2503) );
  OA21X1 U1704 ( .IN1(\fpu_add_frac_dp/n666 ), .IN2(n34), .IN3(
        \fpu_add_frac_dp/n5610 ), .Q(n2495) );
  OA221X1 U1705 ( .IN1(n2504), .IN2(n87), .IN3(n2505), .IN4(n2506), .IN5(n2507), .Q(n2463) );
  OA21X1 U1706 ( .IN1(n2508), .IN2(n2509), .IN3(n2510), .Q(n2507) );
  NAND4X0 U1707 ( .IN1(n2511), .IN2(\fpu_add_frac_dp/n2394 ), .IN3(n2512), 
        .IN4(n2513), .QN(n2510) );
  NAND2X0 U1708 ( .IN1(\fpu_add_frac_dp/n2343 ), .IN2(\fpu_add_frac_dp/n654 ), 
        .QN(n2512) );
  NOR2X0 U1709 ( .IN1(\fpu_add_frac_dp/n2386 ), .IN2(n22), .QN(n2508) );
  OA21X1 U1710 ( .IN1(\fpu_add_frac_dp/n2416 ), .IN2(n92), .IN3(
        \fpu_add_frac_dp/n2290 ), .Q(n2505) );
  OA21X1 U1711 ( .IN1(n94), .IN2(n654), .IN3(\fpu_add_frac_dp/n5618 ), .Q(
        n2504) );
  AO222X1 U1712 ( .IN1(n2460), .IN2(n72), .IN3(n1321), .IN4(n2514), .IN5(n1388), .IN6(n582), .Q(\fpu_add_frac_dp/n3665 ) );
  AO221X1 U1713 ( .IN1(n2515), .IN2(n2516), .IN3(n2468), .IN4(n2517), .IN5(
        n2518), .Q(n2514) );
  NAND2X0 U1714 ( .IN1(n2519), .IN2(n2520), .QN(n2518) );
  NAND4X0 U1715 ( .IN1(n2521), .IN2(\fpu_add_frac_dp/n2363 ), .IN3(n2522), 
        .IN4(n839), .QN(n2520) );
  NAND2X0 U1716 ( .IN1(n2494), .IN2(n2523), .QN(n2522) );
  NAND3X0 U1717 ( .IN1(n346), .IN2(n710), .IN3(n2524), .QN(n2523) );
  NAND2X0 U1718 ( .IN1(n2492), .IN2(n2525), .QN(n2524) );
  NAND3X0 U1719 ( .IN1(\fpu_add_frac_dp/n2409 ), .IN2(n2526), .IN3(
        \fpu_add_frac_dp/n662 ), .QN(n2525) );
  NAND3X0 U1720 ( .IN1(n447), .IN2(n1087), .IN3(n2527), .QN(n2526) );
  NAND2X0 U1721 ( .IN1(\fpu_add_frac_dp/n2344 ), .IN2(\fpu_add_frac_dp/n2411 ), 
        .QN(n2527) );
  AO21X1 U1722 ( .IN1(n2528), .IN2(n2529), .IN3(n2462), .Q(n2519) );
  NAND3X0 U1723 ( .IN1(n2530), .IN2(n2531), .IN3(\fpu_add_frac_dp/n2290 ), 
        .QN(n2529) );
  NAND3X0 U1724 ( .IN1(\fpu_add_frac_dp/n2345 ), .IN2(n2532), .IN3(
        \fpu_add_frac_dp/n2416 ), .QN(n2531) );
  NAND2X0 U1725 ( .IN1(\fpu_add_frac_dp/n5631 ), .IN2(\fpu_add_frac_dp/n2378 ), 
        .QN(n2532) );
  NAND3X0 U1726 ( .IN1(\fpu_add_frac_dp/n2440 ), .IN2(n2533), .IN3(
        \fpu_add_frac_dp/n5618 ), .QN(n2528) );
  NAND3X0 U1727 ( .IN1(n2534), .IN2(n654), .IN3(\fpu_add_frac_dp/n2288 ), .QN(
        n2533) );
  OR3X1 U1728 ( .IN1(n82), .IN2(n2535), .IN3(n171), .Q(n2534) );
  AO222X1 U1729 ( .IN1(n2476), .IN2(n2536), .IN3(n2537), .IN4(n2538), .IN5(
        n2539), .IN6(n2540), .Q(n2517) );
  INVX0 U1730 ( .INP(n2470), .ZN(n2538) );
  NAND3X0 U1731 ( .IN1(n2541), .IN2(n2542), .IN3(n2476), .QN(n2470) );
  NAND3X0 U1732 ( .IN1(\fpu_add_frac_dp/n2336 ), .IN2(n716), .IN3(
        \fpu_add_frac_dp/n659 ), .QN(n2542) );
  NOR2X0 U1733 ( .IN1(n86), .IN2(n19), .QN(n2537) );
  NAND2X0 U1734 ( .IN1(n2478), .IN2(n2543), .QN(n2536) );
  NAND3X0 U1735 ( .IN1(\fpu_add_frac_dp/n2481 ), .IN2(n2479), .IN3(
        \fpu_add_frac_dp/n2537 ), .QN(n2543) );
  INVX0 U1736 ( .INP(n2544), .ZN(n2478) );
  NAND3X0 U1737 ( .IN1(n2545), .IN2(n2546), .IN3(n2547), .QN(n2516) );
  NAND3X0 U1738 ( .IN1(n2548), .IN2(n2549), .IN3(\fpu_add_frac_dp/n5610 ), 
        .QN(n2547) );
  NAND3X0 U1739 ( .IN1(\fpu_add_frac_dp/n2494 ), .IN2(n2550), .IN3(
        \fpu_add_frac_dp/n666 ), .QN(n2549) );
  OR3X1 U1740 ( .IN1(n33), .IN2(n2551), .IN3(n173), .Q(n2550) );
  INVX0 U1741 ( .INP(n2496), .ZN(n2548) );
  OR3X1 U1742 ( .IN1(\fpu_add_frac_dp/n2330 ), .IN2(\fpu_add_frac_dp/n2400 ), 
        .IN3(n2552), .Q(n2545) );
  AO222X1 U1743 ( .IN1(n2460), .IN2(n159), .IN3(n1319), .IN4(n2553), .IN5(
        n1388), .IN6(n63), .Q(\fpu_add_frac_dp/n3664 ) );
  NAND2X0 U1744 ( .IN1(n2554), .IN2(n2555), .QN(n2553) );
  NAND3X0 U1745 ( .IN1(n2556), .IN2(n2557), .IN3(n2515), .QN(n2555) );
  NAND2X0 U1746 ( .IN1(n2502), .IN2(n2558), .QN(n2557) );
  NAND3X0 U1747 ( .IN1(\fpu_add_frac_dp/n2513 ), .IN2(n2551), .IN3(
        \fpu_add_frac_dp/n668 ), .QN(n2558) );
  MUX21X1 U1748 ( .IN1(n2559), .IN2(n2560), .S(n2481), .Q(n2554) );
  NAND2X0 U1749 ( .IN1(n2561), .IN2(n2562), .QN(n2560) );
  AO21X1 U1750 ( .IN1(n2563), .IN2(n2564), .IN3(n2565), .Q(n2562) );
  OA22X1 U1751 ( .IN1(n2566), .IN2(n2567), .IN3(n2568), .IN4(n2569), .Q(n2559)
         );
  NOR4X0 U1752 ( .IN1(n2570), .IN2(n22), .IN3(n175), .IN4(n104), .QN(n2566) );
  AO221X1 U1753 ( .IN1(n2571), .IN2(n2476), .IN3(n2539), .IN4(n716), .IN5(n85), 
        .Q(n2570) );
  INVX0 U1754 ( .INP(n2473), .ZN(n2539) );
  NOR2X0 U1755 ( .IN1(n2541), .IN2(n2544), .QN(n2571) );
  AO222X1 U1756 ( .IN1(n2460), .IN2(n178), .IN3(n1322), .IN4(n2572), .IN5(
        n1388), .IN6(n584), .Q(\fpu_add_frac_dp/n3663 ) );
  NAND4X0 U1757 ( .IN1(n2573), .IN2(n2574), .IN3(n2575), .IN4(n2576), .QN(
        n2572) );
  NAND3X0 U1758 ( .IN1(n2561), .IN2(n2492), .IN3(n2521), .QN(n2576) );
  NOR2X0 U1759 ( .IN1(n2577), .IN2(n2500), .QN(n2521) );
  NAND3X0 U1760 ( .IN1(n2476), .IN2(n2541), .IN3(n2468), .QN(n2575) );
  NAND3X0 U1761 ( .IN1(n2568), .IN2(n2578), .IN3(n2511), .QN(n2574) );
  INVX0 U1762 ( .INP(n2569), .ZN(n2511) );
  INVX0 U1763 ( .INP(n2513), .ZN(n2568) );
  NAND2X0 U1764 ( .IN1(n2515), .IN2(n2502), .QN(n2573) );
  AO222X1 U1765 ( .IN1(n2460), .IN2(n67), .IN3(n1321), .IN4(n2579), .IN5(n1388), .IN6(n762), .Q(\fpu_add_frac_dp/n3662 ) );
  NAND3X0 U1766 ( .IN1(n2580), .IN2(n2581), .IN3(n2582), .QN(
        \fpu_add_frac_dp/n3661 ) );
  OR2X1 U1767 ( .IN1(n2046), .IN2(\fpu_add_frac_dp/n593 ), .Q(n2582) );
  AO222X1 U1768 ( .IN1(n2583), .IN2(n67), .IN3(n2584), .IN4(n2579), .IN5(n1388), .IN6(n2), .Q(\fpu_add_frac_dp/n3660 ) );
  AO222X1 U1769 ( .IN1(\fpu_add_exp_dp/n432 ), .IN2(n2583), .IN3(n2585), .IN4(
        n2584), .IN5(n1379), .IN6(n2586), .Q(\fpu_add_frac_dp/n3659 ) );
  INVX0 U1770 ( .INP(n2580), .ZN(n2584) );
  NAND2X0 U1771 ( .IN1(n1320), .IN2(n2481), .QN(n2580) );
  INVX0 U1772 ( .INP(n2577), .ZN(n2481) );
  INVX0 U1773 ( .INP(n2581), .ZN(n2583) );
  NAND2X0 U1774 ( .IN1(n2460), .IN2(n69), .QN(n2581) );
  OAI22X1 U1775 ( .IN1(n2046), .IN2(\fpu_add_frac_dp/n5633 ), .IN3(n1745), 
        .IN4(n2587), .QN(\fpu_add_frac_dp/n3658 ) );
  OAI22X1 U1776 ( .IN1(n2046), .IN2(\fpu_add_frac_dp/n589 ), .IN3(n1745), 
        .IN4(n2587), .QN(\fpu_add_frac_dp/n3657 ) );
  MUX21X1 U1777 ( .IN1(n2588), .IN2(n2589), .S(n2590), .Q(n2587) );
  NAND2X0 U1778 ( .IN1(\fpu_add_exp_dp/n433 ), .IN2(n67), .QN(n2589) );
  NAND2X0 U1779 ( .IN1(n2579), .IN2(n2577), .QN(n2588) );
  INVX0 U1780 ( .INP(n2585), .ZN(n2579) );
  AO21X1 U1781 ( .IN1(n1397), .IN2(n2591), .IN3(n2592), .Q(
        \fpu_add_frac_dp/n3656 ) );
  AO21X1 U1782 ( .IN1(n1396), .IN2(n596), .IN3(n2592), .Q(
        \fpu_add_frac_dp/n3655 ) );
  AO21X1 U1783 ( .IN1(n1397), .IN2(n1144), .IN3(n2592), .Q(
        \fpu_add_frac_dp/n3654 ) );
  NAND2X0 U1784 ( .IN1(n2593), .IN2(n2594), .QN(n2592) );
  NAND3X0 U1785 ( .IN1(n1320), .IN2(n2577), .IN3(n2585), .QN(n2594) );
  NOR2X0 U1786 ( .IN1(n2468), .IN2(n2515), .QN(n2585) );
  NOR2X0 U1787 ( .IN1(n2564), .IN2(n2577), .QN(n2515) );
  INVX0 U1788 ( .INP(n2500), .ZN(n2564) );
  NOR2X0 U1789 ( .IN1(n2493), .IN2(n2595), .QN(n2500) );
  NOR2X0 U1790 ( .IN1(n2578), .IN2(n2596), .QN(n2468) );
  NAND3X0 U1791 ( .IN1(\fpu_add_exp_dp/n432 ), .IN2(n2460), .IN3(
        \fpu_add_exp_dp/n433 ), .QN(n2593) );
  AO21X1 U1792 ( .IN1(n1396), .IN2(n641), .IN3(n2597), .Q(
        \fpu_add_frac_dp/n3653 ) );
  AO21X1 U1793 ( .IN1(n1397), .IN2(n166), .IN3(n2597), .Q(
        \fpu_add_frac_dp/n3652 ) );
  AO21X1 U1794 ( .IN1(n1396), .IN2(n1145), .IN3(n2598), .Q(
        \fpu_add_frac_dp/n3651 ) );
  AO21X1 U1795 ( .IN1(n1397), .IN2(n311), .IN3(n2598), .Q(
        \fpu_add_frac_dp/n3650 ) );
  AO21X1 U1796 ( .IN1(n1397), .IN2(n653), .IN3(n2599), .Q(
        \fpu_add_frac_dp/n3649 ) );
  AO21X1 U1797 ( .IN1(n1404), .IN2(n746), .IN3(n2599), .Q(
        \fpu_add_frac_dp/n3648 ) );
  AO22X1 U1798 ( .IN1(n1421), .IN2(n296), .IN3(n1442), .IN4(n2600), .Q(
        \fpu_add_frac_dp/n3647 ) );
  NAND2X0 U1799 ( .IN1(n2601), .IN2(n2602), .QN(n2600) );
  AO21X1 U1800 ( .IN1(n1404), .IN2(n962), .IN3(n2597), .Q(
        \fpu_add_frac_dp/n3646 ) );
  AND2X1 U1801 ( .IN1(n1442), .IN2(n2603), .Q(n2597) );
  AO221X1 U1802 ( .IN1(n2604), .IN2(n2605), .IN3(n2606), .IN4(n2058), .IN5(
        n2607), .Q(n2603) );
  AO21X1 U1803 ( .IN1(n2608), .IN2(n2609), .IN3(n2610), .Q(n2607) );
  AO21X1 U1804 ( .IN1(n2057), .IN2(n2608), .IN3(a1stg_fsdtoix), .Q(n2606) );
  NAND2X0 U1805 ( .IN1(n2052), .IN2(n2051), .QN(n2605) );
  NAND2X0 U1806 ( .IN1(n2611), .IN2(n2612), .QN(n2051) );
  AO21X1 U1807 ( .IN1(n1404), .IN2(n255), .IN3(n2598), .Q(
        \fpu_add_frac_dp/n3645 ) );
  AND2X1 U1808 ( .IN1(n1442), .IN2(n2613), .Q(n2598) );
  AO221X1 U1809 ( .IN1(a1stg_fsdtoix), .IN2(n2614), .IN3(n2604), .IN4(n2615), 
        .IN5(n2616), .Q(n2613) );
  AO21X1 U1810 ( .IN1(n2608), .IN2(n2617), .IN3(n2610), .Q(n2616) );
  XOR3X1 U1811 ( .IN1(n2618), .IN2(n2619), .IN3(n2609), .Q(n2617) );
  XOR3X1 U1812 ( .IN1(n2620), .IN2(n2621), .IN3(n2052), .Q(n2615) );
  AO21X1 U1813 ( .IN1(n2619), .IN2(n2622), .IN3(n2623), .Q(n2614) );
  AO21X1 U1814 ( .IN1(n1404), .IN2(n755), .IN3(n2599), .Q(
        \fpu_add_frac_dp/n3644 ) );
  AND2X1 U1815 ( .IN1(n1442), .IN2(n2624), .Q(n2599) );
  AO221X1 U1816 ( .IN1(n2625), .IN2(n2604), .IN3(n2608), .IN4(n2626), .IN5(
        n2627), .Q(n2624) );
  AO21X1 U1817 ( .IN1(a1stg_fsdtoix), .IN2(n2628), .IN3(n2610), .Q(n2627) );
  INVX0 U1818 ( .INP(n2629), .ZN(n2628) );
  XOR3X1 U1819 ( .IN1(n2630), .IN2(n2631), .IN3(n2632), .Q(n2626) );
  XOR3X1 U1820 ( .IN1(n2633), .IN2(n2634), .IN3(n2635), .Q(n2625) );
  AO21X1 U1821 ( .IN1(n1404), .IN2(n693), .IN3(n2636), .Q(
        \fpu_add_frac_dp/n3643 ) );
  AO21X1 U1822 ( .IN1(\fpu_add_frac_dp/n2306 ), .IN2(n1415), .IN3(n2637), .Q(
        \fpu_add_frac_dp/n3642 ) );
  AO21X1 U1823 ( .IN1(n1404), .IN2(n2638), .IN3(n2639), .Q(
        \fpu_add_frac_dp/n3641 ) );
  AO21X1 U1824 ( .IN1(n1405), .IN2(n1063), .IN3(n2636), .Q(
        \fpu_add_frac_dp/n3640 ) );
  AO21X1 U1825 ( .IN1(\fpu_add_frac_dp/n2399 ), .IN2(n1415), .IN3(n2636), .Q(
        \fpu_add_frac_dp/n3639 ) );
  AO21X1 U1826 ( .IN1(n1405), .IN2(n581), .IN3(n2636), .Q(
        \fpu_add_frac_dp/n3638 ) );
  AO21X1 U1827 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n1416), .IN3(n2636), .Q(
        \fpu_add_frac_dp/n3637 ) );
  AO21X1 U1828 ( .IN1(\fpu_add_frac_dp/n2322 ), .IN2(n1415), .IN3(n2636), .Q(
        \fpu_add_frac_dp/n3636 ) );
  AND2X1 U1829 ( .IN1(n1443), .IN2(n2640), .Q(n2636) );
  AO221X1 U1830 ( .IN1(a1stg_fsdtoix), .IN2(n2641), .IN3(n2608), .IN4(n2642), 
        .IN5(n2643), .Q(n2640) );
  AO21X1 U1831 ( .IN1(n2644), .IN2(n2604), .IN3(n2610), .Q(n2643) );
  XNOR3X1 U1832 ( .IN1(n2645), .IN2(n2646), .IN3(n2647), .Q(n2644) );
  XOR3X1 U1833 ( .IN1(n2648), .IN2(n2649), .IN3(n2650), .Q(n2642) );
  OR2X1 U1834 ( .IN1(n2651), .IN2(n2652), .Q(n2641) );
  AO21X1 U1835 ( .IN1(n1405), .IN2(n1220), .IN3(n2637), .Q(
        \fpu_add_frac_dp/n3635 ) );
  AO21X1 U1836 ( .IN1(n1405), .IN2(n1221), .IN3(n2637), .Q(
        \fpu_add_frac_dp/n3634 ) );
  AO21X1 U1837 ( .IN1(n1405), .IN2(n1126), .IN3(n2637), .Q(
        \fpu_add_frac_dp/n3633 ) );
  AO21X1 U1838 ( .IN1(n1405), .IN2(n2653), .IN3(n2637), .Q(
        \fpu_add_frac_dp/n3632 ) );
  AO21X1 U1839 ( .IN1(\fpu_add_frac_dp/n2382 ), .IN2(n1416), .IN3(n2637), .Q(
        \fpu_add_frac_dp/n3631 ) );
  AND2X1 U1840 ( .IN1(n1442), .IN2(n2654), .Q(n2637) );
  AO221X1 U1841 ( .IN1(a1stg_fsdtoix), .IN2(n2655), .IN3(n2608), .IN4(n2656), 
        .IN5(n2657), .Q(n2654) );
  AO21X1 U1842 ( .IN1(n2658), .IN2(n2604), .IN3(n2610), .Q(n2657) );
  XNOR3X1 U1843 ( .IN1(n2659), .IN2(n2660), .IN3(n2661), .Q(n2658) );
  XOR3X1 U1844 ( .IN1(n2662), .IN2(n2663), .IN3(n2664), .Q(n2656) );
  OR2X1 U1845 ( .IN1(n2665), .IN2(n2666), .Q(n2655) );
  AO21X1 U1846 ( .IN1(n1405), .IN2(n47), .IN3(n2639), .Q(
        \fpu_add_frac_dp/n3630 ) );
  AO21X1 U1847 ( .IN1(n1405), .IN2(n5), .IN3(n2639), .Q(
        \fpu_add_frac_dp/n3629 ) );
  AO21X1 U1848 ( .IN1(n1405), .IN2(n1222), .IN3(n2639), .Q(
        \fpu_add_frac_dp/n3628 ) );
  AND2X1 U1849 ( .IN1(n1442), .IN2(n2667), .Q(n2639) );
  AO21X1 U1850 ( .IN1(n1405), .IN2(n1124), .IN3(n1930), .Q(
        \fpu_add_frac_dp/n3627 ) );
  AO21X1 U1851 ( .IN1(n1405), .IN2(n118), .IN3(n1930), .Q(
        \fpu_add_frac_dp/n3626 ) );
  AO21X1 U1852 ( .IN1(n1406), .IN2(n20), .IN3(n1930), .Q(
        \fpu_add_frac_dp/n3625 ) );
  NOR2X0 U1853 ( .IN1(n2667), .IN2(n1745), .QN(n1930) );
  AO221X1 U1854 ( .IN1(n2668), .IN2(n2669), .IN3(n2608), .IN4(n2670), .IN5(
        n2671), .Q(n2667) );
  AO21X1 U1855 ( .IN1(n2672), .IN2(n2604), .IN3(n2610), .Q(n2671) );
  AO22X1 U1856 ( .IN1(n2608), .IN2(n2059), .IN3(n2604), .IN4(n2054), .Q(n2610)
         );
  NAND4X0 U1857 ( .IN1(n2673), .IN2(n2674), .IN3(n2675), .IN4(n2676), .QN(
        n2054) );
  NOR2X0 U1858 ( .IN1(n2677), .IN2(n2678), .QN(n2676) );
  XNOR3X1 U1859 ( .IN1(n2679), .IN2(n2680), .IN3(n2681), .Q(n2678) );
  XNOR3X1 U1860 ( .IN1(n2682), .IN2(n2683), .IN3(n2684), .Q(n2677) );
  NAND3X0 U1861 ( .IN1(n2685), .IN2(n2686), .IN3(n2687), .QN(n2675) );
  XOR3X1 U1862 ( .IN1(n2688), .IN2(n2689), .IN3(n2690), .Q(n2674) );
  XOR3X1 U1863 ( .IN1(n2691), .IN2(n2692), .IN3(n2693), .Q(n2673) );
  NAND4X0 U1864 ( .IN1(n2694), .IN2(n2695), .IN3(n2696), .IN4(n2697), .QN(
        n2059) );
  NOR2X0 U1865 ( .IN1(n2698), .IN2(n2699), .QN(n2697) );
  XOR3X1 U1866 ( .IN1(n2700), .IN2(n2701), .IN3(n2702), .Q(n2699) );
  OA22X1 U1867 ( .IN1(\fpu_add_exp_dp/n205 ), .IN2(\fpu_add_exp_dp/n235 ), 
        .IN3(\fpu_add_exp_dp/n189 ), .IN4(\fpu_add_exp_dp/n238 ), .Q(n2701) );
  XOR3X1 U1868 ( .IN1(n2703), .IN2(n2704), .IN3(n2705), .Q(n2698) );
  OA22X1 U1869 ( .IN1(\fpu_add_exp_dp/n204 ), .IN2(\fpu_add_exp_dp/n234 ), 
        .IN3(\fpu_add_exp_dp/n188 ), .IN4(\fpu_add_exp_dp/n237 ), .Q(n2704) );
  XOR3X1 U1870 ( .IN1(n2706), .IN2(n2707), .IN3(n2708), .Q(n2696) );
  NAND2X0 U1871 ( .IN1(n2709), .IN2(n2710), .QN(n2708) );
  NOR2X0 U1872 ( .IN1(\fpu_add_exp_dp/n234 ), .IN2(\fpu_add_exp_dp/n185 ), 
        .QN(n2707) );
  XOR3X1 U1873 ( .IN1(n2710), .IN2(n2711), .IN3(n2709), .Q(n2695) );
  NOR2X0 U1874 ( .IN1(n2712), .IN2(n2713), .QN(n2709) );
  NOR2X0 U1875 ( .IN1(\fpu_add_exp_dp/n186 ), .IN2(\fpu_add_exp_dp/n235 ), 
        .QN(n2711) );
  XOR3X1 U1876 ( .IN1(n2713), .IN2(n2714), .IN3(n2712), .Q(n2694) );
  NAND2X0 U1877 ( .IN1(n2703), .IN2(n2705), .QN(n2712) );
  NOR2X0 U1878 ( .IN1(n2702), .IN2(n2700), .QN(n2705) );
  AO22X1 U1879 ( .IN1(n2715), .IN2(n2716), .IN3(n2717), .IN4(n2718), .Q(n2702)
         );
  OR2X1 U1880 ( .IN1(n2716), .IN2(n2715), .Q(n2717) );
  NOR2X0 U1881 ( .IN1(\fpu_add_exp_dp/n236 ), .IN2(\fpu_add_exp_dp/n187 ), 
        .QN(n2714) );
  AND2X1 U1882 ( .IN1(n2050), .IN2(n2719), .Q(n2604) );
  XNOR3X1 U1883 ( .IN1(n2720), .IN2(n2721), .IN3(n2722), .Q(n2672) );
  XOR3X1 U1884 ( .IN1(n2718), .IN2(n2715), .IN3(n2716), .Q(n2670) );
  AO22X1 U1885 ( .IN1(n2663), .IN2(n2664), .IN3(n2723), .IN4(n2662), .Q(n2716)
         );
  OR2X1 U1886 ( .IN1(n2664), .IN2(n2663), .Q(n2723) );
  AO22X1 U1887 ( .IN1(n2648), .IN2(n2650), .IN3(n2724), .IN4(n2649), .Q(n2664)
         );
  OR2X1 U1888 ( .IN1(n2650), .IN2(n2648), .Q(n2724) );
  AO22X1 U1889 ( .IN1(n2630), .IN2(n2632), .IN3(n2725), .IN4(n2631), .Q(n2650)
         );
  OR2X1 U1890 ( .IN1(n2632), .IN2(n2630), .Q(n2725) );
  AO22X1 U1891 ( .IN1(n2618), .IN2(n2726), .IN3(n2727), .IN4(n2728), .Q(n2632)
         );
  INVX0 U1892 ( .INP(n2619), .ZN(n2728) );
  OR2X1 U1893 ( .IN1(n2726), .IN2(n2618), .Q(n2727) );
  INVX0 U1894 ( .INP(n2609), .ZN(n2726) );
  NOR2X0 U1895 ( .IN1(n2058), .IN2(n2057), .QN(n2609) );
  OA22X1 U1896 ( .IN1(\fpu_add_exp_dp/n211 ), .IN2(\fpu_add_exp_dp/n241 ), 
        .IN3(\fpu_add_exp_dp/n195 ), .IN4(\fpu_add_exp_dp/n244 ), .Q(n2057) );
  INVX0 U1897 ( .INP(n2622), .ZN(n2058) );
  OA22X1 U1898 ( .IN1(\fpu_add_exp_dp/n243 ), .IN2(\fpu_add_exp_dp/n194 ), 
        .IN3(\fpu_add_exp_dp/n240 ), .IN4(\fpu_add_exp_dp/n210 ), .Q(n2618) );
  OA22X1 U1899 ( .IN1(\fpu_add_exp_dp/n242 ), .IN2(\fpu_add_exp_dp/n193 ), 
        .IN3(\fpu_add_exp_dp/n239 ), .IN4(\fpu_add_exp_dp/n209 ), .Q(n2630) );
  OA22X1 U1900 ( .IN1(\fpu_add_exp_dp/n241 ), .IN2(\fpu_add_exp_dp/n192 ), 
        .IN3(\fpu_add_exp_dp/n238 ), .IN4(\fpu_add_exp_dp/n208 ), .Q(n2648) );
  OA22X1 U1901 ( .IN1(\fpu_add_exp_dp/n240 ), .IN2(\fpu_add_exp_dp/n191 ), 
        .IN3(\fpu_add_exp_dp/n237 ), .IN4(\fpu_add_exp_dp/n207 ), .Q(n2663) );
  OA22X1 U1902 ( .IN1(\fpu_add_exp_dp/n239 ), .IN2(\fpu_add_exp_dp/n190 ), 
        .IN3(\fpu_add_exp_dp/n236 ), .IN4(\fpu_add_exp_dp/n206 ), .Q(n2715) );
  NOR2X0 U1903 ( .IN1(n1867), .IN2(n2050), .QN(n2608) );
  OR2X1 U1904 ( .IN1(n2729), .IN2(n2730), .Q(n2669) );
  AO222X1 U1905 ( .IN1(n1322), .IN2(n652), .IN3(n2460), .IN4(n103), .IN5(n1388), .IN6(n219), .Q(\fpu_add_frac_dp/n3624 ) );
  AO222X1 U1906 ( .IN1(n1321), .IN2(n103), .IN3(n2460), .IN4(n282), .IN5(n1388), .IN6(n48), .Q(\fpu_add_frac_dp/n3623 ) );
  AO222X1 U1907 ( .IN1(n1319), .IN2(n282), .IN3(n2460), .IN4(n671), .IN5(n1388), .IN6(n115), .Q(\fpu_add_frac_dp/n3622 ) );
  AO222X1 U1908 ( .IN1(n1320), .IN2(n671), .IN3(n2460), .IN4(n90), .IN5(n1388), 
        .IN6(n50), .Q(\fpu_add_frac_dp/n3621 ) );
  AO222X1 U1909 ( .IN1(n1322), .IN2(n90), .IN3(n2460), .IN4(n626), .IN5(n1388), 
        .IN6(n284), .Q(\fpu_add_frac_dp/n3620 ) );
  AO222X1 U1910 ( .IN1(n1321), .IN2(n626), .IN3(n2460), .IN4(n173), .IN5(n1388), .IN6(n51), .Q(\fpu_add_frac_dp/n3619 ) );
  AO222X1 U1911 ( .IN1(n1319), .IN2(n173), .IN3(n2460), .IN4(n33), .IN5(n1387), 
        .IN6(n124), .Q(\fpu_add_frac_dp/n3618 ) );
  AO222X1 U1912 ( .IN1(n1320), .IN2(n33), .IN3(n2460), .IN4(n623), .IN5(n1387), 
        .IN6(n286), .Q(\fpu_add_frac_dp/n3617 ) );
  AO222X1 U1913 ( .IN1(n1322), .IN2(n623), .IN3(n2460), .IN4(n34), .IN5(n1387), 
        .IN6(n123), .Q(\fpu_add_frac_dp/n3616 ) );
  AO222X1 U1914 ( .IN1(n1321), .IN2(n34), .IN3(n2460), .IN4(n12), .IN5(n1387), 
        .IN6(n285), .Q(\fpu_add_frac_dp/n3615 ) );
  AO222X1 U1915 ( .IN1(n1319), .IN2(n12), .IN3(n2460), .IN4(n691), .IN5(n1387), 
        .IN6(n119), .Q(\fpu_add_frac_dp/n3614 ) );
  AO222X1 U1916 ( .IN1(n1320), .IN2(n691), .IN3(n2460), .IN4(n37), .IN5(n1387), 
        .IN6(n264), .Q(\fpu_add_frac_dp/n3613 ) );
  AO222X1 U1917 ( .IN1(n1322), .IN2(n37), .IN3(n2460), .IN4(n597), .IN5(n1387), 
        .IN6(n107), .Q(\fpu_add_frac_dp/n3612 ) );
  AO222X1 U1918 ( .IN1(n1321), .IN2(n597), .IN3(n2460), .IN4(
        \fpu_add_frac_dp/n2330 ), .IN5(n1387), .IN6(n257), .Q(
        \fpu_add_frac_dp/n3611 ) );
  AO222X1 U1919 ( .IN1(n1319), .IN2(\fpu_add_frac_dp/n2330 ), .IN3(n2460), 
        .IN4(\fpu_add_frac_dp/n2400 ), .IN5(n1387), .IN6(n45), .Q(
        \fpu_add_frac_dp/n3610 ) );
  AO222X1 U1920 ( .IN1(n1320), .IN2(\fpu_add_frac_dp/n2400 ), .IN3(n2460), 
        .IN4(n328), .IN5(n1387), .IN6(n130), .Q(\fpu_add_frac_dp/n3609 ) );
  AO222X1 U1921 ( .IN1(n1322), .IN2(n328), .IN3(n2460), .IN4(n43), .IN5(n1387), 
        .IN6(n756), .Q(\fpu_add_frac_dp/n3608 ) );
  AO222X1 U1922 ( .IN1(n1321), .IN2(n43), .IN3(n2460), .IN4(n111), .IN5(n1387), 
        .IN6(n430), .Q(\fpu_add_frac_dp/n3607 ) );
  AO222X1 U1923 ( .IN1(n1319), .IN2(n111), .IN3(n2460), .IN4(n664), .IN5(n1386), .IN6(n429), .Q(\fpu_add_frac_dp/n3606 ) );
  AO222X1 U1924 ( .IN1(n1320), .IN2(n664), .IN3(n2460), .IN4(
        \fpu_add_frac_dp/n2339 ), .IN5(n1386), .IN6(n431), .Q(
        \fpu_add_frac_dp/n3605 ) );
  AO222X1 U1925 ( .IN1(n1322), .IN2(\fpu_add_frac_dp/n2339 ), .IN3(n2460), 
        .IN4(\fpu_add_frac_dp/n2405 ), .IN5(n1386), .IN6(n432), .Q(
        \fpu_add_frac_dp/n3604 ) );
  AO222X1 U1926 ( .IN1(n1321), .IN2(\fpu_add_frac_dp/n2405 ), .IN3(n2460), 
        .IN4(n594), .IN5(n1386), .IN6(n450), .Q(\fpu_add_frac_dp/n3603 ) );
  AO222X1 U1927 ( .IN1(n1319), .IN2(n594), .IN3(n2460), .IN4(n74), .IN5(n1386), 
        .IN6(n449), .Q(\fpu_add_frac_dp/n3602 ) );
  AO222X1 U1928 ( .IN1(n1320), .IN2(n74), .IN3(n2460), .IN4(n331), .IN5(n1386), 
        .IN6(n750), .Q(\fpu_add_frac_dp/n3601 ) );
  AO222X1 U1929 ( .IN1(n1322), .IN2(n331), .IN3(n2460), .IN4(n116), .IN5(n1386), .IN6(n752), .Q(\fpu_add_frac_dp/n3600 ) );
  AO222X1 U1930 ( .IN1(n1321), .IN2(n116), .IN3(n2460), .IN4(
        \fpu_add_frac_dp/n2402 ), .IN5(n1386), .IN6(n748), .Q(
        \fpu_add_frac_dp/n3599 ) );
  AO222X1 U1931 ( .IN1(n1319), .IN2(\fpu_add_frac_dp/n2402 ), .IN3(n2460), 
        .IN4(\fpu_add_frac_dp/n2313 ), .IN5(n1386), .IN6(n448), .Q(
        \fpu_add_frac_dp/n3598 ) );
  AO222X1 U1932 ( .IN1(n1320), .IN2(\fpu_add_frac_dp/n2313 ), .IN3(n2460), 
        .IN4(n329), .IN5(n1386), .IN6(n749), .Q(\fpu_add_frac_dp/n3597 ) );
  AO222X1 U1933 ( .IN1(n1322), .IN2(n329), .IN3(n2460), .IN4(n101), .IN5(n1386), .IN6(n751), .Q(\fpu_add_frac_dp/n3596 ) );
  AO222X1 U1934 ( .IN1(n1321), .IN2(n101), .IN3(n2460), .IN4(n262), .IN5(n1386), .IN6(n727), .Q(\fpu_add_frac_dp/n3595 ) );
  AO222X1 U1935 ( .IN1(n1319), .IN2(n262), .IN3(n2460), .IN4(
        \fpu_add_frac_dp/n2335 ), .IN5(n1385), .IN6(n726), .Q(
        \fpu_add_frac_dp/n3594 ) );
  AO222X1 U1936 ( .IN1(n1320), .IN2(\fpu_add_frac_dp/n2335 ), .IN3(n2460), 
        .IN4(\fpu_add_frac_dp/n2403 ), .IN5(n1385), .IN6(n729), .Q(
        \fpu_add_frac_dp/n3593 ) );
  AO222X1 U1937 ( .IN1(n1322), .IN2(\fpu_add_frac_dp/n2403 ), .IN3(n2460), 
        .IN4(\fpu_add_frac_dp/n2342 ), .IN5(n1385), .IN6(n1090), .Q(
        \fpu_add_frac_dp/n3592 ) );
  AO222X1 U1938 ( .IN1(n1321), .IN2(\fpu_add_frac_dp/n2342 ), .IN3(n2460), 
        .IN4(\fpu_add_frac_dp/n2289 ), .IN5(n1385), .IN6(n740), .Q(
        \fpu_add_frac_dp/n3591 ) );
  AO222X1 U1939 ( .IN1(n1319), .IN2(\fpu_add_frac_dp/n2289 ), .IN3(n2460), 
        .IN4(\fpu_add_frac_dp/n2406 ), .IN5(n1385), .IN6(n739), .Q(
        \fpu_add_frac_dp/n3590 ) );
  AO222X1 U1940 ( .IN1(n1320), .IN2(\fpu_add_frac_dp/n2406 ), .IN3(n2460), 
        .IN4(\fpu_add_frac_dp/n2332 ), .IN5(n1385), .IN6(n741), .Q(
        \fpu_add_frac_dp/n3589 ) );
  AO222X1 U1941 ( .IN1(n1322), .IN2(\fpu_add_frac_dp/n2332 ), .IN3(n2460), 
        .IN4(n177), .IN5(n1385), .IN6(n742), .Q(\fpu_add_frac_dp/n3588 ) );
  AO222X1 U1942 ( .IN1(n1321), .IN2(n177), .IN3(n2460), .IN4(n86), .IN5(n1385), 
        .IN6(n765), .Q(\fpu_add_frac_dp/n3587 ) );
  AO222X1 U1943 ( .IN1(n1319), .IN2(n86), .IN3(n2460), .IN4(n19), .IN5(n1385), 
        .IN6(n767), .Q(\fpu_add_frac_dp/n3586 ) );
  AO222X1 U1944 ( .IN1(n1320), .IN2(n19), .IN3(n2460), .IN4(n673), .IN5(n1385), 
        .IN6(n459), .Q(\fpu_add_frac_dp/n3585 ) );
  AO222X1 U1945 ( .IN1(n1322), .IN2(n673), .IN3(n2460), .IN4(n117), .IN5(n1385), .IN6(n458), .Q(\fpu_add_frac_dp/n3584 ) );
  AO222X1 U1946 ( .IN1(n1321), .IN2(n117), .IN3(n2460), .IN4(n38), .IN5(n1385), 
        .IN6(n462), .Q(\fpu_add_frac_dp/n3583 ) );
  AO222X1 U1947 ( .IN1(n1319), .IN2(n38), .IN3(n2460), .IN4(n83), .IN5(n1384), 
        .IN6(n766), .Q(\fpu_add_frac_dp/n3582 ) );
  AO222X1 U1948 ( .IN1(n1320), .IN2(n83), .IN3(n2460), .IN4(n665), .IN5(n1384), 
        .IN6(n461), .Q(\fpu_add_frac_dp/n3581 ) );
  AO222X1 U1949 ( .IN1(n1322), .IN2(n665), .IN3(n2460), .IN4(n100), .IN5(n1384), .IN6(n464), .Q(\fpu_add_frac_dp/n3580 ) );
  AO222X1 U1950 ( .IN1(n1321), .IN2(n100), .IN3(n2460), .IN4(n667), .IN5(n1384), .IN6(n457), .Q(\fpu_add_frac_dp/n3579 ) );
  AO222X1 U1951 ( .IN1(n1319), .IN2(n667), .IN3(n2460), .IN4(n40), .IN5(n1384), 
        .IN6(n456), .Q(\fpu_add_frac_dp/n3578 ) );
  AO222X1 U1952 ( .IN1(n1320), .IN2(n40), .IN3(n2460), .IN4(n104), .IN5(n1384), 
        .IN6(n451), .Q(\fpu_add_frac_dp/n3577 ) );
  AO222X1 U1953 ( .IN1(n1322), .IN2(n104), .IN3(n2460), .IN4(n175), .IN5(n1384), .IN6(n914), .Q(\fpu_add_frac_dp/n3576 ) );
  AO222X1 U1954 ( .IN1(n1321), .IN2(n175), .IN3(n2460), .IN4(n22), .IN5(n1384), 
        .IN6(n838), .Q(\fpu_add_frac_dp/n3575 ) );
  AO222X1 U1955 ( .IN1(n1319), .IN2(n22), .IN3(n2460), .IN4(n85), .IN5(n1384), 
        .IN6(n837), .Q(\fpu_add_frac_dp/n3574 ) );
  AO222X1 U1956 ( .IN1(n1320), .IN2(n85), .IN3(n2460), .IN4(n313), .IN5(n1384), 
        .IN6(n842), .Q(\fpu_add_frac_dp/n3573 ) );
  AO222X1 U1957 ( .IN1(n1322), .IN2(n313), .IN3(n2460), .IN4(n92), .IN5(n1383), 
        .IN6(n845), .Q(\fpu_add_frac_dp/n3572 ) );
  AO222X1 U1958 ( .IN1(n1321), .IN2(n92), .IN3(n2460), .IN4(n265), .IN5(n1383), 
        .IN6(n836), .Q(\fpu_add_frac_dp/n3571 ) );
  AO222X1 U1959 ( .IN1(n1319), .IN2(n265), .IN3(n2460), .IN4(
        \fpu_add_frac_dp/n2338 ), .IN5(n1383), .IN6(n835), .Q(
        \fpu_add_frac_dp/n3570 ) );
  AO222X1 U1960 ( .IN1(n1320), .IN2(\fpu_add_frac_dp/n2338 ), .IN3(n2460), 
        .IN4(\fpu_add_frac_dp/n2407 ), .IN5(n1383), .IN6(n841), .Q(
        \fpu_add_frac_dp/n3569 ) );
  AO222X1 U1961 ( .IN1(n1322), .IN2(\fpu_add_frac_dp/n2407 ), .IN3(n2460), 
        .IN4(\fpu_add_frac_dp/n2343 ), .IN5(n1383), .IN6(n844), .Q(
        \fpu_add_frac_dp/n3568 ) );
  AO222X1 U1962 ( .IN1(n1321), .IN2(\fpu_add_frac_dp/n2343 ), .IN3(n2460), 
        .IN4(n171), .IN5(n1383), .IN6(n834), .Q(\fpu_add_frac_dp/n3567 ) );
  AO222X1 U1963 ( .IN1(n1319), .IN2(n171), .IN3(n2460), .IN4(n82), .IN5(n1383), 
        .IN6(n833), .Q(\fpu_add_frac_dp/n3566 ) );
  AO222X1 U1964 ( .IN1(n1320), .IN2(n82), .IN3(n2460), .IN4(
        \fpu_add_frac_dp/n2337 ), .IN5(n1383), .IN6(n840), .Q(
        \fpu_add_frac_dp/n3565 ) );
  AO222X1 U1965 ( .IN1(n1322), .IN2(\fpu_add_frac_dp/n2337 ), .IN3(n2460), 
        .IN4(n94), .IN5(n1379), .IN6(n843), .Q(\fpu_add_frac_dp/n3564 ) );
  AO222X1 U1966 ( .IN1(n1321), .IN2(n94), .IN3(n2460), .IN4(n266), .IN5(n1379), 
        .IN6(n832), .Q(\fpu_add_frac_dp/n3563 ) );
  AO222X1 U1967 ( .IN1(n1319), .IN2(n266), .IN3(n2460), .IN4(n87), .IN5(n1379), 
        .IN6(n831), .Q(\fpu_add_frac_dp/n3562 ) );
  AND2X1 U1968 ( .IN1(n1442), .IN2(n2590), .Q(n2460) );
  AO22X1 U1969 ( .IN1(n1426), .IN2(n846), .IN3(n1320), .IN4(n87), .Q(
        \fpu_add_frac_dp/n3561 ) );
  NAND4X0 U1970 ( .IN1(\fpu_add_frac_dp/n599 ), .IN2(n2731), .IN3(n2732), 
        .IN4(n2733), .QN(n2590) );
  OA221X1 U1971 ( .IN1(n2734), .IN2(n2506), .IN3(n2735), .IN4(n2578), .IN5(
        n2736), .Q(n2733) );
  OA22X1 U1972 ( .IN1(n2737), .IN2(n87), .IN3(n2738), .IN4(n2509), .Q(n2736)
         );
  INVX0 U1973 ( .INP(n2739), .ZN(n2509) );
  OA21X1 U1974 ( .IN1(n2740), .IN2(n22), .IN3(\fpu_add_frac_dp/n612 ), .Q(
        n2738) );
  OA21X1 U1975 ( .IN1(\fpu_add_frac_dp/n614 ), .IN2(n175), .IN3(
        \fpu_add_frac_dp/n613 ), .Q(n2740) );
  OA21X1 U1976 ( .IN1(n2741), .IN2(n266), .IN3(\fpu_add_frac_dp/n600 ), .Q(
        n2737) );
  OA21X1 U1977 ( .IN1(\fpu_add_frac_dp/n602 ), .IN2(n94), .IN3(
        \fpu_add_frac_dp/n601 ), .Q(n2741) );
  OA221X1 U1978 ( .IN1(n2742), .IN2(n2743), .IN3(n2744), .IN4(n2473), .IN5(
        n2745), .Q(n2735) );
  OA21X1 U1979 ( .IN1(\fpu_add_frac_dp/n616 ), .IN2(n40), .IN3(
        \fpu_add_frac_dp/n615 ), .Q(n2745) );
  OA221X1 U1980 ( .IN1(\fpu_add_frac_dp/n628 ), .IN2(n2480), .IN3(n2746), 
        .IN4(n2747), .IN5(n2748), .Q(n2744) );
  OA21X1 U1981 ( .IN1(\fpu_add_frac_dp/n627 ), .IN2(\fpu_add_frac_dp/n2332 ), 
        .IN3(\fpu_add_frac_dp/n626 ), .Q(n2748) );
  OA21X1 U1982 ( .IN1(\fpu_add_frac_dp/n630 ), .IN2(\fpu_add_frac_dp/n2342 ), 
        .IN3(\fpu_add_frac_dp/n629 ), .Q(n2746) );
  OA221X1 U1983 ( .IN1(n2749), .IN2(n2544), .IN3(n2750), .IN4(n2751), .IN5(
        n2752), .Q(n2742) );
  OA21X1 U1984 ( .IN1(\fpu_add_frac_dp/n618 ), .IN2(n100), .IN3(
        \fpu_add_frac_dp/n617 ), .Q(n2752) );
  INVX0 U1985 ( .INP(n2541), .ZN(n2751) );
  OA21X1 U1986 ( .IN1(n2753), .IN2(n19), .IN3(\fpu_add_frac_dp/n623 ), .Q(
        n2750) );
  OA21X1 U1987 ( .IN1(\fpu_add_frac_dp/n625 ), .IN2(n86), .IN3(
        \fpu_add_frac_dp/n624 ), .Q(n2753) );
  OA21X1 U1988 ( .IN1(n2754), .IN2(n83), .IN3(\fpu_add_frac_dp/n619 ), .Q(
        n2749) );
  OA21X1 U1989 ( .IN1(n2755), .IN2(n38), .IN3(\fpu_add_frac_dp/n620 ), .Q(
        n2754) );
  OA21X1 U1990 ( .IN1(\fpu_add_frac_dp/n622 ), .IN2(n117), .IN3(
        \fpu_add_frac_dp/n621 ), .Q(n2755) );
  INVX0 U1991 ( .INP(n2530), .ZN(n2506) );
  OA21X1 U1992 ( .IN1(n2756), .IN2(n265), .IN3(\fpu_add_frac_dp/n608 ), .Q(
        n2734) );
  OA21X1 U1993 ( .IN1(\fpu_add_frac_dp/n610 ), .IN2(n92), .IN3(
        \fpu_add_frac_dp/n609 ), .Q(n2756) );
  OA22X1 U1994 ( .IN1(n2757), .IN2(n2577), .IN3(n2758), .IN4(n2569), .Q(n2732)
         );
  OA221X1 U1995 ( .IN1(\fpu_add_frac_dp/n607 ), .IN2(n2513), .IN3(n2759), 
        .IN4(n82), .IN5(\fpu_add_frac_dp/n603 ), .Q(n2758) );
  OA21X1 U1996 ( .IN1(n2760), .IN2(n171), .IN3(\fpu_add_frac_dp/n604 ), .Q(
        n2759) );
  OA21X1 U1997 ( .IN1(\fpu_add_frac_dp/n606 ), .IN2(\fpu_add_frac_dp/n2343 ), 
        .IN3(\fpu_add_frac_dp/n605 ), .Q(n2760) );
  NAND2X0 U1998 ( .IN1(n2596), .IN2(n2462), .QN(n2577) );
  INVX0 U1999 ( .INP(n2578), .ZN(n2462) );
  NAND4X0 U2000 ( .IN1(\fpu_add_frac_dp/n5631 ), .IN2(\fpu_add_frac_dp/n5630 ), 
        .IN3(\fpu_add_frac_dp/n2386 ), .IN4(n2739), .QN(n2578) );
  NOR2X0 U2001 ( .IN1(n85), .IN2(n2567), .QN(n2739) );
  NOR4X0 U2002 ( .IN1(n2473), .IN2(n2747), .IN3(\fpu_add_frac_dp/n2342 ), 
        .IN4(\fpu_add_frac_dp/n2403 ), .QN(n2596) );
  INVX0 U2003 ( .INP(n2540), .ZN(n2747) );
  NOR2X0 U2004 ( .IN1(n2480), .IN2(\fpu_add_frac_dp/n2289 ), .QN(n2540) );
  OR2X1 U2005 ( .IN1(\fpu_add_frac_dp/n2332 ), .IN2(\fpu_add_frac_dp/n2406 ), 
        .Q(n2480) );
  NAND4X0 U2006 ( .IN1(n2476), .IN2(n2541), .IN3(\fpu_add_frac_dp/n2336 ), 
        .IN4(n2761), .QN(n2473) );
  NOR2X0 U2007 ( .IN1(n19), .IN2(n177), .QN(n2761) );
  NOR3X0 U2008 ( .IN1(n2479), .IN2(n2544), .IN3(n83), .QN(n2541) );
  NAND2X0 U2009 ( .IN1(\fpu_add_frac_dp/n5609 ), .IN2(\fpu_add_frac_dp/n2387 ), 
        .QN(n2544) );
  NAND3X0 U2010 ( .IN1(\fpu_add_frac_dp/n2481 ), .IN2(\fpu_add_frac_dp/n2361 ), 
        .IN3(\fpu_add_frac_dp/n658 ), .QN(n2479) );
  INVX0 U2011 ( .INP(n2743), .ZN(n2476) );
  NAND2X0 U2012 ( .IN1(\fpu_add_frac_dp/n5632 ), .IN2(\fpu_add_frac_dp/n2333 ), 
        .QN(n2743) );
  OA221X1 U2013 ( .IN1(\fpu_add_frac_dp/n2335 ), .IN2(n2762), .IN3(n2763), 
        .IN4(n2493), .IN5(\fpu_add_frac_dp/n631 ), .Q(n2757) );
  NAND4X0 U2014 ( .IN1(\fpu_add_frac_dp/n2411 ), .IN2(n2561), .IN3(n2492), 
        .IN4(n2563), .QN(n2493) );
  NOR4X0 U2015 ( .IN1(n594), .IN2(n74), .IN3(\fpu_add_frac_dp/n2339 ), .IN4(
        \fpu_add_frac_dp/n2405 ), .QN(n2563) );
  INVX0 U2016 ( .INP(n2565), .ZN(n2492) );
  INVX0 U2017 ( .INP(n2490), .ZN(n2561) );
  NAND2X0 U2018 ( .IN1(n2494), .IN2(n839), .QN(n2490) );
  INVX0 U2019 ( .INP(n2764), .ZN(n2494) );
  OA221X1 U2020 ( .IN1(n2765), .IN2(n2595), .IN3(n2766), .IN4(n111), .IN5(
        \fpu_add_frac_dp/n644 ), .Q(n2763) );
  OA21X1 U2021 ( .IN1(\fpu_add_frac_dp/n646 ), .IN2(n43), .IN3(
        \fpu_add_frac_dp/n645 ), .Q(n2766) );
  NAND3X0 U2022 ( .IN1(\fpu_add_frac_dp/n2344 ), .IN2(\fpu_add_frac_dp/n2495 ), 
        .IN3(\fpu_add_frac_dp/n664 ), .QN(n2595) );
  AND3X1 U2023 ( .IN1(\fpu_add_frac_dp/n647 ), .IN2(n2767), .IN3(n2768), .Q(
        n2765) );
  OA221X1 U2024 ( .IN1(\fpu_add_frac_dp/n2400 ), .IN2(n2769), .IN3(n2770), 
        .IN4(n2496), .IN5(n2771), .Q(n2768) );
  OR3X1 U2025 ( .IN1(n103), .IN2(n2546), .IN3(n652), .Q(n2771) );
  NAND4X0 U2026 ( .IN1(n2502), .IN2(n2551), .IN3(\fpu_add_frac_dp/n2447 ), 
        .IN4(n2772), .QN(n2546) );
  AND3X1 U2027 ( .IN1(\fpu_add_frac_dp/n668 ), .IN2(\fpu_add_frac_dp/n2513 ), 
        .IN3(\fpu_add_frac_dp/n670 ), .Q(n2772) );
  NOR2X0 U2028 ( .IN1(n90), .IN2(n626), .QN(n2551) );
  NOR4X0 U2029 ( .IN1(n623), .IN2(n12), .IN3(n34), .IN4(n2496), .QN(n2502) );
  NAND2X0 U2030 ( .IN1(\fpu_add_frac_dp/n2519 ), .IN2(n2556), .QN(n2496) );
  OA21X1 U2031 ( .IN1(\fpu_add_ctl/n140 ), .IN2(n12), .IN3(
        \fpu_add_frac_dp/n652 ), .Q(n2770) );
  OA21X1 U2032 ( .IN1(\fpu_add_frac_dp/n2330 ), .IN2(n2773), .IN3(
        \fpu_add_frac_dp/n648 ), .Q(n2769) );
  OA21X1 U2033 ( .IN1(\fpu_add_frac_dp/n650 ), .IN2(n597), .IN3(
        \fpu_add_frac_dp/n649 ), .Q(n2773) );
  NAND2X0 U2034 ( .IN1(n2556), .IN2(n1081), .QN(n2767) );
  NOR3X0 U2035 ( .IN1(\fpu_add_frac_dp/n2330 ), .IN2(\fpu_add_frac_dp/n2400 ), 
        .IN3(n2774), .QN(n2556) );
  INVX0 U2036 ( .INP(n2552), .ZN(n2774) );
  NOR2X0 U2037 ( .IN1(n37), .IN2(n597), .QN(n2552) );
  OA221X1 U2038 ( .IN1(n2775), .IN2(n2764), .IN3(n2776), .IN4(n262), .IN5(
        \fpu_add_frac_dp/n632 ), .Q(n2762) );
  OA21X1 U2039 ( .IN1(\fpu_add_frac_dp/n634 ), .IN2(n101), .IN3(
        \fpu_add_frac_dp/n633 ), .Q(n2776) );
  NAND3X0 U2040 ( .IN1(\fpu_add_frac_dp/n2496 ), .IN2(\fpu_add_frac_dp/n2363 ), 
        .IN3(\fpu_add_frac_dp/n660 ), .QN(n2764) );
  OA221X1 U2041 ( .IN1(n2777), .IN2(n2565), .IN3(\fpu_add_frac_dp/n2313 ), 
        .IN4(n2778), .IN5(\fpu_add_frac_dp/n635 ), .Q(n2775) );
  OA21X1 U2042 ( .IN1(\fpu_add_frac_dp/n2402 ), .IN2(n2779), .IN3(
        \fpu_add_frac_dp/n636 ), .Q(n2778) );
  OA21X1 U2043 ( .IN1(\fpu_add_frac_dp/n638 ), .IN2(n116), .IN3(
        \fpu_add_frac_dp/n637 ), .Q(n2779) );
  NAND4X0 U2044 ( .IN1(\fpu_add_frac_dp/n5619 ), .IN2(\fpu_add_frac_dp/n2470 ), 
        .IN3(n346), .IN4(n710), .QN(n2565) );
  OA21X1 U2045 ( .IN1(n2780), .IN2(n74), .IN3(\fpu_add_frac_dp/n639 ), .Q(
        n2777) );
  OA21X1 U2046 ( .IN1(n2781), .IN2(n594), .IN3(\fpu_add_frac_dp/n640 ), .Q(
        n2780) );
  OA21X1 U2047 ( .IN1(n2782), .IN2(\fpu_add_frac_dp/n2405 ), .IN3(
        \fpu_add_frac_dp/n641 ), .Q(n2781) );
  OA21X1 U2048 ( .IN1(\fpu_add_frac_dp/n2339 ), .IN2(\fpu_add_frac_dp/n643 ), 
        .IN3(\fpu_add_frac_dp/n642 ), .Q(n2782) );
  OR2X1 U2049 ( .IN1(n2567), .IN2(\fpu_add_frac_dp/n611 ), .Q(n2731) );
  NAND4X0 U2050 ( .IN1(\fpu_add_frac_dp/n2416 ), .IN2(\fpu_add_frac_dp/n2345 ), 
        .IN3(\fpu_add_frac_dp/n2290 ), .IN4(n2530), .QN(n2567) );
  NOR3X0 U2051 ( .IN1(n2513), .IN2(\fpu_add_frac_dp/n2338 ), .IN3(n2569), .QN(
        n2530) );
  NAND4X0 U2052 ( .IN1(\fpu_add_frac_dp/n5618 ), .IN2(\fpu_add_frac_dp/n2440 ), 
        .IN3(\fpu_add_frac_dp/n2288 ), .IN4(n654), .QN(n2569) );
  NAND3X0 U2053 ( .IN1(\fpu_add_frac_dp/n2394 ), .IN2(n2535), .IN3(
        \fpu_add_frac_dp/n654 ), .QN(n2513) );
  NOR2X0 U2054 ( .IN1(\fpu_add_frac_dp/n2407 ), .IN2(\fpu_add_frac_dp/n2343 ), 
        .QN(n2535) );
  AO22X1 U2055 ( .IN1(n1426), .IN2(n987), .IN3(n2783), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3560 ) );
  NOR2X0 U2056 ( .IN1(n2784), .IN2(n2785), .QN(n2783) );
  NOR3X0 U2057 ( .IN1(n2786), .IN2(n21), .IN3(n108), .QN(n2785) );
  AO22X1 U2058 ( .IN1(n1426), .IN2(n986), .IN3(n2787), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3559 ) );
  XOR2X1 U2059 ( .IN1(n2788), .IN2(n2784), .Q(n2787) );
  AO22X1 U2060 ( .IN1(n1426), .IN2(n985), .IN3(n2789), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3558 ) );
  NOR2X0 U2061 ( .IN1(n2790), .IN2(n2791), .QN(n2789) );
  AOI21X1 U2062 ( .IN1(n2788), .IN2(n2784), .IN3(n2792), .QN(n2791) );
  AO22X1 U2063 ( .IN1(n1426), .IN2(n984), .IN3(n2793), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3557 ) );
  XOR2X1 U2064 ( .IN1(n2790), .IN2(n2794), .Q(n2793) );
  AO22X1 U2065 ( .IN1(n1426), .IN2(n983), .IN3(n2795), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3556 ) );
  NOR2X0 U2066 ( .IN1(n2796), .IN2(n2797), .QN(n2795) );
  AOI21X1 U2067 ( .IN1(n2794), .IN2(n2790), .IN3(n2798), .QN(n2797) );
  AO22X1 U2068 ( .IN1(n1427), .IN2(n982), .IN3(n2799), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3555 ) );
  XOR2X1 U2069 ( .IN1(n2800), .IN2(n2796), .Q(n2799) );
  AO22X1 U2070 ( .IN1(n1427), .IN2(n981), .IN3(n2801), .IN4(n1435), .Q(
        \fpu_add_frac_dp/n3554 ) );
  NOR2X0 U2071 ( .IN1(n2802), .IN2(n2803), .QN(n2801) );
  OA21X1 U2072 ( .IN1(n2804), .IN2(n2805), .IN3(n2806), .Q(n2803) );
  AO22X1 U2073 ( .IN1(n1427), .IN2(n980), .IN3(n2807), .IN4(n1435), .Q(
        \fpu_add_frac_dp/n3553 ) );
  XOR2X1 U2074 ( .IN1(n2808), .IN2(n2809), .Q(n2807) );
  AO22X1 U2075 ( .IN1(n1427), .IN2(n979), .IN3(n2810), .IN4(n1435), .Q(
        \fpu_add_frac_dp/n3552 ) );
  NOR2X0 U2076 ( .IN1(n2811), .IN2(n2812), .QN(n2810) );
  OA21X1 U2077 ( .IN1(n2809), .IN2(n2808), .IN3(n2813), .Q(n2812) );
  AO22X1 U2078 ( .IN1(n1427), .IN2(n977), .IN3(n2814), .IN4(n1435), .Q(
        \fpu_add_frac_dp/n3551 ) );
  XOR2X1 U2079 ( .IN1(n2815), .IN2(n2811), .Q(n2814) );
  AO22X1 U2080 ( .IN1(n1427), .IN2(n976), .IN3(n2816), .IN4(n1435), .Q(
        \fpu_add_frac_dp/n3550 ) );
  NOR2X0 U2081 ( .IN1(n2817), .IN2(n2818), .QN(n2816) );
  OA21X1 U2082 ( .IN1(n2819), .IN2(n2820), .IN3(n2821), .Q(n2818) );
  AO22X1 U2083 ( .IN1(n1427), .IN2(n975), .IN3(n2822), .IN4(n1435), .Q(
        \fpu_add_frac_dp/n3549 ) );
  XOR2X1 U2084 ( .IN1(n2823), .IN2(n2824), .Q(n2822) );
  AO22X1 U2085 ( .IN1(n1427), .IN2(n974), .IN3(n2825), .IN4(n1435), .Q(
        \fpu_add_frac_dp/n3548 ) );
  NOR2X0 U2086 ( .IN1(n2826), .IN2(n2827), .QN(n2825) );
  OA21X1 U2087 ( .IN1(n2824), .IN2(n2823), .IN3(n2828), .Q(n2827) );
  AO22X1 U2088 ( .IN1(n1427), .IN2(n973), .IN3(n2829), .IN4(n1435), .Q(
        \fpu_add_frac_dp/n3547 ) );
  XOR2X1 U2089 ( .IN1(n2830), .IN2(n2826), .Q(n2829) );
  AO22X1 U2090 ( .IN1(n1427), .IN2(n972), .IN3(n2831), .IN4(n1435), .Q(
        \fpu_add_frac_dp/n3546 ) );
  NOR2X0 U2091 ( .IN1(n2832), .IN2(n2833), .QN(n2831) );
  AOI21X1 U2092 ( .IN1(n2830), .IN2(n2826), .IN3(n2834), .QN(n2833) );
  AO22X1 U2093 ( .IN1(n1427), .IN2(n971), .IN3(n2835), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3545 ) );
  XOR2X1 U2094 ( .IN1(n2832), .IN2(n2836), .Q(n2835) );
  AO22X1 U2095 ( .IN1(n1428), .IN2(n970), .IN3(n2837), .IN4(n1435), .Q(
        \fpu_add_frac_dp/n3544 ) );
  NOR2X0 U2096 ( .IN1(n2838), .IN2(n2839), .QN(n2837) );
  AOI21X1 U2097 ( .IN1(n2836), .IN2(n2832), .IN3(n2840), .QN(n2839) );
  AO22X1 U2098 ( .IN1(n1427), .IN2(n969), .IN3(n2841), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3543 ) );
  XOR2X1 U2099 ( .IN1(n2842), .IN2(n2838), .Q(n2841) );
  AO22X1 U2100 ( .IN1(n1428), .IN2(n1062), .IN3(n2843), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3542 ) );
  NOR2X0 U2101 ( .IN1(n2844), .IN2(n2845), .QN(n2843) );
  AOI21X1 U2102 ( .IN1(n2842), .IN2(n2838), .IN3(n2846), .QN(n2845) );
  AO22X1 U2103 ( .IN1(n1428), .IN2(n1061), .IN3(n2847), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3541 ) );
  XOR2X1 U2104 ( .IN1(n2844), .IN2(n2848), .Q(n2847) );
  AO22X1 U2105 ( .IN1(n1428), .IN2(n1060), .IN3(n2849), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3540 ) );
  NOR2X0 U2106 ( .IN1(n2850), .IN2(n2851), .QN(n2849) );
  AOI21X1 U2107 ( .IN1(n2848), .IN2(n2844), .IN3(n2852), .QN(n2851) );
  AO22X1 U2108 ( .IN1(n1427), .IN2(n1059), .IN3(n2853), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3539 ) );
  XOR2X1 U2109 ( .IN1(n2854), .IN2(n2850), .Q(n2853) );
  AO22X1 U2110 ( .IN1(n1427), .IN2(n1058), .IN3(n2855), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3538 ) );
  NOR2X0 U2111 ( .IN1(n2856), .IN2(n2857), .QN(n2855) );
  AOI21X1 U2112 ( .IN1(n2854), .IN2(n2850), .IN3(n2858), .QN(n2857) );
  AO22X1 U2113 ( .IN1(n1428), .IN2(n1057), .IN3(n2859), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3537 ) );
  XOR2X1 U2114 ( .IN1(n2860), .IN2(n2861), .Q(n2859) );
  AO22X1 U2115 ( .IN1(n1428), .IN2(n1056), .IN3(n2862), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3536 ) );
  NOR2X0 U2116 ( .IN1(n2863), .IN2(n2864), .QN(n2862) );
  OA21X1 U2117 ( .IN1(n2861), .IN2(n2860), .IN3(n2865), .Q(n2864) );
  AO22X1 U2118 ( .IN1(n1428), .IN2(n1055), .IN3(n2866), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3535 ) );
  XOR2X1 U2119 ( .IN1(n2867), .IN2(n2863), .Q(n2866) );
  AO22X1 U2120 ( .IN1(n1428), .IN2(n1054), .IN3(n2868), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3534 ) );
  NOR2X0 U2121 ( .IN1(n2869), .IN2(n2870), .QN(n2868) );
  OA21X1 U2122 ( .IN1(n2871), .IN2(n2872), .IN3(n2873), .Q(n2870) );
  AO22X1 U2123 ( .IN1(n1429), .IN2(n1053), .IN3(n2874), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3533 ) );
  XOR2X1 U2124 ( .IN1(n2875), .IN2(n2876), .Q(n2874) );
  AO22X1 U2125 ( .IN1(n1427), .IN2(n1052), .IN3(n2877), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3532 ) );
  NOR2X0 U2126 ( .IN1(n2878), .IN2(n2879), .QN(n2877) );
  OA21X1 U2127 ( .IN1(n2876), .IN2(n2875), .IN3(n2880), .Q(n2879) );
  INVX0 U2128 ( .INP(n2881), .ZN(n2876) );
  AO22X1 U2129 ( .IN1(n1429), .IN2(n1051), .IN3(n1442), .IN4(n2882), .Q(
        \fpu_add_frac_dp/n3531 ) );
  XOR3X1 U2130 ( .IN1(n2883), .IN2(n2884), .IN3(n2885), .Q(n2882) );
  AO22X1 U2131 ( .IN1(n1428), .IN2(n1050), .IN3(n2886), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3530 ) );
  OA21X1 U2132 ( .IN1(n2887), .IN2(n2888), .IN3(n2889), .Q(n2886) );
  AO22X1 U2133 ( .IN1(n1429), .IN2(n1049), .IN3(n2890), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3529 ) );
  XOR2X1 U2134 ( .IN1(n2891), .IN2(n2892), .Q(n2890) );
  AO22X1 U2135 ( .IN1(n1428), .IN2(n1048), .IN3(n2893), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3528 ) );
  NOR2X0 U2136 ( .IN1(n2894), .IN2(n2895), .QN(n2893) );
  AOI21X1 U2137 ( .IN1(n2891), .IN2(n2892), .IN3(n2896), .QN(n2895) );
  AO22X1 U2138 ( .IN1(n1429), .IN2(n1047), .IN3(n2897), .IN4(n1436), .Q(
        \fpu_add_frac_dp/n3527 ) );
  XOR2X1 U2139 ( .IN1(n2894), .IN2(n2898), .Q(n2897) );
  AO22X1 U2140 ( .IN1(n1428), .IN2(n1046), .IN3(n2899), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3526 ) );
  NOR2X0 U2141 ( .IN1(n2900), .IN2(n2901), .QN(n2899) );
  AOI21X1 U2142 ( .IN1(n2898), .IN2(n2894), .IN3(n2902), .QN(n2901) );
  AO22X1 U2143 ( .IN1(n1429), .IN2(n1045), .IN3(n2903), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3525 ) );
  XOR2X1 U2144 ( .IN1(n2904), .IN2(n2900), .Q(n2903) );
  AO22X1 U2145 ( .IN1(n1428), .IN2(n1044), .IN3(n2905), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3524 ) );
  NOR2X0 U2146 ( .IN1(n2906), .IN2(n2907), .QN(n2905) );
  AOI21X1 U2147 ( .IN1(n2904), .IN2(n2900), .IN3(n2908), .QN(n2907) );
  AO22X1 U2148 ( .IN1(n1429), .IN2(n1043), .IN3(n2909), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3523 ) );
  XOR2X1 U2149 ( .IN1(n2906), .IN2(n2910), .Q(n2909) );
  AO22X1 U2150 ( .IN1(n1429), .IN2(n1042), .IN3(n2911), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3522 ) );
  NOR2X0 U2151 ( .IN1(n2912), .IN2(n2913), .QN(n2911) );
  AOI21X1 U2152 ( .IN1(n2910), .IN2(n2906), .IN3(n2914), .QN(n2913) );
  AO22X1 U2153 ( .IN1(n1428), .IN2(n968), .IN3(n2915), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3521 ) );
  XOR2X1 U2154 ( .IN1(n2916), .IN2(n2912), .Q(n2915) );
  AO22X1 U2155 ( .IN1(n1429), .IN2(n967), .IN3(n2917), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3520 ) );
  NOR2X0 U2156 ( .IN1(n2918), .IN2(n2919), .QN(n2917) );
  AOI21X1 U2157 ( .IN1(n2916), .IN2(n2912), .IN3(n2920), .QN(n2919) );
  AO22X1 U2158 ( .IN1(n1419), .IN2(n966), .IN3(n2921), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3519 ) );
  XOR2X1 U2159 ( .IN1(n2918), .IN2(n2922), .Q(n2921) );
  AO22X1 U2160 ( .IN1(n1416), .IN2(n965), .IN3(n2923), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3518 ) );
  NOR2X0 U2161 ( .IN1(n2924), .IN2(n2925), .QN(n2923) );
  AOI21X1 U2162 ( .IN1(n2922), .IN2(n2918), .IN3(n2926), .QN(n2925) );
  AO22X1 U2163 ( .IN1(n1416), .IN2(n964), .IN3(n2927), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3517 ) );
  XOR2X1 U2164 ( .IN1(n2928), .IN2(n2924), .Q(n2927) );
  AO22X1 U2165 ( .IN1(n1416), .IN2(n1041), .IN3(n2929), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3516 ) );
  NOR2X0 U2166 ( .IN1(n2930), .IN2(n2931), .QN(n2929) );
  AOI21X1 U2167 ( .IN1(n2928), .IN2(n2924), .IN3(n2932), .QN(n2931) );
  AO22X1 U2168 ( .IN1(n1416), .IN2(n1040), .IN3(n2933), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3515 ) );
  XOR2X1 U2169 ( .IN1(n2934), .IN2(n2935), .Q(n2933) );
  AO22X1 U2170 ( .IN1(n1416), .IN2(n1039), .IN3(n2936), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3514 ) );
  NOR2X0 U2171 ( .IN1(n2937), .IN2(n2938), .QN(n2936) );
  OA21X1 U2172 ( .IN1(n2935), .IN2(n2934), .IN3(n2939), .Q(n2938) );
  INVX0 U2173 ( .INP(n2940), .ZN(n2935) );
  AO22X1 U2174 ( .IN1(n1416), .IN2(n1038), .IN3(n2941), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3513 ) );
  XOR2X1 U2175 ( .IN1(n2942), .IN2(n2937), .Q(n2941) );
  AO22X1 U2176 ( .IN1(n1416), .IN2(n1037), .IN3(n2943), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3512 ) );
  NOR2X0 U2177 ( .IN1(n2944), .IN2(n2945), .QN(n2943) );
  AOI21X1 U2178 ( .IN1(n2942), .IN2(n2937), .IN3(n2946), .QN(n2945) );
  AO22X1 U2179 ( .IN1(n1416), .IN2(n1036), .IN3(n2947), .IN4(n1437), .Q(
        \fpu_add_frac_dp/n3511 ) );
  XOR2X1 U2180 ( .IN1(n2944), .IN2(n2948), .Q(n2947) );
  AO22X1 U2181 ( .IN1(n1416), .IN2(n1035), .IN3(n2949), .IN4(n1438), .Q(
        \fpu_add_frac_dp/n3510 ) );
  NOR2X0 U2182 ( .IN1(n2950), .IN2(n2951), .QN(n2949) );
  AOI21X1 U2183 ( .IN1(n2948), .IN2(n2944), .IN3(n2952), .QN(n2951) );
  AO21X1 U2184 ( .IN1(n1406), .IN2(n1006), .IN3(n2953), .Q(
        \fpu_add_frac_dp/n3509 ) );
  MUX21X1 U2185 ( .IN1(n2954), .IN2(n2955), .S(n2950), .Q(n2953) );
  NOR2X0 U2186 ( .IN1(n1745), .IN2(n2956), .QN(n2955) );
  AO22X1 U2187 ( .IN1(n1443), .IN2(n2957), .IN3(n1410), .IN4(n1186), .Q(
        \fpu_add_frac_dp/n3508 ) );
  AO22X1 U2188 ( .IN1(n1416), .IN2(n65), .IN3(n1442), .IN4(n2958), .Q(
        \fpu_add_frac_dp/n3507 ) );
  AO21X1 U2189 ( .IN1(n2959), .IN2(n2960), .IN3(n492), .Q(n2958) );
  OAI22X1 U2190 ( .IN1(n1745), .IN2(n2959), .IN3(n2046), .IN4(
        \fpu_add_frac_dp/n132 ), .QN(\fpu_add_frac_dp/n3506 ) );
  AO22X1 U2191 ( .IN1(n1416), .IN2(n1305), .IN3(n1442), .IN4(n2961), .Q(
        \fpu_add_frac_dp/n3505 ) );
  NAND2X0 U2192 ( .IN1(\fpu_add_ctl/n85 ), .IN2(n2962), .QN(n2961) );
  AO22X1 U2193 ( .IN1(n1448), .IN2(n2963), .IN3(n1410), .IN4(n579), .Q(
        \fpu_add_frac_dp/n3504 ) );
  AO22X1 U2194 ( .IN1(n1417), .IN2(n1248), .IN3(n2954), .IN4(n2950), .Q(
        \fpu_add_frac_dp/n3503 ) );
  AO22X1 U2195 ( .IN1(n1448), .IN2(n956), .IN3(n1410), .IN4(n544), .Q(
        \fpu_add_frac_dp/n3502 ) );
  AO22X1 U2196 ( .IN1(n1417), .IN2(n978), .IN3(n1442), .IN4(n2964), .Q(
        \fpu_add_frac_dp/n3501 ) );
  AO22X1 U2197 ( .IN1(n1449), .IN2(n2965), .IN3(n1410), .IN4(n543), .Q(
        \fpu_add_frac_dp/n3500 ) );
  AO22X1 U2198 ( .IN1(n1448), .IN2(n2966), .IN3(n1410), .IN4(n542), .Q(
        \fpu_add_frac_dp/n3499 ) );
  AO22X1 U2199 ( .IN1(n1449), .IN2(n2967), .IN3(n1410), .IN4(n541), .Q(
        \fpu_add_frac_dp/n3498 ) );
  AO22X1 U2200 ( .IN1(n1448), .IN2(n2968), .IN3(n1410), .IN4(n540), .Q(
        \fpu_add_frac_dp/n3497 ) );
  AO22X1 U2201 ( .IN1(n1448), .IN2(n2969), .IN3(n1410), .IN4(n539), .Q(
        \fpu_add_frac_dp/n3496 ) );
  AO22X1 U2202 ( .IN1(n1448), .IN2(n2970), .IN3(n1410), .IN4(n538), .Q(
        \fpu_add_frac_dp/n3495 ) );
  AO22X1 U2203 ( .IN1(n1448), .IN2(n2971), .IN3(n1410), .IN4(n537), .Q(
        \fpu_add_frac_dp/n3494 ) );
  AO22X1 U2204 ( .IN1(n1448), .IN2(n2972), .IN3(n1410), .IN4(n536), .Q(
        \fpu_add_frac_dp/n3493 ) );
  AO22X1 U2205 ( .IN1(n1448), .IN2(n2973), .IN3(n1411), .IN4(n908), .Q(
        \fpu_add_frac_dp/n3492 ) );
  AO22X1 U2206 ( .IN1(n1746), .IN2(n2786), .IN3(n1411), .IN4(n955), .Q(
        \fpu_add_frac_dp/n3491 ) );
  AO22X1 U2207 ( .IN1(n1448), .IN2(n2788), .IN3(n1411), .IN4(n954), .Q(
        \fpu_add_frac_dp/n3490 ) );
  AO22X1 U2208 ( .IN1(n1448), .IN2(n2792), .IN3(n1411), .IN4(n953), .Q(
        \fpu_add_frac_dp/n3489 ) );
  AO22X1 U2209 ( .IN1(n1448), .IN2(n2794), .IN3(n1411), .IN4(n952), .Q(
        \fpu_add_frac_dp/n3488 ) );
  AO22X1 U2210 ( .IN1(n1448), .IN2(n2798), .IN3(n1411), .IN4(n951), .Q(
        \fpu_add_frac_dp/n3487 ) );
  AO22X1 U2211 ( .IN1(n1448), .IN2(n2800), .IN3(n1411), .IN4(n950), .Q(
        \fpu_add_frac_dp/n3486 ) );
  AO22X1 U2212 ( .IN1(n1746), .IN2(n2974), .IN3(n1411), .IN4(n949), .Q(
        \fpu_add_frac_dp/n3485 ) );
  AO22X1 U2213 ( .IN1(n1448), .IN2(n2975), .IN3(n1411), .IN4(n948), .Q(
        \fpu_add_frac_dp/n3484 ) );
  AO22X1 U2214 ( .IN1(n1448), .IN2(n2976), .IN3(n1411), .IN4(n947), .Q(
        \fpu_add_frac_dp/n3483 ) );
  AO22X1 U2215 ( .IN1(n1448), .IN2(n2815), .IN3(n1411), .IN4(n946), .Q(
        \fpu_add_frac_dp/n3482 ) );
  AO22X1 U2216 ( .IN1(n1746), .IN2(n2977), .IN3(n1411), .IN4(n945), .Q(
        \fpu_add_frac_dp/n3481 ) );
  AO22X1 U2217 ( .IN1(n1448), .IN2(n2978), .IN3(n1411), .IN4(n944), .Q(
        \fpu_add_frac_dp/n3480 ) );
  AO22X1 U2218 ( .IN1(n1746), .IN2(n2979), .IN3(n1411), .IN4(n943), .Q(
        \fpu_add_frac_dp/n3479 ) );
  AO22X1 U2219 ( .IN1(n1746), .IN2(n2830), .IN3(n1412), .IN4(n942), .Q(
        \fpu_add_frac_dp/n3478 ) );
  AO22X1 U2220 ( .IN1(n1746), .IN2(n2834), .IN3(n1412), .IN4(n941), .Q(
        \fpu_add_frac_dp/n3477 ) );
  AO22X1 U2221 ( .IN1(n1746), .IN2(n2836), .IN3(n1412), .IN4(n940), .Q(
        \fpu_add_frac_dp/n3476 ) );
  AO22X1 U2222 ( .IN1(n1746), .IN2(n2840), .IN3(n1412), .IN4(n939), .Q(
        \fpu_add_frac_dp/n3475 ) );
  AO22X1 U2223 ( .IN1(n1746), .IN2(n2842), .IN3(n1412), .IN4(n938), .Q(
        \fpu_add_frac_dp/n3474 ) );
  AO22X1 U2224 ( .IN1(n1447), .IN2(n2846), .IN3(n1412), .IN4(n881), .Q(
        \fpu_add_frac_dp/n3473 ) );
  AO22X1 U2225 ( .IN1(n1449), .IN2(n2848), .IN3(n1412), .IN4(n880), .Q(
        \fpu_add_frac_dp/n3472 ) );
  AO22X1 U2226 ( .IN1(n1746), .IN2(n2852), .IN3(n1412), .IN4(n879), .Q(
        \fpu_add_frac_dp/n3471 ) );
  AO22X1 U2227 ( .IN1(n1449), .IN2(n2854), .IN3(n1412), .IN4(n878), .Q(
        \fpu_add_frac_dp/n3470 ) );
  AO22X1 U2228 ( .IN1(n1746), .IN2(n2858), .IN3(n1412), .IN4(n877), .Q(
        \fpu_add_frac_dp/n3469 ) );
  AO22X1 U2229 ( .IN1(n1449), .IN2(n2980), .IN3(n1412), .IN4(n876), .Q(
        \fpu_add_frac_dp/n3468 ) );
  AO22X1 U2230 ( .IN1(n1449), .IN2(n2981), .IN3(n1412), .IN4(n875), .Q(
        \fpu_add_frac_dp/n3467 ) );
  AO22X1 U2231 ( .IN1(n1746), .IN2(n2867), .IN3(n1412), .IN4(n874), .Q(
        \fpu_add_frac_dp/n3466 ) );
  AO22X1 U2232 ( .IN1(n1449), .IN2(n2982), .IN3(n1412), .IN4(n873), .Q(
        \fpu_add_frac_dp/n3465 ) );
  AO22X1 U2233 ( .IN1(n1447), .IN2(n2881), .IN3(n1413), .IN4(n872), .Q(
        \fpu_add_frac_dp/n3464 ) );
  AO22X1 U2234 ( .IN1(n1449), .IN2(n2983), .IN3(n1413), .IN4(n871), .Q(
        \fpu_add_frac_dp/n3463 ) );
  AO22X1 U2235 ( .IN1(n1447), .IN2(n2984), .IN3(n1413), .IN4(n870), .Q(
        \fpu_add_frac_dp/n3462 ) );
  AO22X1 U2236 ( .IN1(n1447), .IN2(n2888), .IN3(n1413), .IN4(n869), .Q(
        \fpu_add_frac_dp/n3461 ) );
  AO22X1 U2237 ( .IN1(n1447), .IN2(n2891), .IN3(n1413), .IN4(n868), .Q(
        \fpu_add_frac_dp/n3460 ) );
  AO22X1 U2238 ( .IN1(n1447), .IN2(n2896), .IN3(n1413), .IN4(n867), .Q(
        \fpu_add_frac_dp/n3459 ) );
  AO22X1 U2239 ( .IN1(n1447), .IN2(n2898), .IN3(n1413), .IN4(n866), .Q(
        \fpu_add_frac_dp/n3458 ) );
  AO22X1 U2240 ( .IN1(n1447), .IN2(n2902), .IN3(n1413), .IN4(n865), .Q(
        \fpu_add_frac_dp/n3457 ) );
  AO22X1 U2241 ( .IN1(n1447), .IN2(n2904), .IN3(n1413), .IN4(n864), .Q(
        \fpu_add_frac_dp/n3456 ) );
  AO22X1 U2242 ( .IN1(n1447), .IN2(n2908), .IN3(n1413), .IN4(n863), .Q(
        \fpu_add_frac_dp/n3455 ) );
  AO22X1 U2243 ( .IN1(n1447), .IN2(n2910), .IN3(n1413), .IN4(n862), .Q(
        \fpu_add_frac_dp/n3454 ) );
  AO22X1 U2244 ( .IN1(n1447), .IN2(n2914), .IN3(n1413), .IN4(n861), .Q(
        \fpu_add_frac_dp/n3453 ) );
  AO22X1 U2245 ( .IN1(n1447), .IN2(n2916), .IN3(n1413), .IN4(n503), .Q(
        \fpu_add_frac_dp/n3452 ) );
  AO22X1 U2246 ( .IN1(n1447), .IN2(n2920), .IN3(n1413), .IN4(n502), .Q(
        \fpu_add_frac_dp/n3451 ) );
  AO22X1 U2247 ( .IN1(n1446), .IN2(n2922), .IN3(n1414), .IN4(n501), .Q(
        \fpu_add_frac_dp/n3450 ) );
  AO22X1 U2248 ( .IN1(n1447), .IN2(n2926), .IN3(n1414), .IN4(n500), .Q(
        \fpu_add_frac_dp/n3449 ) );
  AO22X1 U2249 ( .IN1(n1447), .IN2(n2928), .IN3(n1414), .IN4(n499), .Q(
        \fpu_add_frac_dp/n3448 ) );
  AO22X1 U2250 ( .IN1(n1447), .IN2(n2932), .IN3(n1414), .IN4(n498), .Q(
        \fpu_add_frac_dp/n3447 ) );
  AO22X1 U2251 ( .IN1(n1446), .IN2(n2940), .IN3(n1414), .IN4(n497), .Q(
        \fpu_add_frac_dp/n3446 ) );
  AO22X1 U2252 ( .IN1(n1447), .IN2(n2985), .IN3(n1414), .IN4(n496), .Q(
        \fpu_add_frac_dp/n3445 ) );
  AO22X1 U2253 ( .IN1(n1446), .IN2(n2942), .IN3(n1414), .IN4(n495), .Q(
        \fpu_add_frac_dp/n3444 ) );
  AO22X1 U2254 ( .IN1(n1446), .IN2(n2946), .IN3(n1414), .IN4(n494), .Q(
        \fpu_add_frac_dp/n3443 ) );
  AO22X1 U2255 ( .IN1(n1446), .IN2(n2948), .IN3(n1414), .IN4(n860), .Q(
        \fpu_add_frac_dp/n3442 ) );
  AO22X1 U2256 ( .IN1(n1446), .IN2(n2952), .IN3(n1414), .IN4(n493), .Q(
        \fpu_add_frac_dp/n3441 ) );
  AO21X1 U2257 ( .IN1(n1405), .IN2(n907), .IN3(n2954), .Q(
        \fpu_add_frac_dp/n3440 ) );
  NOR2X0 U2258 ( .IN1(n1745), .IN2(n2986), .QN(n2954) );
  AO22X1 U2259 ( .IN1(n1446), .IN2(n2987), .IN3(n1406), .IN4(n859), .Q(
        \fpu_add_frac_dp/n3439 ) );
  AO22X1 U2260 ( .IN1(n1421), .IN2(n925), .IN3(n2988), .IN4(n2989), .Q(
        \fpu_add_frac_dp/n3438 ) );
  AO22X1 U2261 ( .IN1(n1421), .IN2(n551), .IN3(n2990), .IN4(n2989), .Q(
        \fpu_add_frac_dp/n3437 ) );
  AO22X1 U2262 ( .IN1(n1421), .IN2(n924), .IN3(n2991), .IN4(n2989), .Q(
        \fpu_add_frac_dp/n3436 ) );
  AO22X1 U2263 ( .IN1(n1421), .IN2(n923), .IN3(n2992), .IN4(n2989), .Q(
        \fpu_add_frac_dp/n3435 ) );
  AO22X1 U2264 ( .IN1(n1421), .IN2(n922), .IN3(n2993), .IN4(n2994), .Q(
        \fpu_add_frac_dp/n3434 ) );
  AO22X1 U2265 ( .IN1(n1421), .IN2(n921), .IN3(n2995), .IN4(n2994), .Q(
        \fpu_add_frac_dp/n3433 ) );
  AO22X1 U2266 ( .IN1(n1421), .IN2(n920), .IN3(n2996), .IN4(n2994), .Q(
        \fpu_add_frac_dp/n3432 ) );
  AO22X1 U2267 ( .IN1(n1421), .IN2(n919), .IN3(n2997), .IN4(n2994), .Q(
        \fpu_add_frac_dp/n3431 ) );
  AO21X1 U2268 ( .IN1(n1405), .IN2(n1003), .IN3(n2998), .Q(
        \fpu_add_frac_dp/n3430 ) );
  AO21X1 U2269 ( .IN1(n1405), .IN2(n1002), .IN3(n2999), .Q(
        \fpu_add_frac_dp/n3429 ) );
  AO222X1 U2270 ( .IN1(n3000), .IN2(n2994), .IN3(n3001), .IN4(n2991), .IN5(
        n1379), .IN6(n535), .Q(\fpu_add_frac_dp/n3428 ) );
  AO222X1 U2271 ( .IN1(n3002), .IN2(n2994), .IN3(n3001), .IN4(n2992), .IN5(
        n1379), .IN6(n534), .Q(\fpu_add_frac_dp/n3427 ) );
  AO222X1 U2272 ( .IN1(n3003), .IN2(n2993), .IN3(n3004), .IN4(n2994), .IN5(
        n1379), .IN6(n533), .Q(\fpu_add_frac_dp/n3426 ) );
  AO222X1 U2273 ( .IN1(n3003), .IN2(n2995), .IN3(n3005), .IN4(n2994), .IN5(
        n1379), .IN6(n532), .Q(\fpu_add_frac_dp/n3425 ) );
  AO222X1 U2274 ( .IN1(n3003), .IN2(n2996), .IN3(n3006), .IN4(n2994), .IN5(
        n1379), .IN6(n531), .Q(\fpu_add_frac_dp/n3424 ) );
  AO222X1 U2275 ( .IN1(n3003), .IN2(n2997), .IN3(n3007), .IN4(n2994), .IN5(
        n1379), .IN6(n530), .Q(\fpu_add_frac_dp/n3423 ) );
  AO222X1 U2276 ( .IN1(n3008), .IN2(n3003), .IN3(n3009), .IN4(n2994), .IN5(
        n1379), .IN6(n529), .Q(\fpu_add_frac_dp/n3422 ) );
  AO222X1 U2277 ( .IN1(n3010), .IN2(n3003), .IN3(n3011), .IN4(n2994), .IN5(
        n1379), .IN6(n528), .Q(\fpu_add_frac_dp/n3421 ) );
  AO222X1 U2278 ( .IN1(n3000), .IN2(n3003), .IN3(n3012), .IN4(n2994), .IN5(
        n1380), .IN6(n527), .Q(\fpu_add_frac_dp/n3420 ) );
  AO222X1 U2279 ( .IN1(n3002), .IN2(n3003), .IN3(n3013), .IN4(n2994), .IN5(
        n1380), .IN6(n526), .Q(\fpu_add_frac_dp/n3419 ) );
  AO222X1 U2280 ( .IN1(n3004), .IN2(n3003), .IN3(n3014), .IN4(n2994), .IN5(
        n1380), .IN6(n525), .Q(\fpu_add_frac_dp/n3418 ) );
  AO222X1 U2281 ( .IN1(n3005), .IN2(n3003), .IN3(n2994), .IN4(n3015), .IN5(
        n1380), .IN6(n524), .Q(\fpu_add_frac_dp/n3417 ) );
  AO222X1 U2282 ( .IN1(n3006), .IN2(n3003), .IN3(n2994), .IN4(n3016), .IN5(
        n1380), .IN6(n523), .Q(\fpu_add_frac_dp/n3416 ) );
  AO222X1 U2283 ( .IN1(n3007), .IN2(n3003), .IN3(n2994), .IN4(n3017), .IN5(
        n1380), .IN6(n522), .Q(\fpu_add_frac_dp/n3415 ) );
  AO222X1 U2284 ( .IN1(n3009), .IN2(n3003), .IN3(n2994), .IN4(n3018), .IN5(
        n1380), .IN6(n521), .Q(\fpu_add_frac_dp/n3414 ) );
  AO222X1 U2285 ( .IN1(n3011), .IN2(n3003), .IN3(n2994), .IN4(n3019), .IN5(
        n1380), .IN6(n520), .Q(\fpu_add_frac_dp/n3413 ) );
  AO222X1 U2286 ( .IN1(n3012), .IN2(n3003), .IN3(n2994), .IN4(n3020), .IN5(
        n1380), .IN6(n519), .Q(\fpu_add_frac_dp/n3412 ) );
  AO222X1 U2287 ( .IN1(n3013), .IN2(n3003), .IN3(n2994), .IN4(n3021), .IN5(
        n1380), .IN6(n518), .Q(\fpu_add_frac_dp/n3411 ) );
  AO222X1 U2288 ( .IN1(n3014), .IN2(n3003), .IN3(n2994), .IN4(n3022), .IN5(
        n1380), .IN6(n517), .Q(\fpu_add_frac_dp/n3410 ) );
  AO222X1 U2289 ( .IN1(n3003), .IN2(n3015), .IN3(n2994), .IN4(n3023), .IN5(
        n1380), .IN6(n489), .Q(\fpu_add_frac_dp/n3409 ) );
  AO222X1 U2290 ( .IN1(n3003), .IN2(n3016), .IN3(n2994), .IN4(n3024), .IN5(
        n1381), .IN6(n488), .Q(\fpu_add_frac_dp/n3408 ) );
  AO222X1 U2291 ( .IN1(n3003), .IN2(n3017), .IN3(n2994), .IN4(n3025), .IN5(
        n1381), .IN6(n487), .Q(\fpu_add_frac_dp/n3407 ) );
  AO222X1 U2292 ( .IN1(n3003), .IN2(n3018), .IN3(n2994), .IN4(n3026), .IN5(
        n1381), .IN6(n486), .Q(\fpu_add_frac_dp/n3406 ) );
  AO222X1 U2293 ( .IN1(n3003), .IN2(n3019), .IN3(n2994), .IN4(n3027), .IN5(
        n1381), .IN6(n485), .Q(\fpu_add_frac_dp/n3405 ) );
  AO222X1 U2294 ( .IN1(n3003), .IN2(n3020), .IN3(n2994), .IN4(n3028), .IN5(
        n1381), .IN6(n484), .Q(\fpu_add_frac_dp/n3404 ) );
  AO222X1 U2295 ( .IN1(n3003), .IN2(n3021), .IN3(n2994), .IN4(n3029), .IN5(
        n1381), .IN6(n483), .Q(\fpu_add_frac_dp/n3403 ) );
  AO222X1 U2296 ( .IN1(n3003), .IN2(n3022), .IN3(n2994), .IN4(n3030), .IN5(
        n1381), .IN6(n482), .Q(\fpu_add_frac_dp/n3402 ) );
  AO222X1 U2297 ( .IN1(n3003), .IN2(n3023), .IN3(n2994), .IN4(n3031), .IN5(
        n1381), .IN6(n481), .Q(\fpu_add_frac_dp/n3401 ) );
  AO222X1 U2298 ( .IN1(n3003), .IN2(n3024), .IN3(n2994), .IN4(n3032), .IN5(
        n1381), .IN6(n480), .Q(\fpu_add_frac_dp/n3400 ) );
  AO222X1 U2299 ( .IN1(n3003), .IN2(n3025), .IN3(n2994), .IN4(n3033), .IN5(
        n1381), .IN6(n479), .Q(\fpu_add_frac_dp/n3399 ) );
  AO222X1 U2300 ( .IN1(n3003), .IN2(n3026), .IN3(n2994), .IN4(n3034), .IN5(
        n1381), .IN6(n478), .Q(\fpu_add_frac_dp/n3398 ) );
  AO222X1 U2301 ( .IN1(n3003), .IN2(n3027), .IN3(n2994), .IN4(n3035), .IN5(
        n1381), .IN6(n477), .Q(\fpu_add_frac_dp/n3397 ) );
  AO222X1 U2302 ( .IN1(n3003), .IN2(n3028), .IN3(n2994), .IN4(n3036), .IN5(
        n1382), .IN6(n476), .Q(\fpu_add_frac_dp/n3396 ) );
  AO222X1 U2303 ( .IN1(n3003), .IN2(n3029), .IN3(n2994), .IN4(n3037), .IN5(
        n1382), .IN6(n475), .Q(\fpu_add_frac_dp/n3395 ) );
  AO222X1 U2304 ( .IN1(n3003), .IN2(n3030), .IN3(n2994), .IN4(n3038), .IN5(
        n1382), .IN6(n474), .Q(\fpu_add_frac_dp/n3394 ) );
  AO222X1 U2305 ( .IN1(n3003), .IN2(n3031), .IN3(n2994), .IN4(n3039), .IN5(
        n1382), .IN6(n473), .Q(\fpu_add_frac_dp/n3393 ) );
  AO222X1 U2306 ( .IN1(n3003), .IN2(n3032), .IN3(n2994), .IN4(n3040), .IN5(
        n1382), .IN6(n472), .Q(\fpu_add_frac_dp/n3392 ) );
  AO222X1 U2307 ( .IN1(n3003), .IN2(n3033), .IN3(n2994), .IN4(n3041), .IN5(
        n1382), .IN6(n471), .Q(\fpu_add_frac_dp/n3391 ) );
  AO222X1 U2308 ( .IN1(n3003), .IN2(n3034), .IN3(n2994), .IN4(n3042), .IN5(
        n1382), .IN6(n470), .Q(\fpu_add_frac_dp/n3390 ) );
  AO222X1 U2309 ( .IN1(n3003), .IN2(n3035), .IN3(n2994), .IN4(n3043), .IN5(
        n1382), .IN6(n469), .Q(\fpu_add_frac_dp/n3389 ) );
  AO222X1 U2310 ( .IN1(n3003), .IN2(n3036), .IN3(n3044), .IN4(n2994), .IN5(
        n1382), .IN6(n913), .Q(\fpu_add_frac_dp/n3388 ) );
  AO222X1 U2311 ( .IN1(n3003), .IN2(n3037), .IN3(n3045), .IN4(n2994), .IN5(
        n1382), .IN6(n912), .Q(\fpu_add_frac_dp/n3387 ) );
  AO222X1 U2312 ( .IN1(n3003), .IN2(n3038), .IN3(n3046), .IN4(n2994), .IN5(
        n1382), .IN6(n911), .Q(\fpu_add_frac_dp/n3386 ) );
  AO222X1 U2313 ( .IN1(n3003), .IN2(n3039), .IN3(n2994), .IN4(n3047), .IN5(
        n1382), .IN6(n910), .Q(\fpu_add_frac_dp/n3385 ) );
  AO222X1 U2314 ( .IN1(n3003), .IN2(n3040), .IN3(n3048), .IN4(n2994), .IN5(
        n1383), .IN6(n909), .Q(\fpu_add_frac_dp/n3384 ) );
  AO222X1 U2315 ( .IN1(n3003), .IN2(n3041), .IN3(n3049), .IN4(n2994), .IN5(
        n1383), .IN6(n918), .Q(\fpu_add_frac_dp/n3383 ) );
  AO22X1 U2316 ( .IN1(n1421), .IN2(n1064), .IN3(n1442), .IN4(n3050), .Q(
        \fpu_add_frac_dp/n3382 ) );
  AO221X1 U2317 ( .IN1(n3003), .IN2(n3043), .IN3(n1393), .IN4(n906), .IN5(
        n3051), .Q(\fpu_add_frac_dp/n3381 ) );
  AO22X1 U2318 ( .IN1(n2989), .IN2(n3052), .IN3(n3053), .IN4(n3054), .Q(n3051)
         );
  AO21X1 U2319 ( .IN1(n1404), .IN2(n1034), .IN3(n3055), .Q(
        \fpu_add_frac_dp/n3380 ) );
  AO21X1 U2320 ( .IN1(n1404), .IN2(n933), .IN3(n3056), .Q(
        \fpu_add_frac_dp/n3379 ) );
  AO221X1 U2321 ( .IN1(n3046), .IN2(n3003), .IN3(n1393), .IN4(n466), .IN5(
        n3057), .Q(\fpu_add_frac_dp/n3378 ) );
  AO22X1 U2322 ( .IN1(n3053), .IN2(n3058), .IN3(n2989), .IN4(n3059), .Q(n3057)
         );
  INVX0 U2323 ( .INP(n3060), .ZN(n3059) );
  AO22X1 U2324 ( .IN1(n1421), .IN2(n963), .IN3(n1442), .IN4(n3061), .Q(
        \fpu_add_frac_dp/n3377 ) );
  AO222X1 U2325 ( .IN1(n3048), .IN2(n3003), .IN3(n1435), .IN4(n3062), .IN5(
        n1383), .IN6(n468), .Q(\fpu_add_frac_dp/n3376 ) );
  AO222X1 U2326 ( .IN1(n3049), .IN2(n3003), .IN3(n1435), .IN4(n3063), .IN5(
        n1383), .IN6(n467), .Q(\fpu_add_frac_dp/n3375 ) );
  INVX0 U2327 ( .INP(n3064), .ZN(\fpu_add_frac_dp/n1574 ) );
  AOI222X1 U2328 ( .IN1(\fpu_add_frac_dp/n1569 ), .IN2(n3065), .IN3(n2997), 
        .IN4(n3066), .IN5(n2970), .IN6(n1389), .QN(\fpu_add_frac_dp/n1007 ) );
  AOI222X1 U2329 ( .IN1(n3065), .IN2(\fpu_add_frac_dp/n1568 ), .IN3(n2998), 
        .IN4(\fpu_add_ctl/n319 ), .IN5(n2971), .IN6(n1389), .QN(
        \fpu_add_frac_dp/n1006 ) );
  AO22X1 U2330 ( .IN1(n3008), .IN2(n2994), .IN3(n3001), .IN4(n2988), .Q(n2998)
         );
  INVX0 U2331 ( .INP(n3067), .ZN(\fpu_add_frac_dp/n1568 ) );
  AOI222X1 U2332 ( .IN1(n3065), .IN2(\fpu_add_frac_dp/n1567 ), .IN3(n2999), 
        .IN4(\fpu_add_ctl/n319 ), .IN5(n2972), .IN6(n1389), .QN(
        \fpu_add_frac_dp/n1005 ) );
  AO22X1 U2333 ( .IN1(n3010), .IN2(n2994), .IN3(n3001), .IN4(n2990), .Q(n2999)
         );
  AND2X1 U2334 ( .IN1(n3003), .IN2(\fpu_add_frac_dp/n2471 ), .Q(n3001) );
  INVX0 U2335 ( .INP(n3068), .ZN(\fpu_add_frac_dp/n1567 ) );
  AOI222X1 U2336 ( .IN1(n3065), .IN2(\fpu_add_frac_dp/a3stg_fracadd[0] ), 
        .IN3(n2990), .IN4(n3069), .IN5(n2964), .IN6(n1389), .QN(
        \fpu_add_frac_dp/n1004 ) );
  INVX0 U2337 ( .INP(n3070), .ZN(n2990) );
  OA222X1 U2338 ( .IN1(n3071), .IN2(n3064), .IN3(n3072), .IN4(n3073), .IN5(
        n3074), .IN6(n2046), .Q(\fpu_add_frac_dp/n1003 ) );
  AOI222X1 U2339 ( .IN1(n3065), .IN2(\fpu_add_frac_dp/n1573 ), .IN3(n2992), 
        .IN4(n3069), .IN5(n2966), .IN6(n1389), .QN(\fpu_add_frac_dp/n1002 ) );
  INVX0 U2340 ( .INP(n3075), .ZN(\fpu_add_frac_dp/n1573 ) );
  AOI222X1 U2341 ( .IN1(n3065), .IN2(\fpu_add_frac_dp/n1572 ), .IN3(n2993), 
        .IN4(n3066), .IN5(n2967), .IN6(n1389), .QN(\fpu_add_frac_dp/n1001 ) );
  INVX0 U2342 ( .INP(n3076), .ZN(\fpu_add_frac_dp/n1572 ) );
  NOR2X0 U2343 ( .IN1(n3077), .IN2(n3078), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N9 ) );
  NOR2X0 U2344 ( .IN1(n3077), .IN2(n3079), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N8 ) );
  NOR2X0 U2345 ( .IN1(n3077), .IN2(n3076), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N7 ) );
  XNOR3X1 U2346 ( .IN1(\fpu_add_frac_dp/n732 ), .IN2(\fpu_add_frac_dp/n505 ), 
        .IN3(n3080), .Q(n3076) );
  INVX0 U2347 ( .INP(n3081), .ZN(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N66 )
         );
  NOR2X0 U2348 ( .IN1(n3077), .IN2(n2602), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N65 ) );
  NOR2X0 U2349 ( .IN1(n3077), .IN2(n3082), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N64 ) );
  NOR2X0 U2350 ( .IN1(n3077), .IN2(n3083), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N63 ) );
  NOR2X0 U2351 ( .IN1(n3077), .IN2(n3084), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N62 ) );
  NOR2X0 U2352 ( .IN1(n3077), .IN2(n3085), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N61 ) );
  NOR2X0 U2353 ( .IN1(n3077), .IN2(n3086), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N60 ) );
  NOR2X0 U2354 ( .IN1(n3077), .IN2(n3075), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N6 ) );
  XNOR3X1 U2355 ( .IN1(\fpu_add_frac_dp/n733 ), .IN2(\fpu_add_frac_dp/n504 ), 
        .IN3(n3087), .Q(n3075) );
  NOR2X0 U2356 ( .IN1(n3077), .IN2(n3088), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N59 ) );
  NOR2X0 U2357 ( .IN1(n3077), .IN2(n3089), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N58 ) );
  NOR2X0 U2358 ( .IN1(n3077), .IN2(n3090), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N57 ) );
  NOR2X0 U2359 ( .IN1(n3077), .IN2(n3091), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N56 ) );
  NOR2X0 U2360 ( .IN1(n3077), .IN2(n3092), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N55 ) );
  NOR2X0 U2361 ( .IN1(n3077), .IN2(n3093), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N54 ) );
  NOR2X0 U2362 ( .IN1(n3077), .IN2(n3094), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N53 ) );
  NOR2X0 U2363 ( .IN1(n3077), .IN2(n3095), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N52 ) );
  NOR2X0 U2364 ( .IN1(n3077), .IN2(n3096), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N51 ) );
  NOR2X0 U2365 ( .IN1(n3077), .IN2(n3097), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N50 ) );
  NOR2X0 U2366 ( .IN1(n3077), .IN2(n3064), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N5 ) );
  XNOR3X1 U2367 ( .IN1(\fpu_add_frac_dp/n734 ), .IN2(\fpu_add_frac_dp/n503 ), 
        .IN3(n3098), .Q(n3064) );
  NOR2X0 U2368 ( .IN1(n3077), .IN2(n3099), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N49 ) );
  NOR2X0 U2369 ( .IN1(n3077), .IN2(n3100), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N48 ) );
  NOR2X0 U2370 ( .IN1(n3077), .IN2(n3101), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N47 ) );
  NOR2X0 U2371 ( .IN1(n3077), .IN2(n3102), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N46 ) );
  NOR2X0 U2372 ( .IN1(n3077), .IN2(n3103), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N45 ) );
  NOR2X0 U2373 ( .IN1(n3077), .IN2(n3104), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N44 ) );
  NOR2X0 U2374 ( .IN1(n3077), .IN2(n3105), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N43 ) );
  NOR2X0 U2375 ( .IN1(n3077), .IN2(n3106), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N42 ) );
  NOR2X0 U2376 ( .IN1(n3077), .IN2(n3107), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N41 ) );
  NOR2X0 U2377 ( .IN1(n3077), .IN2(n3108), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N40 ) );
  NOR2X0 U2378 ( .IN1(n3077), .IN2(n3109), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N4 ) );
  INVX0 U2379 ( .INP(\fpu_add_frac_dp/a3stg_fracadd[0] ), .ZN(n3109) );
  NOR2X0 U2380 ( .IN1(n3077), .IN2(n3110), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N39 ) );
  NOR2X0 U2381 ( .IN1(n3077), .IN2(n3111), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N38 ) );
  NOR2X0 U2382 ( .IN1(n3077), .IN2(n3112), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N37 ) );
  NOR2X0 U2383 ( .IN1(n3077), .IN2(n3113), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N36 ) );
  NOR2X0 U2384 ( .IN1(n3077), .IN2(n3114), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N35 ) );
  NOR2X0 U2385 ( .IN1(n3077), .IN2(n3115), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N34 ) );
  NOR2X0 U2386 ( .IN1(n3077), .IN2(n3116), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N33 ) );
  NOR2X0 U2387 ( .IN1(n3077), .IN2(n3117), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N32 ) );
  NOR2X0 U2388 ( .IN1(n3077), .IN2(n3118), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N31 ) );
  NOR2X0 U2389 ( .IN1(n3077), .IN2(n3119), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N30 ) );
  NOR2X0 U2390 ( .IN1(n3077), .IN2(n3120), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N29 ) );
  NOR2X0 U2391 ( .IN1(n3077), .IN2(n3121), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N28 ) );
  NOR2X0 U2392 ( .IN1(n3077), .IN2(n3122), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N27 ) );
  NOR2X0 U2393 ( .IN1(n3077), .IN2(n3123), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N26 ) );
  NOR2X0 U2394 ( .IN1(n3077), .IN2(n3124), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N25 ) );
  NOR2X0 U2395 ( .IN1(n3077), .IN2(n3125), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N24 ) );
  NOR2X0 U2396 ( .IN1(n3077), .IN2(n3126), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N23 ) );
  NOR2X0 U2397 ( .IN1(n3077), .IN2(n3127), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N22 ) );
  NOR2X0 U2398 ( .IN1(n3077), .IN2(n3128), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N21 ) );
  NOR2X0 U2399 ( .IN1(n3077), .IN2(n3129), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N20 ) );
  NOR2X0 U2400 ( .IN1(n3077), .IN2(n3130), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N19 ) );
  NOR2X0 U2401 ( .IN1(n3077), .IN2(n3131), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N18 ) );
  NOR2X0 U2402 ( .IN1(n3077), .IN2(n3132), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N17 ) );
  NOR2X0 U2403 ( .IN1(n3077), .IN2(n3133), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N16 ) );
  NOR2X0 U2404 ( .IN1(n3077), .IN2(n3134), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N15 ) );
  NOR2X0 U2405 ( .IN1(n3077), .IN2(n3135), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N14 ) );
  NOR2X0 U2406 ( .IN1(n3077), .IN2(n3136), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N13 ) );
  NOR2X0 U2407 ( .IN1(n3077), .IN2(n3068), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N12 ) );
  XNOR3X1 U2408 ( .IN1(\fpu_add_frac_dp/n727 ), .IN2(\fpu_add_frac_dp/n502 ), 
        .IN3(n3137), .Q(n3068) );
  NOR2X0 U2409 ( .IN1(n3077), .IN2(n3067), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N11 ) );
  XNOR3X1 U2410 ( .IN1(\fpu_add_frac_dp/n728 ), .IN2(\fpu_add_frac_dp/n501 ), 
        .IN3(n3138), .Q(n3067) );
  NOR2X0 U2411 ( .IN1(n3077), .IN2(n3139), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre3/N10 ) );
  AND2X1 U2412 ( .IN1(n3140), .IN2(n3081), .Q(n3077) );
  NAND4X0 U2413 ( .IN1(n3141), .IN2(n3142), .IN3(n3143), .IN4(n3144), .QN(
        n3081) );
  NAND4X0 U2414 ( .IN1(n2601), .IN2(n583), .IN3(n3142), .IN4(n3145), .QN(n3140) );
  NOR2X0 U2415 ( .IN1(n3146), .IN2(n2602), .QN(n3145) );
  AO221X1 U2416 ( .IN1(\fpu_add_frac_dp/n1569 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(\fpu_add_frac_dp/n1570 ), .IN4(n3065), .IN5(n3147), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N9 ) );
  AO22X1 U2417 ( .IN1(n1421), .IN2(n2969), .IN3(n3066), .IN4(n2996), .Q(n3147)
         );
  INVX0 U2418 ( .INP(n3139), .ZN(\fpu_add_frac_dp/n1569 ) );
  XNOR3X1 U2419 ( .IN1(\fpu_add_frac_dp/n729 ), .IN2(\fpu_add_frac_dp/n507 ), 
        .IN3(n3148), .Q(n3139) );
  AO221X1 U2420 ( .IN1(\fpu_add_frac_dp/n1570 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(\fpu_add_frac_dp/n1571 ), .IN4(n3065), .IN5(n3149), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N8 ) );
  AO22X1 U2421 ( .IN1(n1421), .IN2(n2968), .IN3(n3066), .IN4(n2995), .Q(n3149)
         );
  INVX0 U2422 ( .INP(n3079), .ZN(\fpu_add_frac_dp/n1571 ) );
  XNOR3X1 U2423 ( .IN1(\fpu_add_frac_dp/n731 ), .IN2(\fpu_add_frac_dp/n506 ), 
        .IN3(n3150), .Q(n3079) );
  INVX0 U2424 ( .INP(n3078), .ZN(\fpu_add_frac_dp/n1570 ) );
  XNOR3X1 U2425 ( .IN1(\fpu_add_frac_dp/n730 ), .IN2(\fpu_add_frac_dp/n508 ), 
        .IN3(n3151), .Q(n3078) );
  NAND2X0 U2426 ( .IN1(n3152), .IN2(n3153), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N66 ) );
  OA221X1 U2427 ( .IN1(n3154), .IN2(n3155), .IN3(n3143), .IN4(n3156), .IN5(
        n3157), .Q(n3153) );
  INVX0 U2428 ( .INP(n3063), .ZN(n3154) );
  AO22X1 U2429 ( .IN1(n3158), .IN2(n3159), .IN3(n3160), .IN4(n3161), .Q(n3063)
         );
  OA22X1 U2430 ( .IN1(n3162), .IN2(n3163), .IN3(n3164), .IN4(n3165), .Q(n3161)
         );
  AO21X1 U2431 ( .IN1(n729), .IN2(n2586), .IN3(n3166), .Q(n3163) );
  AO222X1 U2432 ( .IN1(n451), .IN2(n14), .IN3(n846), .IN4(n2591), .IN5(n130), 
        .IN6(n2), .Q(n3162) );
  NOR2X0 U2433 ( .IN1(n3167), .IN2(n3168), .QN(n3160) );
  OA21X1 U2434 ( .IN1(n3169), .IN2(n3170), .IN3(n582), .Q(n3167) );
  OA222X1 U2435 ( .IN1(n3071), .IN2(n3171), .IN3(n3172), .IN4(n3173), .IN5(
        n3174), .IN6(n2046), .Q(n3152) );
  AO221X1 U2436 ( .IN1(n3141), .IN2(\fpu_add_frac_dp/n1509 ), .IN3(n3175), 
        .IN4(n3065), .IN5(n3176), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N65 ) );
  AO222X1 U2437 ( .IN1(n3177), .IN2(n3048), .IN3(n3178), .IN4(n3062), .IN5(
        n1384), .IN6(n2956), .Q(n3176) );
  AO22X1 U2438 ( .IN1(n3158), .IN2(n3179), .IN3(n3180), .IN4(n3181), .Q(n3062)
         );
  OA22X1 U2439 ( .IN1(n3164), .IN2(n3182), .IN3(n3166), .IN4(n3165), .Q(n3181)
         );
  AO221X1 U2440 ( .IN1(n45), .IN2(n2), .IN3(n726), .IN4(n2586), .IN5(n3183), 
        .Q(n3165) );
  AO22X1 U2441 ( .IN1(n456), .IN2(n14), .IN3(n831), .IN4(n2591), .Q(n3183) );
  NOR2X0 U2442 ( .IN1(n3184), .IN2(n3168), .QN(n3180) );
  AOI21X1 U2443 ( .IN1(n3185), .IN2(n3186), .IN3(\fpu_add_frac_dp/n2460 ), 
        .QN(n3184) );
  AO221X1 U2444 ( .IN1(n1389), .IN2(n2952), .IN3(n3175), .IN4(
        \fpu_add_frac_dp/n1509 ), .IN5(n3187), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N64 ) );
  AO22X1 U2445 ( .IN1(\fpu_add_frac_dp/n1515 ), .IN2(n3065), .IN3(n3178), 
        .IN4(n3061), .Q(n3187) );
  AO222X1 U2446 ( .IN1(n3158), .IN2(n3052), .IN3(n3188), .IN4(n3189), .IN5(
        n3047), .IN6(n584), .Q(n3061) );
  MUX21X1 U2447 ( .IN1(n3190), .IN2(n3191), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n3188) );
  NOR2X0 U2448 ( .IN1(n3169), .IN2(n3170), .QN(n3191) );
  NOR2X0 U2449 ( .IN1(n3182), .IN2(n154), .QN(n3170) );
  AO221X1 U2450 ( .IN1(n257), .IN2(n2), .IN3(n727), .IN4(n2586), .IN5(n3192), 
        .Q(n3182) );
  AO22X1 U2451 ( .IN1(n457), .IN2(n14), .IN3(n832), .IN4(n2591), .Q(n3192) );
  AND2X1 U2452 ( .IN1(n3193), .IN2(n154), .Q(n3169) );
  AND2X1 U2453 ( .IN1(n3194), .IN2(n3195), .Q(n3190) );
  INVX0 U2454 ( .INP(n3196), .ZN(n3052) );
  INVX0 U2455 ( .INP(n3082), .ZN(\fpu_add_frac_dp/n1515 ) );
  AO221X1 U2456 ( .IN1(n3197), .IN2(n3046), .IN3(n1392), .IN4(n2948), .IN5(
        n3198), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N63 ) );
  OAI222X1 U2457 ( .IN1(n3199), .IN2(n3082), .IN3(n3200), .IN4(n3155), .IN5(
        n3071), .IN6(n3083), .QN(n3198) );
  OA22X1 U2458 ( .IN1(n3060), .IN2(n3168), .IN3(n3201), .IN4(n3202), .Q(n3200)
         );
  MUX21X1 U2459 ( .IN1(n3203), .IN2(n3204), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n3060) );
  NAND2X0 U2460 ( .IN1(n3186), .IN2(n3185), .QN(n3204) );
  NAND2X0 U2461 ( .IN1(n3205), .IN2(n154), .QN(n3185) );
  NAND2X0 U2462 ( .IN1(n3193), .IN2(\fpu_add_frac_dp/n2449 ), .QN(n3186) );
  AOI221X1 U2463 ( .IN1(n107), .IN2(n2), .IN3(n751), .IN4(n2586), .IN5(n3206), 
        .QN(n3193) );
  AO22X1 U2464 ( .IN1(n464), .IN2(n14), .IN3(n843), .IN4(n2591), .Q(n3206) );
  XNOR3X1 U2465 ( .IN1(\fpu_add_frac_dp/n675 ), .IN2(\fpu_add_frac_dp/n566 ), 
        .IN3(n3207), .Q(n3082) );
  AO221X1 U2466 ( .IN1(\fpu_add_ctl/n319 ), .IN2(n3056), .IN3(
        \fpu_add_frac_dp/n1516 ), .IN4(\fpu_add_frac_dp/n1509 ), .IN5(n3208), 
        .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N62 ) );
  AO22X1 U2467 ( .IN1(n1421), .IN2(n2946), .IN3(\fpu_add_frac_dp/n1517 ), 
        .IN4(n3065), .Q(n3208) );
  INVX0 U2468 ( .INP(n3083), .ZN(\fpu_add_frac_dp/n1516 ) );
  XNOR3X1 U2469 ( .IN1(\fpu_add_frac_dp/n676 ), .IN2(\fpu_add_frac_dp/n565 ), 
        .IN3(n3209), .Q(n3083) );
  AO222X1 U2470 ( .IN1(n2989), .IN2(n3159), .IN3(n3210), .IN4(n3053), .IN5(
        n3045), .IN6(n3003), .Q(n3056) );
  MUX21X1 U2471 ( .IN1(n3211), .IN2(n3212), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n3210) );
  AND2X1 U2472 ( .IN1(n3213), .IN2(n3214), .Q(n3212) );
  INVX0 U2473 ( .INP(n3215), .ZN(n3159) );
  MUX21X1 U2474 ( .IN1(n3216), .IN2(n3217), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n3215) );
  NAND2X0 U2475 ( .IN1(n3195), .IN2(n3194), .QN(n3217) );
  NAND2X0 U2476 ( .IN1(n3218), .IN2(n154), .QN(n3194) );
  NAND2X0 U2477 ( .IN1(n3205), .IN2(\fpu_add_frac_dp/n2449 ), .QN(n3195) );
  AOI221X1 U2478 ( .IN1(n264), .IN2(n2), .IN3(n749), .IN4(n2586), .IN5(n3219), 
        .QN(n3205) );
  AO22X1 U2479 ( .IN1(n461), .IN2(n14), .IN3(n840), .IN4(n2591), .Q(n3219) );
  AO221X1 U2480 ( .IN1(\fpu_add_ctl/n319 ), .IN2(n3055), .IN3(
        \fpu_add_frac_dp/n1517 ), .IN4(\fpu_add_frac_dp/n1509 ), .IN5(n3220), 
        .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N61 ) );
  AO22X1 U2481 ( .IN1(n1422), .IN2(n2942), .IN3(\fpu_add_frac_dp/n1518 ), 
        .IN4(n3065), .Q(n3220) );
  INVX0 U2482 ( .INP(n3085), .ZN(\fpu_add_frac_dp/n1518 ) );
  INVX0 U2483 ( .INP(n3084), .ZN(\fpu_add_frac_dp/n1517 ) );
  XNOR3X1 U2484 ( .IN1(\fpu_add_frac_dp/n677 ), .IN2(\fpu_add_frac_dp/n564 ), 
        .IN3(n3221), .Q(n3084) );
  AO222X1 U2485 ( .IN1(n2989), .IN2(n3179), .IN3(n3222), .IN4(n3053), .IN5(
        n3044), .IN6(n3003), .Q(n3055) );
  NOR2X0 U2486 ( .IN1(n3202), .IN2(n1745), .QN(n3053) );
  MUX21X1 U2487 ( .IN1(n3223), .IN2(n3224), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n3222) );
  AND2X1 U2488 ( .IN1(n3225), .IN2(n3226), .Q(n3224) );
  INVX0 U2489 ( .INP(n3227), .ZN(n3179) );
  MUX21X1 U2490 ( .IN1(n3228), .IN2(n3203), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n3227) );
  NAND2X0 U2491 ( .IN1(n3229), .IN2(n3230), .QN(n3203) );
  NAND2X0 U2492 ( .IN1(n3231), .IN2(n154), .QN(n3230) );
  NAND2X0 U2493 ( .IN1(n3218), .IN2(\fpu_add_frac_dp/n2449 ), .QN(n3229) );
  AOI221X1 U2494 ( .IN1(n766), .IN2(n14), .IN3(n448), .IN4(n2586), .IN5(n3232), 
        .QN(n3218) );
  AO22X1 U2495 ( .IN1(n119), .IN2(n2), .IN3(n833), .IN4(n2591), .Q(n3232) );
  NAND2X0 U2496 ( .IN1(n3233), .IN2(n3234), .QN(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N60 ) );
  OA222X1 U2497 ( .IN1(n3199), .IN2(n3085), .IN3(n3155), .IN4(n3235), .IN5(
        n3196), .IN6(n3073), .Q(n3234) );
  MUX21X1 U2498 ( .IN1(n3236), .IN2(n3216), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n3196) );
  NAND2X0 U2499 ( .IN1(n3237), .IN2(n3238), .QN(n3216) );
  NAND2X0 U2500 ( .IN1(n3239), .IN2(n154), .QN(n3238) );
  NAND2X0 U2501 ( .IN1(n3231), .IN2(\fpu_add_frac_dp/n2449 ), .QN(n3237) );
  AOI221X1 U2502 ( .IN1(n285), .IN2(n2), .IN3(n748), .IN4(n2586), .IN5(n3240), 
        .QN(n3231) );
  AO22X1 U2503 ( .IN1(n462), .IN2(n14), .IN3(n834), .IN4(n2591), .Q(n3240) );
  NAND2X0 U2504 ( .IN1(n3054), .IN2(n3158), .QN(n3235) );
  XNOR3X1 U2505 ( .IN1(\fpu_add_frac_dp/n678 ), .IN2(\fpu_add_frac_dp/n563 ), 
        .IN3(n3241), .Q(n3085) );
  INVX0 U2506 ( .INP(\fpu_add_frac_dp/n1509 ), .ZN(n3199) );
  OA222X1 U2507 ( .IN1(n2939), .IN2(n2046), .IN3(n3071), .IN4(n3086), .IN5(
        n3242), .IN6(n3173), .Q(n3233) );
  INVX0 U2508 ( .INP(n2985), .ZN(n2939) );
  AO221X1 U2509 ( .IN1(n3178), .IN2(n3050), .IN3(\fpu_add_frac_dp/n1519 ), 
        .IN4(\fpu_add_frac_dp/n1509 ), .IN5(n3243), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N59 ) );
  AO22X1 U2510 ( .IN1(n1422), .IN2(n2940), .IN3(\fpu_add_frac_dp/n1520 ), 
        .IN4(n3065), .Q(n3243) );
  INVX0 U2511 ( .INP(n3086), .ZN(\fpu_add_frac_dp/n1519 ) );
  XNOR3X1 U2512 ( .IN1(\fpu_add_frac_dp/n679 ), .IN2(\fpu_add_frac_dp/n562 ), 
        .IN3(n3244), .Q(n3086) );
  AO222X1 U2513 ( .IN1(n3189), .IN2(n3058), .IN3(n3245), .IN4(n3158), .IN5(
        n3042), .IN6(n584), .Q(n3050) );
  INVX0 U2514 ( .INP(n3202), .ZN(n3158) );
  NAND2X0 U2515 ( .IN1(\fpu_add_frac_dp/n2307 ), .IN2(n63), .QN(n3202) );
  MUX21X1 U2516 ( .IN1(n3246), .IN2(n3223), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n3245) );
  INVX0 U2517 ( .INP(n3201), .ZN(n3058) );
  MUX21X1 U2518 ( .IN1(n3247), .IN2(n3228), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n3201) );
  NAND2X0 U2519 ( .IN1(n3248), .IN2(n3249), .QN(n3228) );
  NAND2X0 U2520 ( .IN1(n3250), .IN2(n154), .QN(n3249) );
  NAND2X0 U2521 ( .IN1(n3239), .IN2(\fpu_add_frac_dp/n2449 ), .QN(n3248) );
  AOI221X1 U2522 ( .IN1(n123), .IN2(n2), .IN3(n752), .IN4(n2586), .IN5(n3251), 
        .QN(n3239) );
  AO22X1 U2523 ( .IN1(n458), .IN2(n14), .IN3(n844), .IN4(n2591), .Q(n3251) );
  INVX0 U2524 ( .INP(n3168), .ZN(n3189) );
  INVX0 U2525 ( .INP(n3155), .ZN(n3178) );
  AO221X1 U2526 ( .IN1(n3177), .IN2(n3041), .IN3(n1392), .IN4(n2932), .IN5(
        n3252), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N58 ) );
  AO222X1 U2527 ( .IN1(\fpu_add_frac_dp/n1520 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3049), .IN5(\fpu_add_frac_dp/n1521 ), .IN6(n3065), 
        .Q(n3252) );
  INVX0 U2528 ( .INP(n3172), .ZN(n3049) );
  AO221X1 U2529 ( .IN1(n3253), .IN2(n3254), .IN3(n3255), .IN4(n3256), .IN5(
        n3257), .Q(n3172) );
  AO22X1 U2530 ( .IN1(n3258), .IN2(n3259), .IN3(n3260), .IN4(n3236), .Q(n3257)
         );
  NAND2X0 U2531 ( .IN1(n3214), .IN2(n3213), .QN(n3236) );
  NAND2X0 U2532 ( .IN1(n3261), .IN2(n154), .QN(n3213) );
  NAND2X0 U2533 ( .IN1(n3250), .IN2(\fpu_add_frac_dp/n2449 ), .QN(n3214) );
  AOI221X1 U2534 ( .IN1(n286), .IN2(n2), .IN3(n750), .IN4(n2586), .IN5(n3262), 
        .QN(n3250) );
  AO22X1 U2535 ( .IN1(n459), .IN2(n14), .IN3(n841), .IN4(n2591), .Q(n3262) );
  OR2X1 U2536 ( .IN1(n3263), .IN2(n3264), .Q(n3256) );
  INVX0 U2537 ( .INP(n3088), .ZN(\fpu_add_frac_dp/n1520 ) );
  XNOR3X1 U2538 ( .IN1(\fpu_add_frac_dp/n680 ), .IN2(\fpu_add_frac_dp/n561 ), 
        .IN3(n3265), .Q(n3088) );
  AO221X1 U2539 ( .IN1(n3177), .IN2(n3040), .IN3(n1393), .IN4(n2928), .IN5(
        n3266), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N57 ) );
  AO222X1 U2540 ( .IN1(\fpu_add_frac_dp/n1521 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3048), .IN5(\fpu_add_frac_dp/n1522 ), .IN6(n3065), 
        .Q(n3266) );
  AOI221X1 U2541 ( .IN1(n3253), .IN2(n3267), .IN3(n3255), .IN4(n3268), .IN5(
        n3269), .QN(n3048) );
  AO22X1 U2542 ( .IN1(n3258), .IN2(n3270), .IN3(n3260), .IN4(n3247), .Q(n3269)
         );
  NAND2X0 U2543 ( .IN1(n3226), .IN2(n3225), .QN(n3247) );
  NAND2X0 U2544 ( .IN1(n3271), .IN2(n154), .QN(n3225) );
  NAND2X0 U2545 ( .IN1(n3261), .IN2(\fpu_add_frac_dp/n2449 ), .QN(n3226) );
  AOI221X1 U2546 ( .IN1(n767), .IN2(n14), .IN3(n449), .IN4(n2586), .IN5(n3272), 
        .QN(n3261) );
  AO22X1 U2547 ( .IN1(n124), .IN2(n2), .IN3(n835), .IN4(n2591), .Q(n3272) );
  INVX0 U2548 ( .INP(n3089), .ZN(\fpu_add_frac_dp/n1521 ) );
  XNOR3X1 U2549 ( .IN1(\fpu_add_frac_dp/n681 ), .IN2(\fpu_add_frac_dp/n560 ), 
        .IN3(n3273), .Q(n3089) );
  AO221X1 U2550 ( .IN1(n3197), .IN2(n3039), .IN3(n1392), .IN4(n2926), .IN5(
        n3274), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N56 ) );
  AO222X1 U2551 ( .IN1(\fpu_add_frac_dp/n1522 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3275), .IN4(n3047), .IN5(\fpu_add_frac_dp/n1523 ), .IN6(n3065), 
        .Q(n3274) );
  MUX21X1 U2552 ( .IN1(n3054), .IN2(n3276), .S(n63), .Q(n3047) );
  INVX0 U2553 ( .INP(n3277), .ZN(n3276) );
  MUX21X1 U2554 ( .IN1(n3278), .IN2(n3211), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n3054) );
  NOR2X0 U2555 ( .IN1(n3264), .IN2(n3263), .QN(n3211) );
  AND2X1 U2556 ( .IN1(n3271), .IN2(\fpu_add_frac_dp/n2449 ), .Q(n3263) );
  AOI221X1 U2557 ( .IN1(n765), .IN2(n14), .IN3(n450), .IN4(n2586), .IN5(n3279), 
        .QN(n3271) );
  AO22X1 U2558 ( .IN1(n51), .IN2(n2), .IN3(n836), .IN4(n2591), .Q(n3279) );
  NOR2X0 U2559 ( .IN1(n3280), .IN2(\fpu_add_frac_dp/n2449 ), .QN(n3264) );
  INVX0 U2560 ( .INP(n3090), .ZN(\fpu_add_frac_dp/n1522 ) );
  XNOR3X1 U2561 ( .IN1(\fpu_add_frac_dp/n682 ), .IN2(\fpu_add_frac_dp/n559 ), 
        .IN3(n3281), .Q(n3090) );
  AO221X1 U2562 ( .IN1(n3177), .IN2(n3038), .IN3(n1392), .IN4(n2922), .IN5(
        n3282), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N55 ) );
  AO222X1 U2563 ( .IN1(\fpu_add_frac_dp/n1523 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3046), .IN5(\fpu_add_frac_dp/n1524 ), .IN6(n3065), 
        .Q(n3282) );
  AOI222X1 U2564 ( .IN1(n3255), .IN2(n3270), .IN3(n63), .IN4(n3283), .IN5(
        n3260), .IN6(n3268), .QN(n3046) );
  INVX0 U2565 ( .INP(n3223), .ZN(n3268) );
  MUX21X1 U2566 ( .IN1(n3284), .IN2(n3280), .S(\fpu_add_frac_dp/n2449 ), .Q(
        n3223) );
  AO221X1 U2567 ( .IN1(n742), .IN2(n14), .IN3(n432), .IN4(n2586), .IN5(n3285), 
        .Q(n3280) );
  AO22X1 U2568 ( .IN1(n284), .IN2(n2), .IN3(n845), .IN4(n2591), .Q(n3285) );
  INVX0 U2569 ( .INP(n3091), .ZN(\fpu_add_frac_dp/n1523 ) );
  XNOR3X1 U2570 ( .IN1(\fpu_add_frac_dp/n683 ), .IN2(\fpu_add_frac_dp/n558 ), 
        .IN3(n3286), .Q(n3091) );
  AO221X1 U2571 ( .IN1(n3177), .IN2(n3037), .IN3(n1392), .IN4(n2920), .IN5(
        n3287), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N54 ) );
  AO222X1 U2572 ( .IN1(\fpu_add_frac_dp/n1524 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3045), .IN5(\fpu_add_frac_dp/n1525 ), .IN6(n3065), 
        .Q(n3287) );
  AOI222X1 U2573 ( .IN1(n3255), .IN2(n3254), .IN3(n63), .IN4(n3288), .IN5(
        n3260), .IN6(n3259), .QN(n3045) );
  INVX0 U2574 ( .INP(n3278), .ZN(n3259) );
  MUX21X1 U2575 ( .IN1(n3289), .IN2(n3284), .S(\fpu_add_frac_dp/n2449 ), .Q(
        n3278) );
  AO221X1 U2576 ( .IN1(n741), .IN2(n14), .IN3(n431), .IN4(n2586), .IN5(n3290), 
        .Q(n3284) );
  AO22X1 U2577 ( .IN1(n50), .IN2(n2), .IN3(n842), .IN4(n2591), .Q(n3290) );
  INVX0 U2578 ( .INP(n3092), .ZN(\fpu_add_frac_dp/n1524 ) );
  XNOR3X1 U2579 ( .IN1(\fpu_add_frac_dp/n684 ), .IN2(\fpu_add_frac_dp/n557 ), 
        .IN3(n3291), .Q(n3092) );
  AO221X1 U2580 ( .IN1(n3177), .IN2(n3036), .IN3(n1393), .IN4(n2916), .IN5(
        n3292), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N53 ) );
  AO222X1 U2581 ( .IN1(\fpu_add_frac_dp/n1525 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3044), .IN5(\fpu_add_frac_dp/n1526 ), .IN6(n3065), 
        .Q(n3292) );
  AOI222X1 U2582 ( .IN1(n3255), .IN2(n3267), .IN3(n63), .IN4(n3293), .IN5(
        n3260), .IN6(n3270), .QN(n3044) );
  INVX0 U2583 ( .INP(n3246), .ZN(n3270) );
  MUX21X1 U2584 ( .IN1(n3294), .IN2(n3289), .S(\fpu_add_frac_dp/n2449 ), .Q(
        n3246) );
  AO221X1 U2585 ( .IN1(n739), .IN2(n14), .IN3(n429), .IN4(n2586), .IN5(n3295), 
        .Q(n3289) );
  AO22X1 U2586 ( .IN1(n115), .IN2(n2), .IN3(n837), .IN4(n2591), .Q(n3295) );
  INVX0 U2587 ( .INP(n3093), .ZN(\fpu_add_frac_dp/n1525 ) );
  XNOR3X1 U2588 ( .IN1(\fpu_add_frac_dp/n685 ), .IN2(\fpu_add_frac_dp/n556 ), 
        .IN3(n3296), .Q(n3093) );
  AO221X1 U2589 ( .IN1(n3177), .IN2(n3035), .IN3(n1392), .IN4(n2914), .IN5(
        n3297), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N52 ) );
  AO222X1 U2590 ( .IN1(\fpu_add_frac_dp/n1526 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3043), .IN5(\fpu_add_frac_dp/n1527 ), .IN6(n3065), 
        .Q(n3297) );
  INVX0 U2591 ( .INP(n3242), .ZN(n3043) );
  MUX21X1 U2592 ( .IN1(n3298), .IN2(n3277), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3242) );
  AO222X1 U2593 ( .IN1(n3299), .IN2(n3300), .IN3(\fpu_add_frac_dp/n2460 ), 
        .IN4(n3254), .IN5(n3301), .IN6(n3302), .Q(n3277) );
  INVX0 U2594 ( .INP(n3303), .ZN(n3254) );
  MUX21X1 U2595 ( .IN1(n3304), .IN2(n3294), .S(\fpu_add_frac_dp/n2449 ), .Q(
        n3303) );
  AO221X1 U2596 ( .IN1(n740), .IN2(n14), .IN3(n430), .IN4(n2586), .IN5(n3305), 
        .Q(n3294) );
  AO22X1 U2597 ( .IN1(n48), .IN2(n2), .IN3(n838), .IN4(n2591), .Q(n3305) );
  NAND3X0 U2598 ( .IN1(n3306), .IN2(n3307), .IN3(n3308), .QN(n3304) );
  INVX0 U2599 ( .INP(n3094), .ZN(\fpu_add_frac_dp/n1526 ) );
  XNOR3X1 U2600 ( .IN1(\fpu_add_frac_dp/n686 ), .IN2(\fpu_add_frac_dp/n555 ), 
        .IN3(n3309), .Q(n3094) );
  AO221X1 U2601 ( .IN1(n3177), .IN2(n3034), .IN3(n1393), .IN4(n2910), .IN5(
        n3310), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N51 ) );
  AO222X1 U2602 ( .IN1(\fpu_add_frac_dp/n1527 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3042), .IN5(\fpu_add_frac_dp/n1528 ), .IN6(n3065), 
        .Q(n3310) );
  INVX0 U2603 ( .INP(n3311), .ZN(n3042) );
  MUX21X1 U2604 ( .IN1(n3312), .IN2(n3283), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3311) );
  AO222X1 U2605 ( .IN1(n3301), .IN2(n3300), .IN3(\fpu_add_frac_dp/n2460 ), 
        .IN4(n3267), .IN5(n3313), .IN6(n3302), .Q(n3283) );
  MUX21X1 U2606 ( .IN1(n3314), .IN2(n3299), .S(n154), .Q(n3267) );
  AND3X1 U2607 ( .IN1(n3306), .IN2(n3307), .IN3(n3308), .Q(n3314) );
  OA22X1 U2608 ( .IN1(\fpu_add_frac_dp/n592 ), .IN2(\fpu_add_frac_dp/n2401 ), 
        .IN3(\fpu_add_frac_dp/n5633 ), .IN4(\fpu_add_frac_dp/n250 ), .Q(n3308)
         );
  NAND2X0 U2609 ( .IN1(n2591), .IN2(n914), .QN(n3307) );
  INVX0 U2610 ( .INP(\fpu_add_frac_dp/n5634 ), .ZN(n2591) );
  NAND2X0 U2611 ( .IN1(n2586), .IN2(n756), .QN(n3306) );
  INVX0 U2612 ( .INP(\fpu_add_frac_dp/n5635 ), .ZN(n2586) );
  INVX0 U2613 ( .INP(n3095), .ZN(\fpu_add_frac_dp/n1527 ) );
  XNOR3X1 U2614 ( .IN1(\fpu_add_frac_dp/n687 ), .IN2(\fpu_add_frac_dp/n554 ), 
        .IN3(n3315), .Q(n3095) );
  AO221X1 U2615 ( .IN1(n3177), .IN2(n3033), .IN3(n1392), .IN4(n2908), .IN5(
        n3316), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N50 ) );
  AO222X1 U2616 ( .IN1(\fpu_add_frac_dp/n1528 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3041), .IN5(\fpu_add_frac_dp/n1529 ), .IN6(n3065), 
        .Q(n3316) );
  INVX0 U2617 ( .INP(n3317), .ZN(n3041) );
  MUX21X1 U2618 ( .IN1(n3318), .IN2(n3288), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3317) );
  AO221X1 U2619 ( .IN1(n3313), .IN2(n3300), .IN3(n3319), .IN4(n3302), .IN5(
        n3320), .Q(n3288) );
  AO22X1 U2620 ( .IN1(n3301), .IN2(n3321), .IN3(n3299), .IN4(n3322), .Q(n3320)
         );
  OA222X1 U2621 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n220 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2417 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n252 ), .Q(n3299) );
  INVX0 U2622 ( .INP(n3096), .ZN(\fpu_add_frac_dp/n1528 ) );
  XNOR3X1 U2623 ( .IN1(\fpu_add_frac_dp/n688 ), .IN2(\fpu_add_frac_dp/n553 ), 
        .IN3(n3323), .Q(n3096) );
  AO221X1 U2624 ( .IN1(n3177), .IN2(n3032), .IN3(n1392), .IN4(n2904), .IN5(
        n3324), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N49 ) );
  AO222X1 U2625 ( .IN1(\fpu_add_frac_dp/n1529 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3040), .IN5(\fpu_add_frac_dp/n1530 ), .IN6(n3065), 
        .Q(n3324) );
  INVX0 U2626 ( .INP(n3325), .ZN(n3040) );
  MUX21X1 U2627 ( .IN1(n3326), .IN2(n3293), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3325) );
  AO221X1 U2628 ( .IN1(n3319), .IN2(n3300), .IN3(n3327), .IN4(n3302), .IN5(
        n3328), .Q(n3293) );
  AO22X1 U2629 ( .IN1(n3313), .IN2(n3321), .IN3(n3301), .IN4(n3322), .Q(n3328)
         );
  OA222X1 U2630 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n222 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2291 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n254 ), .Q(n3301) );
  INVX0 U2631 ( .INP(n3097), .ZN(\fpu_add_frac_dp/n1529 ) );
  XNOR3X1 U2632 ( .IN1(\fpu_add_frac_dp/n689 ), .IN2(\fpu_add_frac_dp/n552 ), 
        .IN3(n3329), .Q(n3097) );
  AO221X1 U2633 ( .IN1(n3177), .IN2(n3031), .IN3(n1391), .IN4(n2902), .IN5(
        n3330), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N48 ) );
  AO222X1 U2634 ( .IN1(\fpu_add_frac_dp/n1530 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3039), .IN5(\fpu_add_frac_dp/n1531 ), .IN6(n3065), 
        .Q(n3330) );
  INVX0 U2635 ( .INP(n3331), .ZN(n3039) );
  MUX21X1 U2636 ( .IN1(n3332), .IN2(n3298), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3331) );
  AO221X1 U2637 ( .IN1(n3327), .IN2(n3300), .IN3(n3333), .IN4(n3302), .IN5(
        n3334), .Q(n3298) );
  AO22X1 U2638 ( .IN1(n3319), .IN2(n3321), .IN3(n3313), .IN4(n3322), .Q(n3334)
         );
  OA222X1 U2639 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n224 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2358 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n256 ), .Q(n3313) );
  INVX0 U2640 ( .INP(n3099), .ZN(\fpu_add_frac_dp/n1530 ) );
  XNOR3X1 U2641 ( .IN1(\fpu_add_frac_dp/n690 ), .IN2(\fpu_add_frac_dp/n551 ), 
        .IN3(n3335), .Q(n3099) );
  AO221X1 U2642 ( .IN1(n3177), .IN2(n3030), .IN3(n1394), .IN4(n2898), .IN5(
        n3336), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N47 ) );
  AO222X1 U2643 ( .IN1(\fpu_add_frac_dp/n1531 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3038), .IN5(\fpu_add_frac_dp/n1532 ), .IN6(n3065), 
        .Q(n3336) );
  INVX0 U2644 ( .INP(n3337), .ZN(n3038) );
  MUX21X1 U2645 ( .IN1(n3338), .IN2(n3312), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3337) );
  AO221X1 U2646 ( .IN1(n3333), .IN2(n3300), .IN3(n3339), .IN4(n3302), .IN5(
        n3340), .Q(n3312) );
  AO22X1 U2647 ( .IN1(n3327), .IN2(n3321), .IN3(n3319), .IN4(n3322), .Q(n3340)
         );
  OA222X1 U2648 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n226 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2292 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n258 ), .Q(n3319) );
  INVX0 U2649 ( .INP(n3100), .ZN(\fpu_add_frac_dp/n1531 ) );
  XNOR3X1 U2650 ( .IN1(\fpu_add_frac_dp/n691 ), .IN2(\fpu_add_frac_dp/n550 ), 
        .IN3(n3341), .Q(n3100) );
  AO221X1 U2651 ( .IN1(n3177), .IN2(n3029), .IN3(n1391), .IN4(n2896), .IN5(
        n3342), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N46 ) );
  AO222X1 U2652 ( .IN1(\fpu_add_frac_dp/n1532 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3037), .IN5(\fpu_add_frac_dp/n1533 ), .IN6(n3065), 
        .Q(n3342) );
  INVX0 U2653 ( .INP(n3343), .ZN(n3037) );
  MUX21X1 U2654 ( .IN1(n3344), .IN2(n3318), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3343) );
  AO221X1 U2655 ( .IN1(n3339), .IN2(n3300), .IN3(n3345), .IN4(n3302), .IN5(
        n3346), .Q(n3318) );
  AO22X1 U2656 ( .IN1(n3333), .IN2(n3321), .IN3(n3327), .IN4(n3322), .Q(n3346)
         );
  OA222X1 U2657 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n228 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2360 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n260 ), .Q(n3327) );
  INVX0 U2658 ( .INP(n3101), .ZN(\fpu_add_frac_dp/n1532 ) );
  XNOR3X1 U2659 ( .IN1(\fpu_add_frac_dp/n692 ), .IN2(\fpu_add_frac_dp/n549 ), 
        .IN3(n3347), .Q(n3101) );
  AO221X1 U2660 ( .IN1(n3197), .IN2(n3028), .IN3(n1391), .IN4(n2891), .IN5(
        n3348), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N45 ) );
  AO222X1 U2661 ( .IN1(\fpu_add_frac_dp/n1533 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3275), .IN4(n3036), .IN5(\fpu_add_frac_dp/n1534 ), .IN6(n3065), 
        .Q(n3348) );
  INVX0 U2662 ( .INP(n3349), .ZN(n3036) );
  MUX21X1 U2663 ( .IN1(n3350), .IN2(n3326), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3349) );
  AO221X1 U2664 ( .IN1(n3345), .IN2(n3300), .IN3(n3351), .IN4(n3302), .IN5(
        n3352), .Q(n3326) );
  AO22X1 U2665 ( .IN1(n3339), .IN2(n3321), .IN3(n3333), .IN4(n3322), .Q(n3352)
         );
  OA222X1 U2666 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n230 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2293 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n262 ), .Q(n3333) );
  INVX0 U2667 ( .INP(n3102), .ZN(\fpu_add_frac_dp/n1533 ) );
  XNOR3X1 U2668 ( .IN1(\fpu_add_frac_dp/n693 ), .IN2(\fpu_add_frac_dp/n548 ), 
        .IN3(n3353), .Q(n3102) );
  AO221X1 U2669 ( .IN1(n3177), .IN2(n3027), .IN3(n1392), .IN4(n2888), .IN5(
        n3354), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N44 ) );
  AO222X1 U2670 ( .IN1(\fpu_add_frac_dp/n1534 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3035), .IN5(\fpu_add_frac_dp/n1535 ), .IN6(n3065), 
        .Q(n3354) );
  INVX0 U2671 ( .INP(n3355), .ZN(n3035) );
  MUX21X1 U2672 ( .IN1(n3356), .IN2(n3332), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3355) );
  AO221X1 U2673 ( .IN1(n3351), .IN2(n3300), .IN3(n3357), .IN4(n3302), .IN5(
        n3358), .Q(n3332) );
  AO22X1 U2674 ( .IN1(n3345), .IN2(n3321), .IN3(n3339), .IN4(n3322), .Q(n3358)
         );
  OA222X1 U2675 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n232 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2410 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n264 ), .Q(n3339) );
  INVX0 U2676 ( .INP(n3103), .ZN(\fpu_add_frac_dp/n1534 ) );
  XNOR3X1 U2677 ( .IN1(\fpu_add_frac_dp/n694 ), .IN2(\fpu_add_frac_dp/n547 ), 
        .IN3(n3359), .Q(n3103) );
  AO221X1 U2678 ( .IN1(n3177), .IN2(n3026), .IN3(n1391), .IN4(n2984), .IN5(
        n3360), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N43 ) );
  AO222X1 U2679 ( .IN1(\fpu_add_frac_dp/n1535 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3034), .IN5(\fpu_add_frac_dp/n1536 ), .IN6(n3065), 
        .Q(n3360) );
  INVX0 U2680 ( .INP(n3361), .ZN(n3034) );
  MUX21X1 U2681 ( .IN1(n3362), .IN2(n3338), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3361) );
  AO221X1 U2682 ( .IN1(n3357), .IN2(n3300), .IN3(n3363), .IN4(n3302), .IN5(
        n3364), .Q(n3338) );
  AO22X1 U2683 ( .IN1(n3351), .IN2(n3321), .IN3(n3345), .IN4(n3322), .Q(n3364)
         );
  OA222X1 U2684 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n234 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2346 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n266 ), .Q(n3345) );
  INVX0 U2685 ( .INP(n3104), .ZN(\fpu_add_frac_dp/n1535 ) );
  XNOR3X1 U2686 ( .IN1(\fpu_add_frac_dp/n695 ), .IN2(\fpu_add_frac_dp/n546 ), 
        .IN3(n3365), .Q(n3104) );
  AO221X1 U2687 ( .IN1(n3177), .IN2(n3025), .IN3(n1391), .IN4(n2983), .IN5(
        n3366), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N42 ) );
  AO222X1 U2688 ( .IN1(\fpu_add_frac_dp/n1536 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3033), .IN5(\fpu_add_frac_dp/n1537 ), .IN6(n3065), 
        .Q(n3366) );
  INVX0 U2689 ( .INP(n3367), .ZN(n3033) );
  MUX21X1 U2690 ( .IN1(n3368), .IN2(n3344), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3367) );
  AO221X1 U2691 ( .IN1(n3363), .IN2(n3300), .IN3(n3369), .IN4(n3302), .IN5(
        n3370), .Q(n3344) );
  AO22X1 U2692 ( .IN1(n3357), .IN2(n3321), .IN3(n3351), .IN4(n3322), .Q(n3370)
         );
  OA222X1 U2693 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n236 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2413 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n268 ), .Q(n3351) );
  INVX0 U2694 ( .INP(n3105), .ZN(\fpu_add_frac_dp/n1536 ) );
  XNOR3X1 U2695 ( .IN1(\fpu_add_frac_dp/n696 ), .IN2(\fpu_add_frac_dp/n544 ), 
        .IN3(n3371), .Q(n3105) );
  AO221X1 U2696 ( .IN1(n3177), .IN2(n3024), .IN3(n1391), .IN4(n2881), .IN5(
        n3372), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N41 ) );
  AO222X1 U2697 ( .IN1(\fpu_add_frac_dp/n1537 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3032), .IN5(\fpu_add_frac_dp/n1538 ), .IN6(n3065), 
        .Q(n3372) );
  INVX0 U2698 ( .INP(n3373), .ZN(n3032) );
  MUX21X1 U2699 ( .IN1(n3374), .IN2(n3350), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3373) );
  AO221X1 U2700 ( .IN1(n3369), .IN2(n3300), .IN3(n3375), .IN4(n3302), .IN5(
        n3376), .Q(n3350) );
  AO22X1 U2701 ( .IN1(n3363), .IN2(n3321), .IN3(n3357), .IN4(n3322), .Q(n3376)
         );
  OA222X1 U2702 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n238 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2349 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n270 ), .Q(n3357) );
  INVX0 U2703 ( .INP(n3106), .ZN(\fpu_add_frac_dp/n1537 ) );
  XNOR3X1 U2704 ( .IN1(\fpu_add_frac_dp/n697 ), .IN2(\fpu_add_frac_dp/n543 ), 
        .IN3(n3377), .Q(n3106) );
  AO221X1 U2705 ( .IN1(n3177), .IN2(n3023), .IN3(n1391), .IN4(n2982), .IN5(
        n3378), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N40 ) );
  AO222X1 U2706 ( .IN1(\fpu_add_frac_dp/n1538 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3031), .IN5(\fpu_add_frac_dp/n1539 ), .IN6(n3065), 
        .Q(n3378) );
  INVX0 U2707 ( .INP(n3379), .ZN(n3031) );
  MUX21X1 U2708 ( .IN1(n3380), .IN2(n3356), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3379) );
  AO221X1 U2709 ( .IN1(n3375), .IN2(n3300), .IN3(n3381), .IN4(n3302), .IN5(
        n3382), .Q(n3356) );
  AO22X1 U2710 ( .IN1(n3369), .IN2(n3321), .IN3(n3363), .IN4(n3322), .Q(n3382)
         );
  OA222X1 U2711 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n240 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2294 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n272 ), .Q(n3363) );
  INVX0 U2712 ( .INP(n3107), .ZN(\fpu_add_frac_dp/n1538 ) );
  XNOR3X1 U2713 ( .IN1(\fpu_add_frac_dp/n698 ), .IN2(\fpu_add_frac_dp/n542 ), 
        .IN3(n3383), .Q(n3107) );
  AO221X1 U2714 ( .IN1(n3177), .IN2(n3022), .IN3(n1391), .IN4(n2867), .IN5(
        n3384), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N39 ) );
  AO222X1 U2715 ( .IN1(\fpu_add_frac_dp/n1539 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3030), .IN5(\fpu_add_frac_dp/n1540 ), .IN6(n3065), 
        .Q(n3384) );
  INVX0 U2716 ( .INP(n3385), .ZN(n3030) );
  MUX21X1 U2717 ( .IN1(n3386), .IN2(n3362), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3385) );
  AO221X1 U2718 ( .IN1(n3381), .IN2(n3300), .IN3(n3387), .IN4(n3302), .IN5(
        n3388), .Q(n3362) );
  AO22X1 U2719 ( .IN1(n3375), .IN2(n3321), .IN3(n3369), .IN4(n3322), .Q(n3388)
         );
  OA222X1 U2720 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n242 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2414 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n274 ), .Q(n3369) );
  INVX0 U2721 ( .INP(n3108), .ZN(\fpu_add_frac_dp/n1539 ) );
  XNOR3X1 U2722 ( .IN1(\fpu_add_frac_dp/n699 ), .IN2(\fpu_add_frac_dp/n541 ), 
        .IN3(n3389), .Q(n3108) );
  AO221X1 U2723 ( .IN1(n3177), .IN2(n3021), .IN3(n1392), .IN4(n2981), .IN5(
        n3390), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N38 ) );
  AO222X1 U2724 ( .IN1(\fpu_add_frac_dp/n1540 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3029), .IN5(\fpu_add_frac_dp/n1541 ), .IN6(n3065), 
        .Q(n3390) );
  INVX0 U2725 ( .INP(n3391), .ZN(n3029) );
  MUX21X1 U2726 ( .IN1(n3392), .IN2(n3368), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3391) );
  AO221X1 U2727 ( .IN1(n3387), .IN2(n3300), .IN3(n3393), .IN4(n3302), .IN5(
        n3394), .Q(n3368) );
  AO22X1 U2728 ( .IN1(n3381), .IN2(n3321), .IN3(n3375), .IN4(n3322), .Q(n3394)
         );
  OA222X1 U2729 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n244 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2347 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n276 ), .Q(n3375) );
  INVX0 U2730 ( .INP(n3110), .ZN(\fpu_add_frac_dp/n1540 ) );
  XNOR3X1 U2731 ( .IN1(\fpu_add_frac_dp/n700 ), .IN2(\fpu_add_frac_dp/n540 ), 
        .IN3(n3395), .Q(n3110) );
  AO221X1 U2732 ( .IN1(n3177), .IN2(n3020), .IN3(n1391), .IN4(n2980), .IN5(
        n3396), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N37 ) );
  AO222X1 U2733 ( .IN1(\fpu_add_frac_dp/n1541 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3028), .IN5(\fpu_add_frac_dp/n1542 ), .IN6(n3065), 
        .Q(n3396) );
  INVX0 U2734 ( .INP(n3397), .ZN(n3028) );
  MUX21X1 U2735 ( .IN1(n3398), .IN2(n3374), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3397) );
  AO221X1 U2736 ( .IN1(n3393), .IN2(n3300), .IN3(n3399), .IN4(n3302), .IN5(
        n3400), .Q(n3374) );
  AO22X1 U2737 ( .IN1(n3387), .IN2(n3321), .IN3(n3381), .IN4(n3322), .Q(n3400)
         );
  OA222X1 U2738 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n246 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2412 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n278 ), .Q(n3381) );
  INVX0 U2739 ( .INP(n3111), .ZN(\fpu_add_frac_dp/n1541 ) );
  XNOR3X1 U2740 ( .IN1(\fpu_add_frac_dp/n701 ), .IN2(\fpu_add_frac_dp/n539 ), 
        .IN3(n3401), .Q(n3111) );
  AO221X1 U2741 ( .IN1(n3177), .IN2(n3019), .IN3(n1391), .IN4(n2858), .IN5(
        n3402), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N36 ) );
  AO222X1 U2742 ( .IN1(\fpu_add_frac_dp/n1542 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3027), .IN5(\fpu_add_frac_dp/n1543 ), .IN6(n3065), 
        .Q(n3402) );
  INVX0 U2743 ( .INP(n3403), .ZN(n3027) );
  MUX21X1 U2744 ( .IN1(n3404), .IN2(n3380), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3403) );
  AO221X1 U2745 ( .IN1(n3399), .IN2(n3300), .IN3(n3405), .IN4(n3302), .IN5(
        n3406), .Q(n3380) );
  AO22X1 U2746 ( .IN1(n3393), .IN2(n3321), .IN3(n3387), .IN4(n3322), .Q(n3406)
         );
  OA222X1 U2747 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n248 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2348 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n280 ), .Q(n3387) );
  INVX0 U2748 ( .INP(n3112), .ZN(\fpu_add_frac_dp/n1542 ) );
  XNOR3X1 U2749 ( .IN1(\fpu_add_frac_dp/n702 ), .IN2(\fpu_add_frac_dp/n538 ), 
        .IN3(n3407), .Q(n3112) );
  AO221X1 U2750 ( .IN1(n3177), .IN2(n3018), .IN3(n1391), .IN4(n2854), .IN5(
        n3408), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N35 ) );
  AO222X1 U2751 ( .IN1(\fpu_add_frac_dp/n1543 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3026), .IN5(\fpu_add_frac_dp/n1544 ), .IN6(n3065), 
        .Q(n3408) );
  INVX0 U2752 ( .INP(n3409), .ZN(n3026) );
  MUX21X1 U2753 ( .IN1(n3410), .IN2(n3386), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3409) );
  AO221X1 U2754 ( .IN1(n3405), .IN2(n3300), .IN3(n3411), .IN4(n3302), .IN5(
        n3412), .Q(n3386) );
  AO22X1 U2755 ( .IN1(n3399), .IN2(n3321), .IN3(n3393), .IN4(n3322), .Q(n3412)
         );
  OA222X1 U2756 ( .IN1(\fpu_add_frac_dp/n5634 ), .IN2(\fpu_add_frac_dp/n250 ), 
        .IN3(\fpu_add_frac_dp/n5635 ), .IN4(\fpu_add_frac_dp/n2401 ), .IN5(
        \fpu_add_frac_dp/n5633 ), .IN6(\fpu_add_frac_dp/n282 ), .Q(n3393) );
  INVX0 U2757 ( .INP(n3113), .ZN(\fpu_add_frac_dp/n1543 ) );
  XNOR3X1 U2758 ( .IN1(\fpu_add_frac_dp/n703 ), .IN2(\fpu_add_frac_dp/n537 ), 
        .IN3(n3413), .Q(n3113) );
  AO221X1 U2759 ( .IN1(n3177), .IN2(n3017), .IN3(n1391), .IN4(n2852), .IN5(
        n3414), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N34 ) );
  AO222X1 U2760 ( .IN1(\fpu_add_frac_dp/n1544 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3025), .IN5(\fpu_add_frac_dp/n1545 ), .IN6(n3065), 
        .Q(n3414) );
  INVX0 U2761 ( .INP(n3415), .ZN(n3025) );
  MUX21X1 U2762 ( .IN1(n3416), .IN2(n3392), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3415) );
  AO221X1 U2763 ( .IN1(n3411), .IN2(n3300), .IN3(n3417), .IN4(n3302), .IN5(
        n3418), .Q(n3392) );
  AO22X1 U2764 ( .IN1(n3405), .IN2(n3321), .IN3(n3399), .IN4(n3322), .Q(n3418)
         );
  OA22X1 U2765 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2417 ), 
        .IN3(\fpu_add_frac_dp/n252 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3399)
         );
  INVX0 U2766 ( .INP(n3114), .ZN(\fpu_add_frac_dp/n1544 ) );
  XNOR3X1 U2767 ( .IN1(\fpu_add_frac_dp/n704 ), .IN2(\fpu_add_frac_dp/n536 ), 
        .IN3(n3419), .Q(n3114) );
  AO221X1 U2768 ( .IN1(n3177), .IN2(n3016), .IN3(n1390), .IN4(n2848), .IN5(
        n3420), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N33 ) );
  AO222X1 U2769 ( .IN1(\fpu_add_frac_dp/n1545 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3024), .IN5(\fpu_add_frac_dp/n1546 ), .IN6(n3065), 
        .Q(n3420) );
  INVX0 U2770 ( .INP(n3421), .ZN(n3024) );
  MUX21X1 U2771 ( .IN1(n3422), .IN2(n3398), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3421) );
  AO221X1 U2772 ( .IN1(n3417), .IN2(n3300), .IN3(n3423), .IN4(n3302), .IN5(
        n3424), .Q(n3398) );
  AO22X1 U2773 ( .IN1(n3411), .IN2(n3321), .IN3(n3405), .IN4(n3322), .Q(n3424)
         );
  OA22X1 U2774 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2291 ), 
        .IN3(\fpu_add_frac_dp/n254 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3405)
         );
  INVX0 U2775 ( .INP(n3115), .ZN(\fpu_add_frac_dp/n1545 ) );
  XNOR3X1 U2776 ( .IN1(\fpu_add_frac_dp/n705 ), .IN2(\fpu_add_frac_dp/n535 ), 
        .IN3(n3425), .Q(n3115) );
  AO221X1 U2777 ( .IN1(n3197), .IN2(n3015), .IN3(n1391), .IN4(n2846), .IN5(
        n3426), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N32 ) );
  AO222X1 U2778 ( .IN1(\fpu_add_frac_dp/n1546 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3275), .IN4(n3023), .IN5(\fpu_add_frac_dp/n1547 ), .IN6(n3065), 
        .Q(n3426) );
  INVX0 U2779 ( .INP(n3427), .ZN(n3023) );
  MUX21X1 U2780 ( .IN1(n3428), .IN2(n3404), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3427) );
  AO221X1 U2781 ( .IN1(n3423), .IN2(n3300), .IN3(n3429), .IN4(n3302), .IN5(
        n3430), .Q(n3404) );
  AO22X1 U2782 ( .IN1(n3417), .IN2(n3321), .IN3(n3411), .IN4(n3322), .Q(n3430)
         );
  OA22X1 U2783 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2358 ), 
        .IN3(\fpu_add_frac_dp/n256 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3411)
         );
  INVX0 U2784 ( .INP(n3116), .ZN(\fpu_add_frac_dp/n1546 ) );
  XNOR3X1 U2785 ( .IN1(\fpu_add_frac_dp/n706 ), .IN2(\fpu_add_frac_dp/n534 ), 
        .IN3(n3431), .Q(n3116) );
  AO221X1 U2786 ( .IN1(n3177), .IN2(n3014), .IN3(n1390), .IN4(n2842), .IN5(
        n3432), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N31 ) );
  AO222X1 U2787 ( .IN1(\fpu_add_frac_dp/n1547 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3022), .IN5(\fpu_add_frac_dp/n1548 ), .IN6(n3065), 
        .Q(n3432) );
  INVX0 U2788 ( .INP(n3433), .ZN(n3022) );
  MUX21X1 U2789 ( .IN1(n3434), .IN2(n3410), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3433) );
  AO221X1 U2790 ( .IN1(n3429), .IN2(n3300), .IN3(n3435), .IN4(n3302), .IN5(
        n3436), .Q(n3410) );
  AO22X1 U2791 ( .IN1(n3423), .IN2(n3321), .IN3(n3417), .IN4(n3322), .Q(n3436)
         );
  OA22X1 U2792 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2292 ), 
        .IN3(\fpu_add_frac_dp/n258 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3417)
         );
  INVX0 U2793 ( .INP(n3117), .ZN(\fpu_add_frac_dp/n1547 ) );
  XNOR3X1 U2794 ( .IN1(\fpu_add_frac_dp/n707 ), .IN2(\fpu_add_frac_dp/n533 ), 
        .IN3(n3437), .Q(n3117) );
  AO221X1 U2795 ( .IN1(n3197), .IN2(n3013), .IN3(n1390), .IN4(n2840), .IN5(
        n3438), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N30 ) );
  AO222X1 U2796 ( .IN1(\fpu_add_frac_dp/n1548 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3275), .IN4(n3021), .IN5(\fpu_add_frac_dp/n1549 ), .IN6(n3065), 
        .Q(n3438) );
  INVX0 U2797 ( .INP(n3439), .ZN(n3021) );
  MUX21X1 U2798 ( .IN1(n3440), .IN2(n3416), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3439) );
  AO221X1 U2799 ( .IN1(n3435), .IN2(n3300), .IN3(n3441), .IN4(n3302), .IN5(
        n3442), .Q(n3416) );
  AO22X1 U2800 ( .IN1(n3429), .IN2(n3321), .IN3(n3423), .IN4(n3322), .Q(n3442)
         );
  OA22X1 U2801 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2360 ), 
        .IN3(\fpu_add_frac_dp/n260 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3423)
         );
  INVX0 U2802 ( .INP(n3118), .ZN(\fpu_add_frac_dp/n1548 ) );
  XNOR3X1 U2803 ( .IN1(\fpu_add_frac_dp/n708 ), .IN2(\fpu_add_frac_dp/n532 ), 
        .IN3(n3443), .Q(n3118) );
  AO222X1 U2804 ( .IN1(n1415), .IN2(n956), .IN3(n3069), .IN4(n2988), .IN5(
        \fpu_add_frac_dp/a3stg_fracadd[0] ), .IN6(\fpu_add_frac_dp/n1509 ), 
        .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N3 ) );
  INVX0 U2805 ( .INP(n3444), .ZN(n2988) );
  INVX0 U2806 ( .INP(n3073), .ZN(n3069) );
  NAND2X0 U2807 ( .IN1(\fpu_add_ctl/n319 ), .IN2(n2989), .QN(n3073) );
  NOR2X0 U2808 ( .IN1(n3168), .IN2(n1745), .QN(n2989) );
  NAND2X0 U2809 ( .IN1(\fpu_add_frac_dp/n2471 ), .IN2(\fpu_add_frac_dp/n2307 ), 
        .QN(n3168) );
  AO221X1 U2810 ( .IN1(n3177), .IN2(n3012), .IN3(n1390), .IN4(n2836), .IN5(
        n3445), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N29 ) );
  AO222X1 U2811 ( .IN1(\fpu_add_frac_dp/n1549 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3020), .IN5(\fpu_add_frac_dp/n1550 ), .IN6(n3065), 
        .Q(n3445) );
  INVX0 U2812 ( .INP(n3446), .ZN(n3020) );
  MUX21X1 U2813 ( .IN1(n3447), .IN2(n3422), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3446) );
  AO221X1 U2814 ( .IN1(n3441), .IN2(n3300), .IN3(n3448), .IN4(n3302), .IN5(
        n3449), .Q(n3422) );
  AO22X1 U2815 ( .IN1(n3435), .IN2(n3321), .IN3(n3429), .IN4(n3322), .Q(n3449)
         );
  OA22X1 U2816 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2293 ), 
        .IN3(\fpu_add_frac_dp/n262 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3429)
         );
  INVX0 U2817 ( .INP(n3119), .ZN(\fpu_add_frac_dp/n1549 ) );
  XNOR3X1 U2818 ( .IN1(\fpu_add_frac_dp/n709 ), .IN2(\fpu_add_frac_dp/n531 ), 
        .IN3(n3450), .Q(n3119) );
  AO221X1 U2819 ( .IN1(n3177), .IN2(n3011), .IN3(n1390), .IN4(n2834), .IN5(
        n3451), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N28 ) );
  AO222X1 U2820 ( .IN1(\fpu_add_frac_dp/n1550 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3019), .IN5(\fpu_add_frac_dp/n1551 ), .IN6(n3065), 
        .Q(n3451) );
  INVX0 U2821 ( .INP(n3452), .ZN(n3019) );
  MUX21X1 U2822 ( .IN1(n3453), .IN2(n3428), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3452) );
  AO221X1 U2823 ( .IN1(n3448), .IN2(n3300), .IN3(n3454), .IN4(n3302), .IN5(
        n3455), .Q(n3428) );
  AO22X1 U2824 ( .IN1(n3441), .IN2(n3321), .IN3(n3435), .IN4(n3322), .Q(n3455)
         );
  OA22X1 U2825 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2410 ), 
        .IN3(\fpu_add_frac_dp/n264 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3435)
         );
  INVX0 U2826 ( .INP(n3120), .ZN(\fpu_add_frac_dp/n1550 ) );
  XNOR3X1 U2827 ( .IN1(\fpu_add_frac_dp/n710 ), .IN2(\fpu_add_frac_dp/n530 ), 
        .IN3(n3456), .Q(n3120) );
  AO221X1 U2828 ( .IN1(n3177), .IN2(n3009), .IN3(n1391), .IN4(n2830), .IN5(
        n3457), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N27 ) );
  AO222X1 U2829 ( .IN1(\fpu_add_frac_dp/n1551 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3018), .IN5(\fpu_add_frac_dp/n1552 ), .IN6(n3065), 
        .Q(n3457) );
  INVX0 U2830 ( .INP(n3458), .ZN(n3018) );
  MUX21X1 U2831 ( .IN1(n3459), .IN2(n3434), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3458) );
  AO221X1 U2832 ( .IN1(n3454), .IN2(n3300), .IN3(n3460), .IN4(n3302), .IN5(
        n3461), .Q(n3434) );
  AO22X1 U2833 ( .IN1(n3448), .IN2(n3321), .IN3(n3441), .IN4(n3322), .Q(n3461)
         );
  OA22X1 U2834 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2346 ), 
        .IN3(\fpu_add_frac_dp/n266 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3441)
         );
  INVX0 U2835 ( .INP(n3121), .ZN(\fpu_add_frac_dp/n1551 ) );
  XNOR3X1 U2836 ( .IN1(\fpu_add_frac_dp/n711 ), .IN2(\fpu_add_frac_dp/n529 ), 
        .IN3(n3462), .Q(n3121) );
  AO221X1 U2837 ( .IN1(n3177), .IN2(n3007), .IN3(n1390), .IN4(n2979), .IN5(
        n3463), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N26 ) );
  AO222X1 U2838 ( .IN1(\fpu_add_frac_dp/n1552 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3017), .IN5(\fpu_add_frac_dp/n1553 ), .IN6(n3065), 
        .Q(n3463) );
  INVX0 U2839 ( .INP(n3464), .ZN(n3017) );
  MUX21X1 U2840 ( .IN1(n3465), .IN2(n3440), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3464) );
  AO221X1 U2841 ( .IN1(n3460), .IN2(n3300), .IN3(n3466), .IN4(n3302), .IN5(
        n3467), .Q(n3440) );
  AO22X1 U2842 ( .IN1(n3454), .IN2(n3321), .IN3(n3448), .IN4(n3322), .Q(n3467)
         );
  OA22X1 U2843 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2413 ), 
        .IN3(\fpu_add_frac_dp/n268 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3448)
         );
  INVX0 U2844 ( .INP(n3122), .ZN(\fpu_add_frac_dp/n1552 ) );
  XNOR3X1 U2845 ( .IN1(\fpu_add_frac_dp/n712 ), .IN2(\fpu_add_frac_dp/n527 ), 
        .IN3(n3468), .Q(n3122) );
  AO221X1 U2846 ( .IN1(n3177), .IN2(n3006), .IN3(n1392), .IN4(n2978), .IN5(
        n3469), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N25 ) );
  AO222X1 U2847 ( .IN1(\fpu_add_frac_dp/n1553 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3016), .IN5(\fpu_add_frac_dp/n1554 ), .IN6(n3065), 
        .Q(n3469) );
  INVX0 U2848 ( .INP(n3470), .ZN(n3016) );
  MUX21X1 U2849 ( .IN1(n3471), .IN2(n3447), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3470) );
  AO221X1 U2850 ( .IN1(n3466), .IN2(n3300), .IN3(n3472), .IN4(n3302), .IN5(
        n3473), .Q(n3447) );
  AO22X1 U2851 ( .IN1(n3460), .IN2(n3321), .IN3(n3454), .IN4(n3322), .Q(n3473)
         );
  OA22X1 U2852 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2349 ), 
        .IN3(\fpu_add_frac_dp/n270 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3454)
         );
  INVX0 U2853 ( .INP(n3123), .ZN(\fpu_add_frac_dp/n1553 ) );
  XNOR3X1 U2854 ( .IN1(\fpu_add_frac_dp/n713 ), .IN2(\fpu_add_frac_dp/n526 ), 
        .IN3(n3474), .Q(n3123) );
  AO221X1 U2855 ( .IN1(n3177), .IN2(n3005), .IN3(n1390), .IN4(n2977), .IN5(
        n3475), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N24 ) );
  AO222X1 U2856 ( .IN1(\fpu_add_frac_dp/n1554 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3015), .IN5(\fpu_add_frac_dp/n1555 ), .IN6(n3065), 
        .Q(n3475) );
  INVX0 U2857 ( .INP(n3476), .ZN(n3015) );
  MUX21X1 U2858 ( .IN1(n3477), .IN2(n3453), .S(\fpu_add_frac_dp/n2471 ), .Q(
        n3476) );
  AO221X1 U2859 ( .IN1(n3302), .IN2(n3478), .IN3(n3472), .IN4(n3300), .IN5(
        n3479), .Q(n3453) );
  AO22X1 U2860 ( .IN1(n3466), .IN2(n3321), .IN3(n3460), .IN4(n3322), .Q(n3479)
         );
  OA22X1 U2861 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2294 ), 
        .IN3(\fpu_add_frac_dp/n272 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3460)
         );
  INVX0 U2862 ( .INP(n3124), .ZN(\fpu_add_frac_dp/n1554 ) );
  XNOR3X1 U2863 ( .IN1(\fpu_add_frac_dp/n714 ), .IN2(\fpu_add_frac_dp/n525 ), 
        .IN3(n3480), .Q(n3124) );
  AO221X1 U2864 ( .IN1(n3197), .IN2(n3004), .IN3(n1390), .IN4(n2815), .IN5(
        n3481), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N23 ) );
  AO222X1 U2865 ( .IN1(\fpu_add_frac_dp/n1555 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3275), .IN4(n3014), .IN5(\fpu_add_frac_dp/n1556 ), .IN6(n3065), 
        .Q(n3481) );
  AOI222X1 U2866 ( .IN1(n3253), .IN2(n3482), .IN3(\fpu_add_frac_dp/n2471 ), 
        .IN4(n3459), .IN5(n3483), .IN6(n3258), .QN(n3014) );
  AO221X1 U2867 ( .IN1(n3466), .IN2(n3322), .IN3(n3302), .IN4(n3484), .IN5(
        n3485), .Q(n3459) );
  AO22X1 U2868 ( .IN1(n3472), .IN2(n3321), .IN3(n3300), .IN4(n3478), .Q(n3485)
         );
  OA22X1 U2869 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2414 ), 
        .IN3(\fpu_add_frac_dp/n274 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3466)
         );
  INVX0 U2870 ( .INP(n3125), .ZN(\fpu_add_frac_dp/n1555 ) );
  XNOR3X1 U2871 ( .IN1(\fpu_add_frac_dp/n715 ), .IN2(\fpu_add_frac_dp/n524 ), 
        .IN3(n3486), .Q(n3125) );
  AO221X1 U2872 ( .IN1(n3177), .IN2(n3002), .IN3(n1390), .IN4(n2976), .IN5(
        n3487), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N22 ) );
  AO222X1 U2873 ( .IN1(\fpu_add_frac_dp/n1556 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3013), .IN5(\fpu_add_frac_dp/n1557 ), .IN6(n3065), 
        .Q(n3487) );
  AOI222X1 U2874 ( .IN1(n3488), .IN2(n3253), .IN3(\fpu_add_frac_dp/n2471 ), 
        .IN4(n3465), .IN5(n3489), .IN6(n3258), .QN(n3013) );
  AO221X1 U2875 ( .IN1(n3302), .IN2(n3490), .IN3(n3300), .IN4(n3484), .IN5(
        n3491), .Q(n3465) );
  AO22X1 U2876 ( .IN1(n3478), .IN2(n3321), .IN3(n3472), .IN4(n3322), .Q(n3491)
         );
  OA22X1 U2877 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2347 ), 
        .IN3(\fpu_add_frac_dp/n276 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3472)
         );
  NOR2X0 U2878 ( .IN1(n154), .IN2(\fpu_add_frac_dp/n2460 ), .QN(n3300) );
  NOR2X0 U2879 ( .IN1(\fpu_add_frac_dp/n2449 ), .IN2(\fpu_add_frac_dp/n2460 ), 
        .QN(n3302) );
  INVX0 U2880 ( .INP(n3126), .ZN(\fpu_add_frac_dp/n1556 ) );
  XNOR3X1 U2881 ( .IN1(\fpu_add_frac_dp/n716 ), .IN2(\fpu_add_frac_dp/n523 ), 
        .IN3(n3492), .Q(n3126) );
  AO221X1 U2882 ( .IN1(n3177), .IN2(n3000), .IN3(n1390), .IN4(n2975), .IN5(
        n3493), .Q(\fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N21 ) );
  AO222X1 U2883 ( .IN1(\fpu_add_frac_dp/n1557 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(n3066), .IN4(n3012), .IN5(\fpu_add_frac_dp/n1558 ), .IN6(n3065), 
        .Q(n3493) );
  AOI222X1 U2884 ( .IN1(n3253), .IN2(n3494), .IN3(\fpu_add_frac_dp/n2471 ), 
        .IN4(n3471), .IN5(n3258), .IN6(n3482), .QN(n3012) );
  AO222X1 U2885 ( .IN1(n3321), .IN2(n3484), .IN3(n3478), .IN4(n3322), .IN5(
        n3483), .IN6(n582), .Q(n3471) );
  OA22X1 U2886 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2412 ), 
        .IN3(\fpu_add_frac_dp/n278 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3478)
         );
  INVX0 U2887 ( .INP(n3127), .ZN(\fpu_add_frac_dp/n1557 ) );
  XNOR3X1 U2888 ( .IN1(\fpu_add_frac_dp/n717 ), .IN2(\fpu_add_frac_dp/n522 ), 
        .IN3(n3495), .Q(n3127) );
  AO221X1 U2889 ( .IN1(\fpu_add_frac_dp/n1559 ), .IN2(n3065), .IN3(n1389), 
        .IN4(n2974), .IN5(n3496), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N20 ) );
  AO222X1 U2890 ( .IN1(n3177), .IN2(n3010), .IN3(n3066), .IN4(n3011), .IN5(
        \fpu_add_frac_dp/n1558 ), .IN6(\fpu_add_frac_dp/n1509 ), .Q(n3496) );
  INVX0 U2891 ( .INP(n3128), .ZN(\fpu_add_frac_dp/n1558 ) );
  XNOR3X1 U2892 ( .IN1(\fpu_add_frac_dp/n718 ), .IN2(\fpu_add_frac_dp/n521 ), 
        .IN3(n3497), .Q(n3128) );
  AOI222X1 U2893 ( .IN1(n3498), .IN2(n3253), .IN3(\fpu_add_frac_dp/n2471 ), 
        .IN4(n3477), .IN5(n3488), .IN6(n3258), .QN(n3011) );
  AO222X1 U2894 ( .IN1(n3490), .IN2(n3321), .IN3(n3484), .IN4(n3322), .IN5(
        n3489), .IN6(n582), .Q(n3477) );
  INVX0 U2895 ( .INP(n3166), .ZN(n3322) );
  NAND2X0 U2896 ( .IN1(\fpu_add_frac_dp/n2460 ), .IN2(\fpu_add_frac_dp/n2449 ), 
        .QN(n3166) );
  OA22X1 U2897 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2348 ), 
        .IN3(\fpu_add_frac_dp/n280 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3484)
         );
  INVX0 U2898 ( .INP(n3164), .ZN(n3321) );
  NAND2X0 U2899 ( .IN1(\fpu_add_frac_dp/n2460 ), .IN2(n154), .QN(n3164) );
  AOI221X1 U2900 ( .IN1(n3253), .IN2(n3499), .IN3(n3500), .IN4(n3255), .IN5(
        n3501), .QN(n3010) );
  AO22X1 U2901 ( .IN1(n3258), .IN2(n3502), .IN3(n3503), .IN4(n3260), .Q(n3501)
         );
  AO221X1 U2902 ( .IN1(\fpu_add_frac_dp/n1560 ), .IN2(n3065), .IN3(n1390), 
        .IN4(n2800), .IN5(n3504), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N19 ) );
  AO222X1 U2903 ( .IN1(n3177), .IN2(n3008), .IN3(n3066), .IN4(n3009), .IN5(
        \fpu_add_frac_dp/n1559 ), .IN6(\fpu_add_frac_dp/n1509 ), .Q(n3504) );
  INVX0 U2904 ( .INP(n3129), .ZN(\fpu_add_frac_dp/n1559 ) );
  XNOR3X1 U2905 ( .IN1(\fpu_add_frac_dp/n719 ), .IN2(\fpu_add_frac_dp/n520 ), 
        .IN3(n3505), .Q(n3129) );
  AOI221X1 U2906 ( .IN1(n3483), .IN2(n3260), .IN3(n3258), .IN4(n3494), .IN5(
        n3506), .QN(n3009) );
  AO22X1 U2907 ( .IN1(n3507), .IN2(n3253), .IN3(n3255), .IN4(n3482), .Q(n3506)
         );
  OA22X1 U2908 ( .IN1(n154), .IN2(n3490), .IN3(n3508), .IN4(
        \fpu_add_frac_dp/n2417 ), .Q(n3483) );
  OA22X1 U2909 ( .IN1(\fpu_add_frac_dp/n589 ), .IN2(\fpu_add_frac_dp/n2401 ), 
        .IN3(\fpu_add_frac_dp/n282 ), .IN4(\fpu_add_frac_dp/n2271 ), .Q(n3490)
         );
  AOI221X1 U2910 ( .IN1(n3253), .IN2(n3509), .IN3(n3510), .IN4(n3255), .IN5(
        n3511), .QN(n3008) );
  AO22X1 U2911 ( .IN1(n3512), .IN2(n3260), .IN3(n3258), .IN4(n3513), .Q(n3511)
         );
  AO221X1 U2912 ( .IN1(\fpu_add_frac_dp/n1561 ), .IN2(n3065), .IN3(n1389), 
        .IN4(n2798), .IN5(n3514), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N18 ) );
  AO222X1 U2913 ( .IN1(n3177), .IN2(n2997), .IN3(n3066), .IN4(n3007), .IN5(
        \fpu_add_frac_dp/n1560 ), .IN6(\fpu_add_frac_dp/n1509 ), .Q(n3514) );
  INVX0 U2914 ( .INP(n3130), .ZN(\fpu_add_frac_dp/n1560 ) );
  XNOR3X1 U2915 ( .IN1(\fpu_add_frac_dp/n720 ), .IN2(\fpu_add_frac_dp/n519 ), 
        .IN3(n3515), .Q(n3130) );
  AOI221X1 U2916 ( .IN1(n3503), .IN2(n3253), .IN3(n3488), .IN4(n3255), .IN5(
        n3516), .QN(n3007) );
  AO22X1 U2917 ( .IN1(n3498), .IN2(n3258), .IN3(n3489), .IN4(n3260), .Q(n3516)
         );
  AOI22X1 U2918 ( .IN1(n3517), .IN2(n130), .IN3(n3518), .IN4(n45), .QN(n3489)
         );
  AOI222X1 U2919 ( .IN1(n3502), .IN2(n3255), .IN3(n3519), .IN4(n63), .IN5(
        n3500), .IN6(n3260), .QN(n2997) );
  AO221X1 U2920 ( .IN1(\fpu_add_frac_dp/n1562 ), .IN2(n3065), .IN3(n1390), 
        .IN4(n2794), .IN5(n3520), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N17 ) );
  AO222X1 U2921 ( .IN1(n3197), .IN2(n2996), .IN3(n3275), .IN4(n3006), .IN5(
        \fpu_add_frac_dp/n1561 ), .IN6(\fpu_add_frac_dp/n1509 ), .Q(n3520) );
  INVX0 U2922 ( .INP(n3131), .ZN(\fpu_add_frac_dp/n1561 ) );
  XNOR3X1 U2923 ( .IN1(\fpu_add_frac_dp/n721 ), .IN2(\fpu_add_frac_dp/n518 ), 
        .IN3(n3521), .Q(n3131) );
  AOI221X1 U2924 ( .IN1(n3253), .IN2(n3512), .IN3(n3255), .IN4(n3494), .IN5(
        n3522), .QN(n3006) );
  AO22X1 U2925 ( .IN1(n3507), .IN2(n3258), .IN3(n3260), .IN4(n3482), .Q(n3522)
         );
  NAND2X0 U2926 ( .IN1(n3523), .IN2(n596), .QN(n3482) );
  MUX21X1 U2927 ( .IN1(n257), .IN2(n45), .S(\fpu_add_frac_dp/n2449 ), .Q(n3523) );
  AOI222X1 U2928 ( .IN1(n3255), .IN2(n3513), .IN3(n3072), .IN4(n63), .IN5(
        n3510), .IN6(n3260), .QN(n2996) );
  AO221X1 U2929 ( .IN1(\fpu_add_frac_dp/n1563 ), .IN2(n3065), .IN3(n1389), 
        .IN4(n2792), .IN5(n3524), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N16 ) );
  AO222X1 U2930 ( .IN1(n3177), .IN2(n2995), .IN3(n3066), .IN4(n3005), .IN5(
        \fpu_add_frac_dp/n1562 ), .IN6(\fpu_add_frac_dp/n1509 ), .Q(n3524) );
  INVX0 U2931 ( .INP(n3132), .ZN(\fpu_add_frac_dp/n1562 ) );
  XNOR3X1 U2932 ( .IN1(\fpu_add_frac_dp/n722 ), .IN2(\fpu_add_frac_dp/n517 ), 
        .IN3(n3525), .Q(n3132) );
  AOI221X1 U2933 ( .IN1(n3253), .IN2(n3500), .IN3(n3498), .IN4(n3255), .IN5(
        n3526), .QN(n3005) );
  AO22X1 U2934 ( .IN1(n3503), .IN2(n3258), .IN3(n3488), .IN4(n3260), .Q(n3526)
         );
  AOI22X1 U2935 ( .IN1(n3517), .IN2(n257), .IN3(n3518), .IN4(n107), .QN(n3488)
         );
  INVX0 U2936 ( .INP(n3508), .ZN(n3518) );
  NAND2X0 U2937 ( .IN1(n154), .IN2(n596), .QN(n3508) );
  AOI222X1 U2938 ( .IN1(n3255), .IN2(n3499), .IN3(n63), .IN4(n3070), .IN5(
        n3502), .IN6(n3260), .QN(n2995) );
  NAND2X0 U2939 ( .IN1(\fpu_add_frac_dp/n2460 ), .IN2(n3527), .QN(n3070) );
  INVX0 U2940 ( .INP(n3528), .ZN(n3499) );
  AO221X1 U2941 ( .IN1(\fpu_add_frac_dp/n1564 ), .IN2(n3065), .IN3(n1390), 
        .IN4(n2788), .IN5(n3529), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N15 ) );
  AO222X1 U2942 ( .IN1(n3177), .IN2(n2993), .IN3(n3066), .IN4(n3004), .IN5(
        \fpu_add_frac_dp/n1563 ), .IN6(\fpu_add_frac_dp/n1509 ), .Q(n3529) );
  INVX0 U2943 ( .INP(n3133), .ZN(\fpu_add_frac_dp/n1563 ) );
  XNOR3X1 U2944 ( .IN1(\fpu_add_frac_dp/n723 ), .IN2(\fpu_add_frac_dp/n516 ), 
        .IN3(n3530), .Q(n3133) );
  AOI221X1 U2945 ( .IN1(n3253), .IN2(n3510), .IN3(n3507), .IN4(n3255), .IN5(
        n3531), .QN(n3004) );
  AO22X1 U2946 ( .IN1(n3512), .IN2(n3258), .IN3(n3260), .IN4(n3494), .Q(n3531)
         );
  NAND2X0 U2947 ( .IN1(n3532), .IN2(n596), .QN(n3494) );
  MUX21X1 U2948 ( .IN1(n264), .IN2(n107), .S(\fpu_add_frac_dp/n2449 ), .Q(
        n3532) );
  AND2X1 U2949 ( .IN1(\fpu_add_ctl/n319 ), .IN2(n2994), .Q(n3066) );
  AOI222X1 U2950 ( .IN1(n3513), .IN2(n3260), .IN3(n63), .IN4(n3444), .IN5(
        n3255), .IN6(n3509), .QN(n2993) );
  INVX0 U2951 ( .INP(n3533), .ZN(n3509) );
  NAND3X0 U2952 ( .IN1(n3534), .IN2(n219), .IN3(\fpu_add_frac_dp/n2460 ), .QN(
        n3444) );
  INVX0 U2953 ( .INP(n3173), .ZN(n3177) );
  NAND2X0 U2954 ( .IN1(\fpu_add_ctl/n319 ), .IN2(n3003), .QN(n3173) );
  NOR2X0 U2955 ( .IN1(n1745), .IN2(\fpu_add_frac_dp/n2307 ), .QN(n3003) );
  AO221X1 U2956 ( .IN1(n1389), .IN2(n2786), .IN3(\fpu_add_frac_dp/n1565 ), 
        .IN4(n3065), .IN5(n3535), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N14 ) );
  AO222X1 U2957 ( .IN1(n3275), .IN2(n3002), .IN3(n3536), .IN4(n3197), .IN5(
        \fpu_add_frac_dp/n1564 ), .IN6(\fpu_add_frac_dp/n1509 ), .Q(n3535) );
  INVX0 U2958 ( .INP(n3134), .ZN(\fpu_add_frac_dp/n1564 ) );
  XNOR3X1 U2959 ( .IN1(\fpu_add_frac_dp/n724 ), .IN2(\fpu_add_frac_dp/n514 ), 
        .IN3(n3537), .Q(n3134) );
  NOR2X0 U2960 ( .IN1(n63), .IN2(n3519), .QN(n3536) );
  INVX0 U2961 ( .INP(n2992), .ZN(n3519) );
  MUX21X1 U2962 ( .IN1(n3527), .IN2(n3528), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n2992) );
  AO22X1 U2963 ( .IN1(n3538), .IN2(n115), .IN3(n3534), .IN4(n50), .Q(n3528) );
  AO22X1 U2964 ( .IN1(n3538), .IN2(n219), .IN3(n3534), .IN4(n48), .Q(n3527) );
  AOI221X1 U2965 ( .IN1(n3253), .IN2(n3502), .IN3(n3503), .IN4(n3255), .IN5(
        n3539), .QN(n3002) );
  AO22X1 U2966 ( .IN1(n3498), .IN2(n3260), .IN3(n3258), .IN4(n3500), .Q(n3539)
         );
  AOI22X1 U2967 ( .IN1(n3534), .IN2(n286), .IN3(n3538), .IN4(n124), .QN(n3500)
         );
  AOI22X1 U2968 ( .IN1(n3517), .IN2(n264), .IN3(n3538), .IN4(n119), .QN(n3498)
         );
  NOR2X0 U2969 ( .IN1(n154), .IN2(\fpu_add_frac_dp/n2271 ), .QN(n3517) );
  AOI22X1 U2970 ( .IN1(n3534), .IN2(n285), .IN3(n3538), .IN4(n123), .QN(n3503)
         );
  AOI22X1 U2971 ( .IN1(n3538), .IN2(n284), .IN3(n3534), .IN4(n51), .QN(n3502)
         );
  AO221X1 U2972 ( .IN1(\fpu_add_frac_dp/n1565 ), .IN2(\fpu_add_frac_dp/n1509 ), 
        .IN3(\fpu_add_frac_dp/n1566 ), .IN4(n3065), .IN5(n3540), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre2/N13 ) );
  AO222X1 U2973 ( .IN1(n1415), .IN2(n2973), .IN3(n3541), .IN4(n3197), .IN5(
        n3275), .IN6(n3000), .Q(n3540) );
  AOI221X1 U2974 ( .IN1(n3253), .IN2(n3513), .IN3(n3512), .IN4(n3255), .IN5(
        n3542), .QN(n3000) );
  AO22X1 U2975 ( .IN1(n3507), .IN2(n3260), .IN3(n3258), .IN4(n3510), .Q(n3542)
         );
  AOI22X1 U2976 ( .IN1(n3534), .IN2(n124), .IN3(n3538), .IN4(n51), .QN(n3510)
         );
  NOR2X0 U2977 ( .IN1(n582), .IN2(\fpu_add_frac_dp/n2471 ), .QN(n3258) );
  NOR2X0 U2978 ( .IN1(n63), .IN2(n582), .QN(n3260) );
  AOI22X1 U2979 ( .IN1(n3538), .IN2(n285), .IN3(n3534), .IN4(n119), .QN(n3507)
         );
  NOR2X0 U2980 ( .IN1(n63), .IN2(\fpu_add_frac_dp/n2460 ), .QN(n3255) );
  AOI22X1 U2981 ( .IN1(n3538), .IN2(n286), .IN3(n3534), .IN4(n123), .QN(n3512)
         );
  AOI22X1 U2982 ( .IN1(n3534), .IN2(n284), .IN3(n3538), .IN4(n50), .QN(n3513)
         );
  NOR2X0 U2983 ( .IN1(\fpu_add_frac_dp/n2460 ), .IN2(\fpu_add_frac_dp/n2471 ), 
        .QN(n3253) );
  NOR2X0 U2984 ( .IN1(n3155), .IN2(n584), .QN(n3275) );
  NOR2X0 U2985 ( .IN1(n3155), .IN2(\fpu_add_frac_dp/n2307 ), .QN(n3197) );
  NAND2X0 U2986 ( .IN1(\fpu_add_ctl/n319 ), .IN2(n1449), .QN(n3155) );
  NOR2X0 U2987 ( .IN1(n63), .IN2(n3072), .QN(n3541) );
  INVX0 U2988 ( .INP(n2991), .ZN(n3072) );
  MUX21X1 U2989 ( .IN1(n3543), .IN2(n3533), .S(\fpu_add_frac_dp/n2460 ), .Q(
        n2991) );
  AO22X1 U2990 ( .IN1(n3534), .IN2(n115), .IN3(n3538), .IN4(n48), .Q(n3533) );
  NOR2X0 U2991 ( .IN1(\fpu_add_frac_dp/n2449 ), .IN2(\fpu_add_frac_dp/n586 ), 
        .QN(n3538) );
  AND2X1 U2992 ( .IN1(n219), .IN2(n3534), .Q(n3543) );
  NOR2X0 U2993 ( .IN1(n154), .IN2(\fpu_add_frac_dp/n586 ), .QN(n3534) );
  NAND2X0 U2994 ( .IN1(\fpu_add_ctl/a3stg_opdec_9_0[3] ), .IN2(n1449), .QN(
        n3071) );
  INVX0 U2995 ( .INP(n3136), .ZN(\fpu_add_frac_dp/n1566 ) );
  XNOR3X1 U2996 ( .IN1(\fpu_add_frac_dp/n726 ), .IN2(\fpu_add_frac_dp/n511 ), 
        .IN3(n3544), .Q(n3136) );
  NAND2X0 U2997 ( .IN1(n3142), .IN2(n3545), .QN(n3157) );
  NAND2X0 U2998 ( .IN1(n1449), .IN2(n3546), .QN(n3156) );
  AO21X1 U2999 ( .IN1(n3547), .IN2(n133), .IN3(n336), .Q(n3546) );
  INVX0 U3000 ( .INP(n3135), .ZN(\fpu_add_frac_dp/n1565 ) );
  XNOR3X1 U3001 ( .IN1(\fpu_add_frac_dp/n725 ), .IN2(\fpu_add_frac_dp/n512 ), 
        .IN3(n3548), .Q(n3135) );
  AND4X1 U3002 ( .IN1(n3146), .IN2(n2601), .IN3(n3142), .IN4(n3175), .Q(
        \fpu_add_frac_dp/i_a4stg_rnd_frac_pre1/N66 ) );
  NOR2X0 U3003 ( .IN1(n1745), .IN2(\fpu_add_ctl/n141 ), .QN(n3142) );
  MUX21X1 U3004 ( .IN1(n3549), .IN2(n1330), .S(n3550), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N9 ) );
  OA221X1 U3005 ( .IN1(\fpu_add_frac_dp/n507 ), .IN2(n1312), .IN3(n3551), 
        .IN4(n3552), .IN5(n3553), .Q(n3550) );
  OA21X1 U3006 ( .IN1(n3554), .IN2(n3555), .IN3(n3556), .Q(n3553) );
  MUX21X1 U3007 ( .IN1(n3549), .IN2(n1331), .S(n3557), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N8 ) );
  OA221X1 U3008 ( .IN1(\fpu_add_frac_dp/n508 ), .IN2(n1313), .IN3(n3558), 
        .IN4(n3555), .IN5(n3559), .Q(n3557) );
  OA21X1 U3009 ( .IN1(n3554), .IN2(n3552), .IN3(n3556), .Q(n3559) );
  AOI221X1 U3010 ( .IN1(n3560), .IN2(n3561), .IN3(n3562), .IN4(n3563), .IN5(
        n3564), .QN(n3554) );
  AO22X1 U3011 ( .IN1(n3565), .IN2(n3566), .IN3(n3567), .IN4(n3568), .Q(n3564)
         );
  MUX21X1 U3012 ( .IN1(n3549), .IN2(n1332), .S(n3569), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N7 ) );
  OA221X1 U3013 ( .IN1(\fpu_add_frac_dp/n506 ), .IN2(n1314), .IN3(n3570), 
        .IN4(n3555), .IN5(n3571), .Q(n3569) );
  OA21X1 U3014 ( .IN1(n3558), .IN2(n3552), .IN3(n3556), .Q(n3571) );
  AOI221X1 U3015 ( .IN1(n3562), .IN2(n3572), .IN3(n3567), .IN4(n3573), .IN5(
        n3574), .QN(n3558) );
  AO22X1 U3016 ( .IN1(n3565), .IN2(n3575), .IN3(n3560), .IN4(n3576), .Q(n3574)
         );
  MUX21X1 U3017 ( .IN1(n3549), .IN2(n1330), .S(n3577), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N66 ) );
  OA22X1 U3018 ( .IN1(n3578), .IN2(n3579), .IN3(\fpu_add_frac_dp/n569 ), .IN4(
        n1312), .Q(n3577) );
  MUX21X1 U3019 ( .IN1(n3549), .IN2(n1331), .S(n3580), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N65 ) );
  OA221X1 U3020 ( .IN1(\fpu_add_frac_dp/n568 ), .IN2(n1311), .IN3(n3581), 
        .IN4(n3582), .IN5(n3583), .Q(n3580) );
  OA21X1 U3021 ( .IN1(n3578), .IN2(n3584), .IN3(n3556), .Q(n3583) );
  MUX21X1 U3022 ( .IN1(n3549), .IN2(n1332), .S(n3585), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N64 ) );
  OA221X1 U3023 ( .IN1(\fpu_add_frac_dp/n567 ), .IN2(n1312), .IN3(n3586), 
        .IN4(n3582), .IN5(n3587), .Q(n3585) );
  OA21X1 U3024 ( .IN1(n3581), .IN2(n3588), .IN3(n3556), .Q(n3587) );
  AOI22X1 U3025 ( .IN1(n3589), .IN2(n166), .IN3(n3590), .IN4(n3591), .QN(n3581) );
  NOR2X0 U3026 ( .IN1(\fpu_add_frac_dp/n2270 ), .IN2(n641), .QN(n3590) );
  INVX0 U3027 ( .INP(n3578), .ZN(n3589) );
  NAND2X0 U3028 ( .IN1(n3591), .IN2(n15), .QN(n3578) );
  MUX21X1 U3029 ( .IN1(n3549), .IN2(n1330), .S(n3592), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N63 ) );
  OA221X1 U3030 ( .IN1(\fpu_add_frac_dp/n566 ), .IN2(n1313), .IN3(n3593), 
        .IN4(n3579), .IN5(n3594), .Q(n3592) );
  OA221X1 U3031 ( .IN1(n3586), .IN2(n3588), .IN3(n3582), .IN4(n3595), .IN5(
        n3556), .Q(n3594) );
  NAND2X0 U3032 ( .IN1(n3596), .IN2(n166), .QN(n3595) );
  AOI22X1 U3033 ( .IN1(\fpu_add_frac_dp/n2385 ), .IN2(n3596), .IN3(n3597), 
        .IN4(n3591), .QN(n3586) );
  NOR2X0 U3034 ( .IN1(\fpu_add_frac_dp/n5641 ), .IN2(\fpu_add_frac_dp/n2270 ), 
        .QN(n3597) );
  MUX21X1 U3035 ( .IN1(n3549), .IN2(n1331), .S(n3598), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N62 ) );
  OA221X1 U3036 ( .IN1(\fpu_add_frac_dp/n565 ), .IN2(n1314), .IN3(n3599), 
        .IN4(n3579), .IN5(n3600), .Q(n3598) );
  OA221X1 U3037 ( .IN1(n3593), .IN2(n3601), .IN3(n3602), .IN4(n3603), .IN5(
        n3556), .Q(n3600) );
  INVX0 U3038 ( .INP(n3596), .ZN(n3602) );
  AO22X1 U3039 ( .IN1(n3604), .IN2(n15), .IN3(n3591), .IN4(n3), .Q(n3596) );
  MUX21X1 U3040 ( .IN1(n3549), .IN2(n1332), .S(n3605), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N61 ) );
  OA221X1 U3041 ( .IN1(\fpu_add_frac_dp/n564 ), .IN2(n1311), .IN3(n3606), 
        .IN4(n3579), .IN5(n3607), .Q(n3605) );
  OA221X1 U3042 ( .IN1(n3601), .IN2(n3599), .IN3(n3593), .IN4(n3603), .IN5(
        n3556), .Q(n3607) );
  AOI22X1 U3043 ( .IN1(n3604), .IN2(n16), .IN3(n3591), .IN4(n156), .QN(n3593)
         );
  MUX21X1 U3044 ( .IN1(n3549), .IN2(n1330), .S(n3608), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N60 ) );
  OA221X1 U3045 ( .IN1(\fpu_add_frac_dp/n563 ), .IN2(n1312), .IN3(n3609), 
        .IN4(n3579), .IN5(n3610), .Q(n3608) );
  OA221X1 U3046 ( .IN1(n3601), .IN2(n3606), .IN3(n3599), .IN4(n3603), .IN5(
        n3556), .Q(n3610) );
  AOI222X1 U3047 ( .IN1(n3604), .IN2(n3), .IN3(n3591), .IN4(n68), .IN5(n3611), 
        .IN6(n15), .QN(n3599) );
  MUX21X1 U3048 ( .IN1(n3549), .IN2(n1331), .S(n3612), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N6 ) );
  OA221X1 U3049 ( .IN1(\fpu_add_frac_dp/n505 ), .IN2(n1313), .IN3(n3613), 
        .IN4(n3555), .IN5(n3614), .Q(n3612) );
  OA21X1 U3050 ( .IN1(n3570), .IN2(n3552), .IN3(n3556), .Q(n3614) );
  AOI221X1 U3051 ( .IN1(n3560), .IN2(n3615), .IN3(n3567), .IN4(n3561), .IN5(
        n3616), .QN(n3570) );
  AO22X1 U3052 ( .IN1(n3562), .IN2(n3568), .IN3(n3565), .IN4(n3563), .Q(n3616)
         );
  MUX21X1 U3053 ( .IN1(n3549), .IN2(n1332), .S(n3617), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N59 ) );
  OA221X1 U3054 ( .IN1(\fpu_add_frac_dp/n562 ), .IN2(n1314), .IN3(n3618), 
        .IN4(n3579), .IN5(n3619), .Q(n3617) );
  OA221X1 U3055 ( .IN1(n3601), .IN2(n3609), .IN3(n3606), .IN4(n3603), .IN5(
        n3556), .Q(n3619) );
  AOI222X1 U3056 ( .IN1(n3604), .IN2(n156), .IN3(n3591), .IN4(n1857), .IN5(
        n3611), .IN6(n16), .QN(n3606) );
  MUX21X1 U3057 ( .IN1(n3549), .IN2(n1330), .S(n3620), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N58 ) );
  OA221X1 U3058 ( .IN1(\fpu_add_frac_dp/n561 ), .IN2(n1311), .IN3(n3621), 
        .IN4(n3579), .IN5(n3622), .Q(n3620) );
  OA221X1 U3059 ( .IN1(n3601), .IN2(n3618), .IN3(n3609), .IN4(n3603), .IN5(
        n3556), .Q(n3622) );
  AOI221X1 U3060 ( .IN1(n3591), .IN2(n157), .IN3(n3604), .IN4(n68), .IN5(n3623), .QN(n3609) );
  AO22X1 U3061 ( .IN1(n3624), .IN2(n15), .IN3(n3611), .IN4(n3), .Q(n3623) );
  MUX21X1 U3062 ( .IN1(n3549), .IN2(n1331), .S(n3625), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N57 ) );
  OA221X1 U3063 ( .IN1(\fpu_add_frac_dp/n560 ), .IN2(n1312), .IN3(n3626), 
        .IN4(n3579), .IN5(n3627), .Q(n3625) );
  OA221X1 U3064 ( .IN1(n3601), .IN2(n3621), .IN3(n3618), .IN4(n3603), .IN5(
        n3556), .Q(n3627) );
  AOI221X1 U3065 ( .IN1(n3591), .IN2(n4), .IN3(n3604), .IN4(n1857), .IN5(n3628), .QN(n3618) );
  AO22X1 U3066 ( .IN1(n3624), .IN2(n16), .IN3(n3611), .IN4(n156), .Q(n3628) );
  AND2X1 U3067 ( .IN1(n3629), .IN2(n3560), .Q(n3591) );
  MUX21X1 U3068 ( .IN1(n3549), .IN2(n1332), .S(n3630), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N56 ) );
  OA221X1 U3069 ( .IN1(\fpu_add_frac_dp/n559 ), .IN2(n1313), .IN3(n3631), 
        .IN4(n3579), .IN5(n3632), .Q(n3630) );
  OA221X1 U3070 ( .IN1(n3601), .IN2(n3626), .IN3(n3621), .IN4(n3603), .IN5(
        n3556), .Q(n3632) );
  AOI221X1 U3071 ( .IN1(n3604), .IN2(n157), .IN3(n3611), .IN4(n68), .IN5(n3633), .QN(n3621) );
  AO22X1 U3072 ( .IN1(n3560), .IN2(n3634), .IN3(n3624), .IN4(n3), .Q(n3633) );
  MUX21X1 U3073 ( .IN1(n3549), .IN2(n1330), .S(n3635), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N55 ) );
  OA221X1 U3074 ( .IN1(\fpu_add_frac_dp/n558 ), .IN2(n1314), .IN3(n3636), 
        .IN4(n3579), .IN5(n3637), .Q(n3635) );
  OA221X1 U3075 ( .IN1(n3601), .IN2(n3631), .IN3(n3626), .IN4(n3603), .IN5(
        n3556), .Q(n3637) );
  AOI221X1 U3076 ( .IN1(n3604), .IN2(n4), .IN3(n3611), .IN4(n1857), .IN5(n3638), .QN(n3626) );
  AO22X1 U3077 ( .IN1(n3560), .IN2(n3639), .IN3(n3624), .IN4(n156), .Q(n3638)
         );
  AND2X1 U3078 ( .IN1(n3629), .IN2(n3567), .Q(n3604) );
  MUX21X1 U3079 ( .IN1(n3549), .IN2(n1331), .S(n3640), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N54 ) );
  OA221X1 U3080 ( .IN1(\fpu_add_frac_dp/n557 ), .IN2(n1311), .IN3(n3641), 
        .IN4(n3579), .IN5(n3642), .Q(n3640) );
  OA221X1 U3081 ( .IN1(n3601), .IN2(n3636), .IN3(n3631), .IN4(n3603), .IN5(
        n3556), .Q(n3642) );
  AOI221X1 U3082 ( .IN1(n3611), .IN2(n157), .IN3(n3624), .IN4(n68), .IN5(n3643), .QN(n3631) );
  AO22X1 U3083 ( .IN1(n3560), .IN2(n3644), .IN3(n3567), .IN4(n3634), .Q(n3643)
         );
  MUX21X1 U3084 ( .IN1(n3549), .IN2(n1332), .S(n3645), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N53 ) );
  OA221X1 U3085 ( .IN1(\fpu_add_frac_dp/n556 ), .IN2(n1312), .IN3(n3646), 
        .IN4(n3579), .IN5(n3647), .Q(n3645) );
  OA221X1 U3086 ( .IN1(n3601), .IN2(n3641), .IN3(n3636), .IN4(n3603), .IN5(
        n3556), .Q(n3647) );
  AOI221X1 U3087 ( .IN1(n3611), .IN2(n4), .IN3(n3624), .IN4(n1857), .IN5(n3648), .QN(n3636) );
  AO22X1 U3088 ( .IN1(n3560), .IN2(n3649), .IN3(n3567), .IN4(n3639), .Q(n3648)
         );
  AND2X1 U3089 ( .IN1(n3629), .IN2(n3562), .Q(n3611) );
  MUX21X1 U3090 ( .IN1(n3549), .IN2(n1330), .S(n3650), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N52 ) );
  OA221X1 U3091 ( .IN1(\fpu_add_frac_dp/n555 ), .IN2(n1313), .IN3(n3651), 
        .IN4(n3579), .IN5(n3652), .Q(n3650) );
  OA221X1 U3092 ( .IN1(n3601), .IN2(n3646), .IN3(n3641), .IN4(n3603), .IN5(
        n3556), .Q(n3652) );
  AOI221X1 U3093 ( .IN1(n3624), .IN2(n157), .IN3(n3562), .IN4(n3634), .IN5(
        n3653), .QN(n3641) );
  AO22X1 U3094 ( .IN1(n3560), .IN2(n3654), .IN3(n3567), .IN4(n3644), .Q(n3653)
         );
  MUX21X1 U3095 ( .IN1(n3549), .IN2(n1331), .S(n3655), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N51 ) );
  OA221X1 U3096 ( .IN1(\fpu_add_frac_dp/n554 ), .IN2(n1314), .IN3(n3656), 
        .IN4(n3579), .IN5(n3657), .Q(n3655) );
  OA221X1 U3097 ( .IN1(n3601), .IN2(n3651), .IN3(n3646), .IN4(n3603), .IN5(
        n3556), .Q(n3657) );
  AOI221X1 U3098 ( .IN1(n3624), .IN2(n4), .IN3(n3562), .IN4(n3639), .IN5(n3658), .QN(n3646) );
  AO22X1 U3099 ( .IN1(n3560), .IN2(n3659), .IN3(n3567), .IN4(n3649), .Q(n3658)
         );
  AND2X1 U3100 ( .IN1(n3629), .IN2(n3565), .Q(n3624) );
  MUX21X1 U3101 ( .IN1(n3549), .IN2(n1332), .S(n3660), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N50 ) );
  OA221X1 U3102 ( .IN1(\fpu_add_frac_dp/n553 ), .IN2(n1311), .IN3(n3661), 
        .IN4(n3579), .IN5(n3662), .Q(n3660) );
  OA221X1 U3103 ( .IN1(n3601), .IN2(n3656), .IN3(n3651), .IN4(n3603), .IN5(
        n3556), .Q(n3662) );
  AOI221X1 U3104 ( .IN1(n3567), .IN2(n3654), .IN3(n3560), .IN4(n3663), .IN5(
        n3664), .QN(n3651) );
  AO22X1 U3105 ( .IN1(n3562), .IN2(n3644), .IN3(n3565), .IN4(n3634), .Q(n3664)
         );
  AO22X1 U3106 ( .IN1(n3665), .IN2(n15), .IN3(n3629), .IN4(n98), .Q(n3634) );
  MUX21X1 U3107 ( .IN1(n3549), .IN2(n1330), .S(n3666), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N5 ) );
  OA221X1 U3108 ( .IN1(\fpu_add_frac_dp/n504 ), .IN2(n1312), .IN3(n3667), 
        .IN4(n3555), .IN5(n3668), .Q(n3666) );
  OA21X1 U3109 ( .IN1(n3613), .IN2(n3552), .IN3(n3556), .Q(n3668) );
  AOI221X1 U3110 ( .IN1(n3560), .IN2(n3669), .IN3(n3567), .IN4(n3576), .IN5(
        n3670), .QN(n3613) );
  AO22X1 U3111 ( .IN1(n3565), .IN2(n3572), .IN3(n3562), .IN4(n3573), .Q(n3670)
         );
  MUX21X1 U3112 ( .IN1(n3549), .IN2(n1331), .S(n3671), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N49 ) );
  OA221X1 U3113 ( .IN1(\fpu_add_frac_dp/n552 ), .IN2(n1313), .IN3(n3672), 
        .IN4(n3579), .IN5(n3673), .Q(n3671) );
  OA221X1 U3114 ( .IN1(n3601), .IN2(n3661), .IN3(n3656), .IN4(n3603), .IN5(
        n3556), .Q(n3673) );
  AOI221X1 U3115 ( .IN1(n3567), .IN2(n3659), .IN3(n3560), .IN4(n3674), .IN5(
        n3675), .QN(n3656) );
  AO22X1 U3116 ( .IN1(n3562), .IN2(n3649), .IN3(n3565), .IN4(n3639), .Q(n3675)
         );
  AO22X1 U3117 ( .IN1(n3665), .IN2(n16), .IN3(n3629), .IN4(n97), .Q(n3639) );
  MUX21X1 U3118 ( .IN1(n3549), .IN2(n1332), .S(n3676), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N48 ) );
  OA221X1 U3119 ( .IN1(\fpu_add_frac_dp/n551 ), .IN2(n1314), .IN3(n3677), 
        .IN4(n3579), .IN5(n3678), .Q(n3676) );
  OA221X1 U3120 ( .IN1(n3601), .IN2(n3672), .IN3(n3661), .IN4(n3603), .IN5(
        n3556), .Q(n3678) );
  AOI221X1 U3121 ( .IN1(n3567), .IN2(n3663), .IN3(n3560), .IN4(n3679), .IN5(
        n3680), .QN(n3661) );
  AO22X1 U3122 ( .IN1(n3562), .IN2(n3654), .IN3(n3565), .IN4(n3644), .Q(n3680)
         );
  AO22X1 U3123 ( .IN1(n3665), .IN2(n3), .IN3(n3629), .IN4(n613), .Q(n3644) );
  MUX21X1 U3124 ( .IN1(n3549), .IN2(n1330), .S(n3681), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N47 ) );
  OA221X1 U3125 ( .IN1(\fpu_add_frac_dp/n550 ), .IN2(n1311), .IN3(n3682), 
        .IN4(n3579), .IN5(n3683), .Q(n3681) );
  OA221X1 U3126 ( .IN1(n3601), .IN2(n3677), .IN3(n3672), .IN4(n3603), .IN5(
        n3556), .Q(n3683) );
  AOI221X1 U3127 ( .IN1(n3567), .IN2(n3674), .IN3(n3560), .IN4(n3684), .IN5(
        n3685), .QN(n3672) );
  AO22X1 U3128 ( .IN1(n3562), .IN2(n3659), .IN3(n3565), .IN4(n3649), .Q(n3685)
         );
  AO22X1 U3129 ( .IN1(n3665), .IN2(n156), .IN3(n3629), .IN4(n95), .Q(n3649) );
  MUX21X1 U3130 ( .IN1(n3549), .IN2(n1331), .S(n3686), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N46 ) );
  OA221X1 U3131 ( .IN1(\fpu_add_frac_dp/n549 ), .IN2(n1312), .IN3(n3687), 
        .IN4(n3579), .IN5(n3688), .Q(n3686) );
  OA221X1 U3132 ( .IN1(n3601), .IN2(n3682), .IN3(n3677), .IN4(n3603), .IN5(
        n3556), .Q(n3688) );
  AOI221X1 U3133 ( .IN1(n3567), .IN2(n3679), .IN3(n3560), .IN4(n3689), .IN5(
        n3690), .QN(n3677) );
  AO22X1 U3134 ( .IN1(n3562), .IN2(n3663), .IN3(n3565), .IN4(n3654), .Q(n3690)
         );
  AO22X1 U3135 ( .IN1(n3665), .IN2(n68), .IN3(n3629), .IN4(n632), .Q(n3654) );
  MUX21X1 U3136 ( .IN1(n3549), .IN2(n1332), .S(n3691), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N45 ) );
  OA221X1 U3137 ( .IN1(\fpu_add_frac_dp/n548 ), .IN2(n1313), .IN3(n3692), 
        .IN4(n3579), .IN5(n3693), .Q(n3691) );
  OA221X1 U3138 ( .IN1(n3601), .IN2(n3687), .IN3(n3682), .IN4(n3603), .IN5(
        n3556), .Q(n3693) );
  AOI221X1 U3139 ( .IN1(n3567), .IN2(n3684), .IN3(n3560), .IN4(n3694), .IN5(
        n3695), .QN(n3682) );
  AO22X1 U3140 ( .IN1(n3562), .IN2(n3674), .IN3(n3565), .IN4(n3659), .Q(n3695)
         );
  AO22X1 U3141 ( .IN1(n3665), .IN2(n1857), .IN3(n3629), .IN4(n630), .Q(n3659)
         );
  MUX21X1 U3142 ( .IN1(n3549), .IN2(n1330), .S(n3696), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N44 ) );
  OA221X1 U3143 ( .IN1(\fpu_add_frac_dp/n547 ), .IN2(n1314), .IN3(n3697), 
        .IN4(n3579), .IN5(n3698), .Q(n3696) );
  OA221X1 U3144 ( .IN1(n3601), .IN2(n3692), .IN3(n3687), .IN4(n3603), .IN5(
        n3556), .Q(n3698) );
  AOI221X1 U3145 ( .IN1(n3567), .IN2(n3689), .IN3(n3560), .IN4(n3699), .IN5(
        n3700), .QN(n3687) );
  AO22X1 U3146 ( .IN1(n3562), .IN2(n3679), .IN3(n3565), .IN4(n3663), .Q(n3700)
         );
  AO22X1 U3147 ( .IN1(n3665), .IN2(n157), .IN3(n3629), .IN4(n631), .Q(n3663)
         );
  MUX21X1 U3148 ( .IN1(n3549), .IN2(n1331), .S(n3701), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N43 ) );
  OA221X1 U3149 ( .IN1(\fpu_add_frac_dp/n546 ), .IN2(n1311), .IN3(n3702), 
        .IN4(n3579), .IN5(n3703), .Q(n3701) );
  OA221X1 U3150 ( .IN1(n3601), .IN2(n3697), .IN3(n3692), .IN4(n3603), .IN5(
        n3556), .Q(n3703) );
  AOI221X1 U3151 ( .IN1(n3567), .IN2(n3694), .IN3(n3560), .IN4(n3704), .IN5(
        n3705), .QN(n3692) );
  AO22X1 U3152 ( .IN1(n3562), .IN2(n3684), .IN3(n3565), .IN4(n3674), .Q(n3705)
         );
  AO22X1 U3153 ( .IN1(n3665), .IN2(n4), .IN3(n3629), .IN4(n96), .Q(n3674) );
  MUX21X1 U3154 ( .IN1(n3549), .IN2(n1332), .S(n3706), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N42 ) );
  OA221X1 U3155 ( .IN1(\fpu_add_frac_dp/n544 ), .IN2(n1312), .IN3(n3707), 
        .IN4(n3579), .IN5(n3708), .Q(n3706) );
  OA221X1 U3156 ( .IN1(n3601), .IN2(n3702), .IN3(n3697), .IN4(n3603), .IN5(
        n3556), .Q(n3708) );
  AOI221X1 U3157 ( .IN1(n3567), .IN2(n3699), .IN3(n3560), .IN4(n3709), .IN5(
        n3710), .QN(n3697) );
  AO22X1 U3158 ( .IN1(n3562), .IN2(n3689), .IN3(n3565), .IN4(n3679), .Q(n3710)
         );
  AO222X1 U3159 ( .IN1(n3629), .IN2(n217), .IN3(n3711), .IN4(n15), .IN5(n3665), 
        .IN6(n98), .Q(n3679) );
  MUX21X1 U3160 ( .IN1(n3549), .IN2(n1330), .S(n3712), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N41 ) );
  OA221X1 U3161 ( .IN1(\fpu_add_frac_dp/n543 ), .IN2(n1313), .IN3(n3713), 
        .IN4(n3579), .IN5(n3714), .Q(n3712) );
  OA221X1 U3162 ( .IN1(n3601), .IN2(n3707), .IN3(n3702), .IN4(n3603), .IN5(
        n3556), .Q(n3714) );
  AOI221X1 U3163 ( .IN1(n3567), .IN2(n3704), .IN3(n3560), .IN4(n3715), .IN5(
        n3716), .QN(n3702) );
  AO22X1 U3164 ( .IN1(n3562), .IN2(n3694), .IN3(n3565), .IN4(n3684), .Q(n3716)
         );
  AO222X1 U3165 ( .IN1(n3629), .IN2(n280), .IN3(n3711), .IN4(n16), .IN5(n3665), 
        .IN6(n97), .Q(n3684) );
  MUX21X1 U3166 ( .IN1(n3549), .IN2(n1331), .S(n3717), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N40 ) );
  OA221X1 U3167 ( .IN1(\fpu_add_frac_dp/n542 ), .IN2(n1314), .IN3(n3718), 
        .IN4(n3579), .IN5(n3719), .Q(n3717) );
  OA221X1 U3168 ( .IN1(n3601), .IN2(n3713), .IN3(n3707), .IN4(n3603), .IN5(
        n3556), .Q(n3719) );
  AOI221X1 U3169 ( .IN1(n3565), .IN2(n3689), .IN3(n3562), .IN4(n3699), .IN5(
        n3720), .QN(n3707) );
  AO22X1 U3170 ( .IN1(n3560), .IN2(n3721), .IN3(n3567), .IN4(n3709), .Q(n3720)
         );
  AO222X1 U3171 ( .IN1(n3629), .IN2(n281), .IN3(n3711), .IN4(n3), .IN5(n3665), 
        .IN6(n613), .Q(n3689) );
  MUX21X1 U3172 ( .IN1(n3549), .IN2(n1332), .S(n3722), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N4 ) );
  OA221X1 U3173 ( .IN1(\fpu_add_frac_dp/n503 ), .IN2(n1311), .IN3(n3723), 
        .IN4(n3555), .IN5(n3724), .Q(n3722) );
  OA21X1 U3174 ( .IN1(n3667), .IN2(n3552), .IN3(n3556), .Q(n3724) );
  AOI221X1 U3175 ( .IN1(n3560), .IN2(n3725), .IN3(n3567), .IN4(n3615), .IN5(
        n3726), .QN(n3667) );
  AO22X1 U3176 ( .IN1(n3565), .IN2(n3568), .IN3(n3562), .IN4(n3561), .Q(n3726)
         );
  MUX21X1 U3177 ( .IN1(n3549), .IN2(n1330), .S(n3727), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N39 ) );
  OA221X1 U3178 ( .IN1(\fpu_add_frac_dp/n541 ), .IN2(n1312), .IN3(n3728), 
        .IN4(n3579), .IN5(n3729), .Q(n3727) );
  OA221X1 U3179 ( .IN1(n3601), .IN2(n3718), .IN3(n3713), .IN4(n3603), .IN5(
        n3556), .Q(n3729) );
  AOI221X1 U3180 ( .IN1(n3565), .IN2(n3694), .IN3(n3562), .IN4(n3704), .IN5(
        n3730), .QN(n3713) );
  AO22X1 U3181 ( .IN1(n3560), .IN2(n3731), .IN3(n3567), .IN4(n3715), .Q(n3730)
         );
  AO222X1 U3182 ( .IN1(n3629), .IN2(n638), .IN3(n3711), .IN4(n156), .IN5(n3665), .IN6(n95), .Q(n3694) );
  MUX21X1 U3183 ( .IN1(n3549), .IN2(n1331), .S(n3732), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N38 ) );
  OA221X1 U3184 ( .IN1(\fpu_add_frac_dp/n540 ), .IN2(n1313), .IN3(n3733), 
        .IN4(n3579), .IN5(n3734), .Q(n3732) );
  OA221X1 U3185 ( .IN1(n3601), .IN2(n3728), .IN3(n3718), .IN4(n3603), .IN5(
        n3556), .Q(n3734) );
  AOI221X1 U3186 ( .IN1(n3565), .IN2(n3699), .IN3(n3562), .IN4(n3709), .IN5(
        n3735), .QN(n3718) );
  AO22X1 U3187 ( .IN1(n3560), .IN2(n3736), .IN3(n3567), .IN4(n3721), .Q(n3735)
         );
  AO222X1 U3188 ( .IN1(n3629), .IN2(n174), .IN3(n3711), .IN4(n68), .IN5(n3665), 
        .IN6(n632), .Q(n3699) );
  MUX21X1 U3189 ( .IN1(n3549), .IN2(n1332), .S(n3737), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N37 ) );
  OA221X1 U3190 ( .IN1(\fpu_add_frac_dp/n539 ), .IN2(n1314), .IN3(n3738), 
        .IN4(n3579), .IN5(n3739), .Q(n3737) );
  OA221X1 U3191 ( .IN1(n3601), .IN2(n3733), .IN3(n3728), .IN4(n3603), .IN5(
        n3556), .Q(n3739) );
  AOI221X1 U3192 ( .IN1(n3565), .IN2(n3704), .IN3(n3562), .IN4(n3715), .IN5(
        n3740), .QN(n3728) );
  AO22X1 U3193 ( .IN1(n3560), .IN2(n3741), .IN3(n3567), .IN4(n3731), .Q(n3740)
         );
  AO222X1 U3194 ( .IN1(n3629), .IN2(n70), .IN3(n3711), .IN4(n1857), .IN5(n3665), .IN6(n630), .Q(n3704) );
  MUX21X1 U3195 ( .IN1(n3549), .IN2(n1330), .S(n3742), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N36 ) );
  OA221X1 U3196 ( .IN1(\fpu_add_frac_dp/n538 ), .IN2(n1311), .IN3(n3743), 
        .IN4(n3579), .IN5(n3744), .Q(n3742) );
  OA221X1 U3197 ( .IN1(n3601), .IN2(n3738), .IN3(n3733), .IN4(n3603), .IN5(
        n3556), .Q(n3744) );
  AOI221X1 U3198 ( .IN1(n3565), .IN2(n3709), .IN3(n3562), .IN4(n3721), .IN5(
        n3745), .QN(n3733) );
  AO22X1 U3199 ( .IN1(n3560), .IN2(n1952), .IN3(n3567), .IN4(n3736), .Q(n3745)
         );
  AO222X1 U3200 ( .IN1(n3629), .IN2(\fpu_add_frac_dp/n2380 ), .IN3(n3711), 
        .IN4(n157), .IN5(n3665), .IN6(n631), .Q(n3709) );
  MUX21X1 U3201 ( .IN1(n3549), .IN2(n1331), .S(n3746), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N35 ) );
  OA221X1 U3202 ( .IN1(\fpu_add_frac_dp/n537 ), .IN2(n1312), .IN3(n3738), 
        .IN4(n3603), .IN5(n3747), .Q(n3746) );
  OA221X1 U3203 ( .IN1(n3748), .IN2(n3579), .IN3(n3601), .IN4(n3743), .IN5(
        n3556), .Q(n3747) );
  OA21X1 U3204 ( .IN1(n3582), .IN2(\fpu_add_frac_dp/n5641 ), .IN3(n3584), .Q(
        n3601) );
  OR2X1 U3205 ( .IN1(n3582), .IN2(n641), .Q(n3579) );
  NAND2X0 U3206 ( .IN1(n3749), .IN2(n3750), .QN(n3582) );
  AO21X1 U3207 ( .IN1(n3751), .IN2(n1313), .IN3(n3752), .Q(n3750) );
  AO22X1 U3208 ( .IN1(n3753), .IN2(n553), .IN3(n3754), .IN4(n1022), .Q(n3751)
         );
  AOI221X1 U3209 ( .IN1(n3565), .IN2(n3715), .IN3(n3562), .IN4(n3731), .IN5(
        n3755), .QN(n3738) );
  AO22X1 U3210 ( .IN1(n3560), .IN2(n1950), .IN3(n3567), .IN4(n3741), .Q(n3755)
         );
  AO222X1 U3211 ( .IN1(n3629), .IN2(n168), .IN3(n3711), .IN4(n4), .IN5(n3665), 
        .IN6(n96), .Q(n3715) );
  AND2X1 U3212 ( .IN1(n3756), .IN2(n1063), .Q(n3665) );
  AND2X1 U3213 ( .IN1(n3757), .IN2(n580), .Q(n3711) );
  AND2X1 U3214 ( .IN1(n3756), .IN2(n580), .Q(n3629) );
  MUX21X1 U3215 ( .IN1(n3549), .IN2(n1332), .S(n3758), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N34 ) );
  OA221X1 U3216 ( .IN1(\fpu_add_frac_dp/n536 ), .IN2(n1313), .IN3(n3759), 
        .IN4(n3555), .IN5(n3760), .Q(n3758) );
  OA221X1 U3217 ( .IN1(n3748), .IN2(n3761), .IN3(n3743), .IN4(n3603), .IN5(
        n3556), .Q(n3760) );
  AOI221X1 U3218 ( .IN1(n3567), .IN2(n1952), .IN3(n3560), .IN4(n1951), .IN5(
        n3762), .QN(n3743) );
  AO22X1 U3219 ( .IN1(n3562), .IN2(n3736), .IN3(n3565), .IN4(n3721), .Q(n3762)
         );
  AO222X1 U3220 ( .IN1(n3763), .IN2(n217), .IN3(n3764), .IN4(n15), .IN5(n3765), 
        .IN6(n580), .Q(n3721) );
  MUX21X1 U3221 ( .IN1(n3549), .IN2(n1330), .S(n3766), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N33 ) );
  OA221X1 U3222 ( .IN1(\fpu_add_frac_dp/n535 ), .IN2(n1314), .IN3(n1954), 
        .IN4(n3555), .IN5(n3767), .Q(n3766) );
  OA221X1 U3223 ( .IN1(n3759), .IN2(n3761), .IN3(n3748), .IN4(n3603), .IN5(
        n3556), .Q(n3767) );
  INVX0 U3224 ( .INP(n1948), .ZN(n3748) );
  AO221X1 U3225 ( .IN1(n3567), .IN2(n1950), .IN3(n3560), .IN4(n1949), .IN5(
        n3768), .Q(n1948) );
  AO22X1 U3226 ( .IN1(n3562), .IN2(n3741), .IN3(n3565), .IN4(n3731), .Q(n3768)
         );
  AO222X1 U3227 ( .IN1(n3763), .IN2(n280), .IN3(n3764), .IN4(n16), .IN5(n3769), 
        .IN6(n580), .Q(n3731) );
  MUX21X1 U3228 ( .IN1(n3549), .IN2(n1331), .S(n3770), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N32 ) );
  OA221X1 U3229 ( .IN1(\fpu_add_frac_dp/n534 ), .IN2(n1311), .IN3(n3771), 
        .IN4(n3555), .IN5(n3772), .Q(n3770) );
  OA221X1 U3230 ( .IN1(n1954), .IN2(n3761), .IN3(n3759), .IN4(n3603), .IN5(
        n3556), .Q(n3772) );
  INVX0 U3231 ( .INP(n1945), .ZN(n3759) );
  AO221X1 U3232 ( .IN1(n3567), .IN2(n1951), .IN3(n3560), .IN4(n1963), .IN5(
        n3773), .Q(n1945) );
  AO22X1 U3233 ( .IN1(n3562), .IN2(n1952), .IN3(n3565), .IN4(n3736), .Q(n3773)
         );
  AO222X1 U3234 ( .IN1(n3763), .IN2(n281), .IN3(n3764), .IN4(n3), .IN5(n3774), 
        .IN6(n580), .Q(n3736) );
  MUX21X1 U3235 ( .IN1(n3549), .IN2(n1332), .S(n3775), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N31 ) );
  OA221X1 U3236 ( .IN1(\fpu_add_frac_dp/n533 ), .IN2(n1312), .IN3(n3776), 
        .IN4(n3555), .IN5(n3777), .Q(n3775) );
  OA221X1 U3237 ( .IN1(n3761), .IN2(n3771), .IN3(n1954), .IN4(n3603), .IN5(
        n3556), .Q(n3777) );
  AOI221X1 U3238 ( .IN1(n3567), .IN2(n1949), .IN3(n3560), .IN4(n1964), .IN5(
        n3778), .QN(n1954) );
  AO22X1 U3239 ( .IN1(n3562), .IN2(n1950), .IN3(n3565), .IN4(n3741), .Q(n3778)
         );
  AO222X1 U3240 ( .IN1(n3763), .IN2(n638), .IN3(n3764), .IN4(n156), .IN5(n3779), .IN6(n580), .Q(n3741) );
  MUX21X1 U3241 ( .IN1(n3549), .IN2(n1330), .S(n3780), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N30 ) );
  OA221X1 U3242 ( .IN1(\fpu_add_frac_dp/n532 ), .IN2(n1313), .IN3(n3781), 
        .IN4(n3555), .IN5(n3782), .Q(n3780) );
  OA221X1 U3243 ( .IN1(n3761), .IN2(n3776), .IN3(n3771), .IN4(n3603), .IN5(
        n3556), .Q(n3782) );
  AOI221X1 U3244 ( .IN1(n3567), .IN2(n1963), .IN3(n3560), .IN4(n1972), .IN5(
        n3783), .QN(n3771) );
  AO22X1 U3245 ( .IN1(n3562), .IN2(n1951), .IN3(n3565), .IN4(n1952), .Q(n3783)
         );
  AO222X1 U3246 ( .IN1(n3763), .IN2(n174), .IN3(n3764), .IN4(n68), .IN5(n1946), 
        .IN6(n580), .Q(n1952) );
  MUX21X1 U3247 ( .IN1(n3549), .IN2(n1331), .S(n3784), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N3 ) );
  OA221X1 U3248 ( .IN1(\fpu_add_frac_dp/n509 ), .IN2(n1314), .IN3(n3723), 
        .IN4(n3552), .IN5(n3785), .Q(n3784) );
  OA21X1 U3249 ( .IN1(n3786), .IN2(n3555), .IN3(n3556), .Q(n3785) );
  AOI221X1 U3250 ( .IN1(n3561), .IN2(n3565), .IN3(n3615), .IN4(n3562), .IN5(
        n3787), .QN(n3786) );
  AO22X1 U3251 ( .IN1(n3788), .IN2(n3560), .IN3(n3725), .IN4(n3567), .Q(n3787)
         );
  AO22X1 U3252 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n1976), .IN3(n1960), 
        .IN4(n580), .Q(n3725) );
  AO222X1 U3253 ( .IN1(n3789), .IN2(n690), .IN3(n3790), .IN4(n2653), .IN5(
        n3791), .IN6(\fpu_add_frac_dp/n2393 ), .Q(n1960) );
  AO22X1 U3254 ( .IN1(n580), .IN2(n1959), .IN3(n1977), .IN4(
        \fpu_add_frac_dp/n2397 ), .Q(n3788) );
  AO222X1 U3255 ( .IN1(n3789), .IN2(n896), .IN3(n3792), .IN4(n2653), .IN5(
        n3791), .IN6(n218), .Q(n1959) );
  AO22X1 U3256 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n2027), .IN3(n1957), 
        .IN4(n580), .Q(n3615) );
  AO222X1 U3257 ( .IN1(n3789), .IN2(n660), .IN3(n3793), .IN4(n2653), .IN5(
        n3791), .IN6(n6), .Q(n1957) );
  AO22X1 U3258 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n1989), .IN3(n1958), 
        .IN4(n580), .Q(n3561) );
  AO222X1 U3259 ( .IN1(n3789), .IN2(n655), .IN3(n3794), .IN4(n2653), .IN5(
        n3791), .IN6(n23), .Q(n1958) );
  AOI221X1 U3260 ( .IN1(n3560), .IN2(n3795), .IN3(n3567), .IN4(n3669), .IN5(
        n3796), .QN(n3723) );
  AO22X1 U3261 ( .IN1(n3565), .IN2(n3573), .IN3(n3562), .IN4(n3576), .Q(n3796)
         );
  AO22X1 U3262 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n2026), .IN3(n1966), 
        .IN4(n580), .Q(n3576) );
  AO222X1 U3263 ( .IN1(n3789), .IN2(n898), .IN3(n3797), .IN4(n2653), .IN5(
        n3791), .IN6(n162), .Q(n1966) );
  AO22X1 U3264 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n1990), .IN3(n1967), 
        .IN4(n580), .Q(n3669) );
  AO222X1 U3265 ( .IN1(n3789), .IN2(n899), .IN3(n3798), .IN4(n2653), .IN5(
        n3791), .IN6(n205), .Q(n1967) );
  AO22X1 U3266 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n1996), .IN3(n1965), 
        .IN4(n580), .Q(n3795) );
  AO222X1 U3267 ( .IN1(n3789), .IN2(n902), .IN3(n3799), .IN4(n2653), .IN5(
        n3791), .IN6(n278), .Q(n1965) );
  MUX21X1 U3268 ( .IN1(n3549), .IN2(n1332), .S(n3800), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N29 ) );
  OA221X1 U3269 ( .IN1(\fpu_add_frac_dp/n531 ), .IN2(n1311), .IN3(n3801), 
        .IN4(n3555), .IN5(n3802), .Q(n3800) );
  OA221X1 U3270 ( .IN1(n3761), .IN2(n3781), .IN3(n3776), .IN4(n3603), .IN5(
        n3556), .Q(n3802) );
  AOI221X1 U3271 ( .IN1(n3567), .IN2(n1964), .IN3(n3560), .IN4(n1973), .IN5(
        n3803), .QN(n3776) );
  AO22X1 U3272 ( .IN1(n3562), .IN2(n1949), .IN3(n3565), .IN4(n1950), .Q(n3803)
         );
  AO222X1 U3273 ( .IN1(n3763), .IN2(n70), .IN3(n3764), .IN4(n1857), .IN5(n3804), .IN6(n580), .Q(n1950) );
  MUX21X1 U3274 ( .IN1(n3549), .IN2(n1330), .S(n3805), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N28 ) );
  OA221X1 U3275 ( .IN1(\fpu_add_frac_dp/n530 ), .IN2(n1312), .IN3(n3806), 
        .IN4(n3555), .IN5(n3807), .Q(n3805) );
  OA221X1 U3276 ( .IN1(n3761), .IN2(n3801), .IN3(n3781), .IN4(n3603), .IN5(
        n3556), .Q(n3807) );
  AOI221X1 U3277 ( .IN1(n3567), .IN2(n1972), .IN3(n3560), .IN4(n3808), .IN5(
        n3809), .QN(n3781) );
  AO22X1 U3278 ( .IN1(n3562), .IN2(n1963), .IN3(n3565), .IN4(n1951), .Q(n3809)
         );
  AO222X1 U3279 ( .IN1(n3763), .IN2(\fpu_add_frac_dp/n2380 ), .IN3(n3764), 
        .IN4(n157), .IN5(n3810), .IN6(n580), .Q(n1951) );
  MUX21X1 U3280 ( .IN1(n3549), .IN2(n1331), .S(n3811), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N27 ) );
  OA221X1 U3281 ( .IN1(\fpu_add_frac_dp/n529 ), .IN2(n1313), .IN3(n3812), 
        .IN4(n3555), .IN5(n3813), .Q(n3811) );
  OA221X1 U3282 ( .IN1(n3761), .IN2(n3806), .IN3(n3801), .IN4(n3603), .IN5(
        n3556), .Q(n3813) );
  AOI221X1 U3283 ( .IN1(n3567), .IN2(n1973), .IN3(n3560), .IN4(n1971), .IN5(
        n3814), .QN(n3801) );
  AO22X1 U3284 ( .IN1(n3562), .IN2(n1964), .IN3(n3565), .IN4(n1949), .Q(n3814)
         );
  AO222X1 U3285 ( .IN1(n3763), .IN2(n168), .IN3(n3764), .IN4(n4), .IN5(n3815), 
        .IN6(n580), .Q(n1949) );
  AND2X1 U3286 ( .IN1(n3757), .IN2(\fpu_add_frac_dp/n2399 ), .Q(n3764) );
  NOR2X0 U3287 ( .IN1(\fpu_add_frac_dp/n570 ), .IN2(\fpu_add_frac_dp/n577 ), 
        .QN(n3757) );
  AND2X1 U3288 ( .IN1(n3756), .IN2(\fpu_add_frac_dp/n2399 ), .Q(n3763) );
  NOR2X0 U3289 ( .IN1(\fpu_add_frac_dp/n2382 ), .IN2(\fpu_add_frac_dp/n570 ), 
        .QN(n3756) );
  MUX21X1 U3290 ( .IN1(n3549), .IN2(n1332), .S(n3816), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N26 ) );
  OA221X1 U3291 ( .IN1(\fpu_add_frac_dp/n527 ), .IN2(n1314), .IN3(n3817), 
        .IN4(n3555), .IN5(n3818), .Q(n3816) );
  OA221X1 U3292 ( .IN1(n3761), .IN2(n3812), .IN3(n3806), .IN4(n3603), .IN5(
        n3556), .Q(n3818) );
  AOI221X1 U3293 ( .IN1(n3567), .IN2(n3808), .IN3(n3560), .IN4(n1969), .IN5(
        n3819), .QN(n3806) );
  AO22X1 U3294 ( .IN1(n3562), .IN2(n1972), .IN3(n3565), .IN4(n1963), .Q(n3819)
         );
  AO22X1 U3295 ( .IN1(n1982), .IN2(n580), .IN3(\fpu_add_frac_dp/n2399 ), .IN4(
        n3765), .Q(n1963) );
  AO22X1 U3296 ( .IN1(n3820), .IN2(n98), .IN3(n3821), .IN4(n271), .Q(n3765) );
  MUX21X1 U3297 ( .IN1(n3549), .IN2(n1329), .S(n3822), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N25 ) );
  OA221X1 U3298 ( .IN1(\fpu_add_frac_dp/n526 ), .IN2(n1311), .IN3(n3823), 
        .IN4(n3555), .IN5(n3824), .Q(n3822) );
  OA221X1 U3299 ( .IN1(n3761), .IN2(n3817), .IN3(n3812), .IN4(n3603), .IN5(
        n3556), .Q(n3824) );
  AOI221X1 U3300 ( .IN1(n3567), .IN2(n1971), .IN3(n3560), .IN4(n1968), .IN5(
        n3825), .QN(n3812) );
  AO22X1 U3301 ( .IN1(n3562), .IN2(n1973), .IN3(n3565), .IN4(n1964), .Q(n3825)
         );
  AO22X1 U3302 ( .IN1(n1981), .IN2(n580), .IN3(\fpu_add_frac_dp/n2399 ), .IN4(
        n3769), .Q(n1964) );
  AO22X1 U3303 ( .IN1(n3820), .IN2(n97), .IN3(n3821), .IN4(n23), .Q(n3769) );
  MUX21X1 U3304 ( .IN1(n3549), .IN2(n1329), .S(n3826), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N24 ) );
  OA221X1 U3305 ( .IN1(\fpu_add_frac_dp/n525 ), .IN2(n1312), .IN3(n3827), 
        .IN4(n3555), .IN5(n3828), .Q(n3826) );
  OA221X1 U3306 ( .IN1(n3761), .IN2(n3823), .IN3(n3817), .IN4(n3603), .IN5(
        n3556), .Q(n3828) );
  AOI221X1 U3307 ( .IN1(n3567), .IN2(n1969), .IN3(n3560), .IN4(n3829), .IN5(
        n3830), .QN(n3817) );
  AO22X1 U3308 ( .IN1(n3562), .IN2(n3808), .IN3(n3565), .IN4(n1972), .Q(n3830)
         );
  AO22X1 U3309 ( .IN1(n1983), .IN2(n580), .IN3(\fpu_add_frac_dp/n2399 ), .IN4(
        n3774), .Q(n1972) );
  AO22X1 U3310 ( .IN1(n3820), .IN2(n613), .IN3(n3821), .IN4(n162), .Q(n3774)
         );
  MUX21X1 U3311 ( .IN1(n3549), .IN2(n1329), .S(n3831), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N23 ) );
  OA221X1 U3312 ( .IN1(\fpu_add_frac_dp/n524 ), .IN2(n1313), .IN3(n3832), 
        .IN4(n3555), .IN5(n3833), .Q(n3831) );
  OA221X1 U3313 ( .IN1(n3761), .IN2(n3827), .IN3(n3823), .IN4(n3603), .IN5(
        n3556), .Q(n3833) );
  AOI221X1 U3314 ( .IN1(n3567), .IN2(n1968), .IN3(n3560), .IN4(n3834), .IN5(
        n3835), .QN(n3823) );
  AO22X1 U3315 ( .IN1(n3562), .IN2(n1971), .IN3(n3565), .IN4(n1973), .Q(n3835)
         );
  AO22X1 U3316 ( .IN1(n1985), .IN2(n580), .IN3(\fpu_add_frac_dp/n2399 ), .IN4(
        n3779), .Q(n1973) );
  AO22X1 U3317 ( .IN1(n3820), .IN2(n95), .IN3(n3821), .IN4(n6), .Q(n3779) );
  MUX21X1 U3318 ( .IN1(n3549), .IN2(n1329), .S(n3836), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N22 ) );
  OA221X1 U3319 ( .IN1(\fpu_add_frac_dp/n523 ), .IN2(n1314), .IN3(n3837), 
        .IN4(n3555), .IN5(n3838), .Q(n3836) );
  OA221X1 U3320 ( .IN1(n3761), .IN2(n3832), .IN3(n3827), .IN4(n3603), .IN5(
        n3556), .Q(n3838) );
  AOI221X1 U3321 ( .IN1(n3567), .IN2(n3829), .IN3(n3560), .IN4(n3839), .IN5(
        n3840), .QN(n3827) );
  AO22X1 U3322 ( .IN1(n3562), .IN2(n1969), .IN3(n3565), .IN4(n3808), .Q(n3840)
         );
  AO22X1 U3323 ( .IN1(n1986), .IN2(n580), .IN3(\fpu_add_frac_dp/n2399 ), .IN4(
        n1946), .Q(n3808) );
  AO22X1 U3324 ( .IN1(n3820), .IN2(n632), .IN3(n3821), .IN4(n205), .Q(n1946)
         );
  MUX21X1 U3325 ( .IN1(n3549), .IN2(n1329), .S(n3841), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N21 ) );
  OA221X1 U3326 ( .IN1(\fpu_add_frac_dp/n522 ), .IN2(n1311), .IN3(n3842), 
        .IN4(n3555), .IN5(n3843), .Q(n3841) );
  OA221X1 U3327 ( .IN1(n3761), .IN2(n3837), .IN3(n3832), .IN4(n3603), .IN5(
        n3556), .Q(n3843) );
  AOI221X1 U3328 ( .IN1(n3567), .IN2(n3834), .IN3(n3560), .IN4(n3844), .IN5(
        n3845), .QN(n3832) );
  AO22X1 U3329 ( .IN1(n3562), .IN2(n1968), .IN3(n3565), .IN4(n1971), .Q(n3845)
         );
  AO22X1 U3330 ( .IN1(n1979), .IN2(n580), .IN3(\fpu_add_frac_dp/n2399 ), .IN4(
        n3804), .Q(n1971) );
  AO22X1 U3331 ( .IN1(n3820), .IN2(n630), .IN3(n3821), .IN4(
        \fpu_add_frac_dp/n2393 ), .Q(n3804) );
  MUX21X1 U3332 ( .IN1(n3549), .IN2(n1329), .S(n3846), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N20 ) );
  OA221X1 U3333 ( .IN1(\fpu_add_frac_dp/n521 ), .IN2(n1312), .IN3(n3847), 
        .IN4(n3555), .IN5(n3848), .Q(n3846) );
  OA221X1 U3334 ( .IN1(n3761), .IN2(n3842), .IN3(n3837), .IN4(n3603), .IN5(
        n3556), .Q(n3848) );
  AOI221X1 U3335 ( .IN1(n3567), .IN2(n3839), .IN3(n3560), .IN4(n3849), .IN5(
        n3850), .QN(n3837) );
  AO22X1 U3336 ( .IN1(n3562), .IN2(n3829), .IN3(n3565), .IN4(n1969), .Q(n3850)
         );
  AO22X1 U3337 ( .IN1(n1978), .IN2(n580), .IN3(\fpu_add_frac_dp/n2399 ), .IN4(
        n3810), .Q(n1969) );
  AO22X1 U3338 ( .IN1(n3820), .IN2(n631), .IN3(n3821), .IN4(n278), .Q(n3810)
         );
  MUX21X1 U3339 ( .IN1(n3549), .IN2(n1329), .S(n3851), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N19 ) );
  OA221X1 U3340 ( .IN1(\fpu_add_frac_dp/n520 ), .IN2(n1313), .IN3(n3852), 
        .IN4(n3555), .IN5(n3853), .Q(n3851) );
  OA221X1 U3341 ( .IN1(n3761), .IN2(n3847), .IN3(n3842), .IN4(n3603), .IN5(
        n3556), .Q(n3853) );
  AOI221X1 U3342 ( .IN1(n3567), .IN2(n3844), .IN3(n3560), .IN4(n3854), .IN5(
        n3855), .QN(n3842) );
  AO22X1 U3343 ( .IN1(n3562), .IN2(n3834), .IN3(n3565), .IN4(n1968), .Q(n3855)
         );
  AO22X1 U3344 ( .IN1(n1980), .IN2(n580), .IN3(\fpu_add_frac_dp/n2399 ), .IN4(
        n3815), .Q(n1968) );
  AO22X1 U3345 ( .IN1(n3820), .IN2(n96), .IN3(n3821), .IN4(n218), .Q(n3815) );
  MUX21X1 U3346 ( .IN1(n3549), .IN2(n1329), .S(n3856), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N18 ) );
  OA221X1 U3347 ( .IN1(\fpu_add_frac_dp/n519 ), .IN2(n1314), .IN3(n3857), 
        .IN4(n3555), .IN5(n3858), .Q(n3856) );
  OA221X1 U3348 ( .IN1(n3761), .IN2(n3852), .IN3(n3847), .IN4(n3603), .IN5(
        n3556), .Q(n3858) );
  AOI221X1 U3349 ( .IN1(n3567), .IN2(n3849), .IN3(n3560), .IN4(n3859), .IN5(
        n3860), .QN(n3847) );
  AO22X1 U3350 ( .IN1(n3562), .IN2(n3839), .IN3(n3565), .IN4(n3829), .Q(n3860)
         );
  AO22X1 U3351 ( .IN1(n1991), .IN2(n580), .IN3(n1982), .IN4(n581), .Q(n3829)
         );
  AO222X1 U3352 ( .IN1(n3821), .IN2(n696), .IN3(n3861), .IN4(n15), .IN5(n3820), 
        .IN6(n217), .Q(n1982) );
  MUX21X1 U3353 ( .IN1(n3549), .IN2(n1329), .S(n3862), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N17 ) );
  OA221X1 U3354 ( .IN1(\fpu_add_frac_dp/n518 ), .IN2(n1311), .IN3(n3863), 
        .IN4(n3555), .IN5(n3864), .Q(n3862) );
  OA221X1 U3355 ( .IN1(n3761), .IN2(n3857), .IN3(n3852), .IN4(n3603), .IN5(
        n3556), .Q(n3864) );
  AOI221X1 U3356 ( .IN1(n3567), .IN2(n3854), .IN3(n3560), .IN4(n3865), .IN5(
        n3866), .QN(n3852) );
  AO22X1 U3357 ( .IN1(n3562), .IN2(n3844), .IN3(n3565), .IN4(n3834), .Q(n3866)
         );
  AO22X1 U3358 ( .IN1(n1993), .IN2(n580), .IN3(n1981), .IN4(n581), .Q(n3834)
         );
  AO222X1 U3359 ( .IN1(n3821), .IN2(n678), .IN3(n3861), .IN4(n16), .IN5(n3820), 
        .IN6(n280), .Q(n1981) );
  MUX21X1 U3360 ( .IN1(n3549), .IN2(n1329), .S(n3867), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N16 ) );
  OA221X1 U3361 ( .IN1(\fpu_add_frac_dp/n517 ), .IN2(n1312), .IN3(n3868), 
        .IN4(n3555), .IN5(n3869), .Q(n3867) );
  OA221X1 U3362 ( .IN1(n3761), .IN2(n3863), .IN3(n3857), .IN4(n3603), .IN5(
        n3556), .Q(n3869) );
  AOI221X1 U3363 ( .IN1(n3567), .IN2(n3859), .IN3(n3560), .IN4(n3870), .IN5(
        n3871), .QN(n3857) );
  AO22X1 U3364 ( .IN1(n3562), .IN2(n3849), .IN3(n3565), .IN4(n3839), .Q(n3871)
         );
  AO22X1 U3365 ( .IN1(n1997), .IN2(n580), .IN3(n1983), .IN4(n581), .Q(n3839)
         );
  AO222X1 U3366 ( .IN1(n3821), .IN2(n679), .IN3(n3861), .IN4(n3), .IN5(n3820), 
        .IN6(n281), .Q(n1983) );
  MUX21X1 U3367 ( .IN1(n3549), .IN2(n1329), .S(n3872), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N15 ) );
  OA221X1 U3368 ( .IN1(\fpu_add_frac_dp/n516 ), .IN2(n1313), .IN3(n3873), 
        .IN4(n3555), .IN5(n3874), .Q(n3872) );
  OA221X1 U3369 ( .IN1(n3761), .IN2(n3868), .IN3(n3863), .IN4(n3603), .IN5(
        n3556), .Q(n3874) );
  AOI221X1 U3370 ( .IN1(n3567), .IN2(n3865), .IN3(n3560), .IN4(n3875), .IN5(
        n3876), .QN(n3863) );
  AO22X1 U3371 ( .IN1(n3562), .IN2(n3854), .IN3(n3565), .IN4(n3844), .Q(n3876)
         );
  AO22X1 U3372 ( .IN1(n1992), .IN2(n580), .IN3(n1985), .IN4(n581), .Q(n3844)
         );
  AO222X1 U3373 ( .IN1(n3821), .IN2(n106), .IN3(n3861), .IN4(n156), .IN5(n3820), .IN6(n638), .Q(n1985) );
  NOR2X0 U3374 ( .IN1(\fpu_add_frac_dp/n2382 ), .IN2(\fpu_add_frac_dp/n573 ), 
        .QN(n3861) );
  NOR2X0 U3375 ( .IN1(\fpu_add_frac_dp/n2382 ), .IN2(\fpu_add_frac_dp/n545 ), 
        .QN(n3821) );
  MUX21X1 U3376 ( .IN1(n3549), .IN2(n1329), .S(n3877), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N14 ) );
  OA221X1 U3377 ( .IN1(\fpu_add_frac_dp/n514 ), .IN2(n1314), .IN3(n3878), 
        .IN4(n3555), .IN5(n3879), .Q(n3877) );
  OA221X1 U3378 ( .IN1(n3761), .IN2(n3873), .IN3(n3868), .IN4(n3603), .IN5(
        n3556), .Q(n3879) );
  AOI221X1 U3379 ( .IN1(n3567), .IN2(n3870), .IN3(n3560), .IN4(n3880), .IN5(
        n3881), .QN(n3868) );
  AO22X1 U3380 ( .IN1(n3562), .IN2(n3859), .IN3(n3565), .IN4(n3849), .Q(n3881)
         );
  AO22X1 U3381 ( .IN1(n3882), .IN2(n580), .IN3(n1986), .IN4(n581), .Q(n3849)
         );
  AO22X1 U3382 ( .IN1(n3883), .IN2(n3884), .IN3(n3820), .IN4(n174), .Q(n1986)
         );
  INVX0 U3383 ( .INP(n3885), .ZN(n3883) );
  MUX21X1 U3384 ( .IN1(n3549), .IN2(n1329), .S(n3886), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N13 ) );
  OA221X1 U3385 ( .IN1(\fpu_add_frac_dp/n512 ), .IN2(n1311), .IN3(n3887), 
        .IN4(n3555), .IN5(n3888), .Q(n3886) );
  OA221X1 U3386 ( .IN1(n3761), .IN2(n3878), .IN3(n3873), .IN4(n3603), .IN5(
        n3556), .Q(n3888) );
  AOI221X1 U3387 ( .IN1(n3560), .IN2(n3566), .IN3(n3567), .IN4(n3875), .IN5(
        n3889), .QN(n3873) );
  AO22X1 U3388 ( .IN1(n3562), .IN2(n3865), .IN3(n3565), .IN4(n3854), .Q(n3889)
         );
  AO22X1 U3389 ( .IN1(n3890), .IN2(n580), .IN3(n1979), .IN4(n581), .Q(n3854)
         );
  AO22X1 U3390 ( .IN1(n3891), .IN2(n3884), .IN3(n3820), .IN4(n70), .Q(n1979)
         );
  MUX21X1 U3391 ( .IN1(n3549), .IN2(n1329), .S(n3892), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N12 ) );
  OA221X1 U3392 ( .IN1(\fpu_add_frac_dp/n511 ), .IN2(n1312), .IN3(n3893), 
        .IN4(n3555), .IN5(n3894), .Q(n3892) );
  OA221X1 U3393 ( .IN1(n3761), .IN2(n3887), .IN3(n3878), .IN4(n3603), .IN5(
        n3556), .Q(n3894) );
  AOI221X1 U3394 ( .IN1(n3560), .IN2(n3575), .IN3(n3567), .IN4(n3880), .IN5(
        n3895), .QN(n3878) );
  AO22X1 U3395 ( .IN1(n3562), .IN2(n3870), .IN3(n3565), .IN4(n3859), .Q(n3895)
         );
  AO22X1 U3396 ( .IN1(n3896), .IN2(n580), .IN3(n1978), .IN4(n581), .Q(n3859)
         );
  AO22X1 U3397 ( .IN1(n3897), .IN2(n3884), .IN3(n3820), .IN4(
        \fpu_add_frac_dp/n2380 ), .Q(n1978) );
  MUX21X1 U3398 ( .IN1(n3549), .IN2(n1329), .S(n3898), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N11 ) );
  OA221X1 U3399 ( .IN1(\fpu_add_frac_dp/n502 ), .IN2(n1313), .IN3(n3899), 
        .IN4(n3555), .IN5(n3900), .Q(n3898) );
  OA221X1 U3400 ( .IN1(n3887), .IN2(n3603), .IN3(n3761), .IN4(n3893), .IN5(
        n3556), .Q(n3900) );
  AOI221X1 U3401 ( .IN1(n3562), .IN2(n3880), .IN3(n3560), .IN4(n3572), .IN5(
        n3901), .QN(n3893) );
  AO22X1 U3402 ( .IN1(n3567), .IN2(n3575), .IN3(n3565), .IN4(n3870), .Q(n3901)
         );
  AND2X1 U3403 ( .IN1(n3552), .IN2(n3584), .Q(n3761) );
  NAND2X0 U3404 ( .IN1(n3902), .IN2(\fpu_add_frac_dp/n2385 ), .QN(n3584) );
  NAND2X0 U3405 ( .IN1(n3902), .IN2(n166), .QN(n3603) );
  INVX0 U3406 ( .INP(n3588), .ZN(n3902) );
  AOI221X1 U3407 ( .IN1(n3565), .IN2(n3865), .IN3(n3560), .IN4(n3563), .IN5(
        n3903), .QN(n3887) );
  AO22X1 U3408 ( .IN1(n3562), .IN2(n3875), .IN3(n3567), .IN4(n3566), .Q(n3903)
         );
  AO22X1 U3409 ( .IN1(n3904), .IN2(n580), .IN3(n1980), .IN4(n581), .Q(n3865)
         );
  AO22X1 U3410 ( .IN1(n3905), .IN2(n3884), .IN3(n3820), .IN4(n168), .Q(n1980)
         );
  NOR2X0 U3411 ( .IN1(\fpu_add_frac_dp/n570 ), .IN2(\fpu_add_frac_dp/n576 ), 
        .QN(n3820) );
  MUX21X1 U3412 ( .IN1(n3549), .IN2(n1329), .S(n3906), .Q(
        \fpu_add_frac_dp/i_a3stg_frac2/N10 ) );
  OA221X1 U3413 ( .IN1(\fpu_add_frac_dp/n501 ), .IN2(n1314), .IN3(n3551), 
        .IN4(n3555), .IN5(n3907), .Q(n3906) );
  OA221X1 U3414 ( .IN1(n3908), .IN2(n3588), .IN3(n3899), .IN4(n3552), .IN5(
        n3556), .Q(n3907) );
  NAND3X0 U3415 ( .IN1(n3909), .IN2(n1311), .IN3(\fpu_add_ctl/n329 ), .QN(
        n3556) );
  INVX0 U3416 ( .INP(n3749), .ZN(n3909) );
  NAND3X0 U3417 ( .IN1(n3749), .IN2(n166), .IN3(n3752), .QN(n3552) );
  AOI221X1 U3418 ( .IN1(n3567), .IN2(n3563), .IN3(n3560), .IN4(n3568), .IN5(
        n3910), .QN(n3899) );
  AO22X1 U3419 ( .IN1(n3565), .IN2(n3875), .IN3(n3562), .IN4(n3566), .Q(n3910)
         );
  AO22X1 U3420 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n3904), .IN3(n1977), 
        .IN4(n580), .Q(n3568) );
  AO222X1 U3421 ( .IN1(n3789), .IN2(n659), .IN3(n3905), .IN4(n2653), .IN5(
        n3791), .IN6(n168), .Q(n1977) );
  AO22X1 U3422 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n3890), .IN3(n1976), 
        .IN4(n580), .Q(n3563) );
  AO222X1 U3423 ( .IN1(n3789), .IN2(n161), .IN3(n3891), .IN4(n2653), .IN5(
        n3791), .IN6(n70), .Q(n1976) );
  NAND2X0 U3424 ( .IN1(n1311), .IN2(n356), .QN(n3588) );
  NOR4X0 U3425 ( .IN1(n3911), .IN2(n3912), .IN3(n2029), .IN4(n2041), .QN(n3908) );
  NAND4X0 U3426 ( .IN1(n3913), .IN2(n3914), .IN3(n3915), .IN4(n2004), .QN(
        n2041) );
  OA21X1 U3427 ( .IN1(\fpu_add_frac_dp/n579 ), .IN2(n3916), .IN3(n3917), .Q(
        n3915) );
  NOR4X0 U3428 ( .IN1(n23), .IN2(n3918), .IN3(n162), .IN4(n6), .QN(n3916) );
  NAND2X0 U3429 ( .IN1(\fpu_add_frac_dp/n2497 ), .IN2(\fpu_add_frac_dp/n2424 ), 
        .QN(n3918) );
  AO221X1 U3430 ( .IN1(\fpu_add_frac_dp/n2306 ), .IN2(n3905), .IN3(n168), 
        .IN4(n2638), .IN5(n659), .Q(n2029) );
  AO22X1 U3431 ( .IN1(n118), .IN2(n929), .IN3(n4), .IN4(n47), .Q(n3905) );
  AO21X1 U3432 ( .IN1(n2008), .IN2(n2638), .IN3(n2033), .Q(n3912) );
  NAND4X0 U3433 ( .IN1(n2038), .IN2(n2015), .IN3(n2005), .IN4(n3919), .QN(
        n2033) );
  NOR3X0 U3434 ( .IN1(n2020), .IN2(n3920), .IN3(n2014), .QN(n3919) );
  MUX21X1 U3435 ( .IN1(n3921), .IN2(n3922), .S(\fpu_add_frac_dp/n2306 ), .Q(
        n2014) );
  NAND3X0 U3436 ( .IN1(n3923), .IN2(n2040), .IN3(n2039), .QN(n3922) );
  NAND4X0 U3437 ( .IN1(n3914), .IN2(\fpu_add_frac_dp/n771 ), .IN3(n2004), 
        .IN4(n3924), .QN(n3921) );
  NAND2X0 U3438 ( .IN1(n205), .IN2(n2638), .QN(n3924) );
  OA21X1 U3439 ( .IN1(\fpu_add_frac_dp/n741 ), .IN2(\fpu_add_frac_dp/n579 ), 
        .IN3(\fpu_add_frac_dp/n773 ), .Q(n2004) );
  INVX0 U3440 ( .INP(n2043), .ZN(n3914) );
  AO21X1 U3441 ( .IN1(\fpu_add_frac_dp/n2393 ), .IN2(n2638), .IN3(n690), .Q(
        n2043) );
  OA21X1 U3442 ( .IN1(n3925), .IN2(n3926), .IN3(n2019), .Q(n3920) );
  NAND3X0 U3443 ( .IN1(n3927), .IN2(n624), .IN3(\fpu_add_frac_dp/n769 ), .QN(
        n2019) );
  NAND2X0 U3444 ( .IN1(n2638), .IN2(n162), .QN(n3927) );
  INVX0 U3445 ( .INP(n2022), .ZN(n3925) );
  NOR2X0 U3446 ( .IN1(n3797), .IN2(n624), .QN(n2022) );
  AO221X1 U3447 ( .IN1(\fpu_add_frac_dp/n2306 ), .IN2(n3793), .IN3(n2638), 
        .IN4(n6), .IN5(n660), .Q(n2020) );
  INVX0 U3448 ( .INP(n2012), .ZN(n2005) );
  NAND3X0 U3449 ( .IN1(n3928), .IN2(n3917), .IN3(\fpu_add_frac_dp/n774 ), .QN(
        n2012) );
  NAND2X0 U3450 ( .IN1(n218), .IN2(n2638), .QN(n3917) );
  NAND2X0 U3451 ( .IN1(\fpu_add_frac_dp/n2306 ), .IN2(n3792), .QN(n3928) );
  AOI221X1 U3452 ( .IN1(\fpu_add_frac_dp/n2306 ), .IN2(n3794), .IN3(n2638), 
        .IN4(n23), .IN5(n655), .QN(n2015) );
  OA21X1 U3453 ( .IN1(\fpu_add_frac_dp/n579 ), .IN2(\fpu_add_frac_dp/n736 ), 
        .IN3(\fpu_add_frac_dp/n767 ), .Q(n2038) );
  NAND4X0 U3454 ( .IN1(n3929), .IN2(n3930), .IN3(n3931), .IN4(n3932), .QN(
        n2008) );
  NOR4X0 U3455 ( .IN1(n3933), .IN2(n627), .IN3(n75), .IN4(n161), .QN(n3932) );
  NAND4X0 U3456 ( .IN1(\fpu_add_frac_dp/n773 ), .IN2(\fpu_add_frac_dp/n772 ), 
        .IN3(\fpu_add_frac_dp/n767 ), .IN4(n3934), .QN(n3933) );
  NAND2X0 U3457 ( .IN1(\fpu_add_frac_dp/n2306 ), .IN2(n3935), .QN(n3934) );
  OR3X1 U3458 ( .IN1(n70), .IN2(\fpu_add_frac_dp/n2380 ), .IN3(n174), .Q(n3935) );
  NOR4X0 U3459 ( .IN1(n3936), .IN2(n312), .IN3(n106), .IN4(n720), .QN(n3931)
         );
  NAND4X0 U3460 ( .IN1(\fpu_add_frac_dp/n745 ), .IN2(\fpu_add_frac_dp/n744 ), 
        .IN3(\fpu_add_frac_dp/n743 ), .IN4(n3913), .QN(n3936) );
  AND4X1 U3461 ( .IN1(\fpu_add_frac_dp/n771 ), .IN2(\fpu_add_frac_dp/n769 ), 
        .IN3(\fpu_add_frac_dp/n766 ), .IN4(n3937), .Q(n3913) );
  AND3X1 U3462 ( .IN1(\fpu_add_frac_dp/n768 ), .IN2(\fpu_add_frac_dp/n774 ), 
        .IN3(\fpu_add_frac_dp/n770 ), .Q(n3937) );
  NOR4X0 U3463 ( .IN1(n3938), .IN2(n717), .IN3(n131), .IN4(n314), .QN(n3930)
         );
  NAND4X0 U3464 ( .IN1(\fpu_add_frac_dp/n752 ), .IN2(\fpu_add_frac_dp/n751 ), 
        .IN3(\fpu_add_frac_dp/n750 ), .IN4(\fpu_add_frac_dp/n749 ), .QN(n3938)
         );
  NOR4X0 U3465 ( .IN1(n3939), .IN2(n150), .IN3(n425), .IN4(n721), .QN(n3929)
         );
  NAND4X0 U3466 ( .IN1(\fpu_add_frac_dp/n759 ), .IN2(\fpu_add_frac_dp/n758 ), 
        .IN3(\fpu_add_frac_dp/n757 ), .IN4(\fpu_add_frac_dp/n756 ), .QN(n3939)
         );
  AO221X1 U3467 ( .IN1(n3940), .IN2(n2021), .IN3(n3941), .IN4(n755), .IN5(
        n3942), .Q(n3911) );
  AO22X1 U3468 ( .IN1(\fpu_add_frac_dp/n2306 ), .IN2(n2042), .IN3(n3943), 
        .IN4(n693), .Q(n3942) );
  NAND4X0 U3469 ( .IN1(n1998), .IN2(n3944), .IN3(n2024), .IN4(n3945), .QN(
        n3943) );
  OA221X1 U3470 ( .IN1(\fpu_add_frac_dp/n2308 ), .IN2(n3946), .IN3(
        \fpu_add_frac_dp/n580 ), .IN4(n3947), .IN5(n3948), .Q(n3945) );
  OA22X1 U3471 ( .IN1(n3949), .IN2(n2016), .IN3(n3950), .IN4(n2006), .Q(n3948)
         );
  INVX0 U3472 ( .INP(n2021), .ZN(n2006) );
  INVX0 U3473 ( .INP(n1944), .ZN(n3947) );
  NAND3X0 U3474 ( .IN1(n3949), .IN2(n3946), .IN3(n3950), .QN(n1944) );
  INVX0 U3475 ( .INP(n3896), .ZN(n3950) );
  INVX0 U3476 ( .INP(n3882), .ZN(n3949) );
  INVX0 U3477 ( .INP(n3890), .ZN(n3946) );
  AO22X1 U3478 ( .IN1(n3951), .IN2(\fpu_add_frac_dp/n2393 ), .IN3(n3790), 
        .IN4(n3884), .Q(n3890) );
  INVX0 U3479 ( .INP(n2039), .ZN(n3790) );
  OA22X1 U3480 ( .IN1(\fpu_add_frac_dp/n756 ), .IN2(\fpu_add_frac_dp/n528 ), 
        .IN3(\fpu_add_frac_dp/n572 ), .IN4(\fpu_add_frac_dp/n2395 ), .Q(n2039)
         );
  INVX0 U3481 ( .INP(n1989), .ZN(n3944) );
  NOR4X0 U3482 ( .IN1(n3952), .IN2(n2026), .IN3(n2027), .IN4(n3904), .QN(n1998) );
  AO22X1 U3483 ( .IN1(n3951), .IN2(n218), .IN3(n3792), .IN4(n3884), .Q(n3904)
         );
  AO22X1 U3484 ( .IN1(n20), .IN2(n930), .IN3(n96), .IN4(n5), .Q(n3792) );
  NAND4X0 U3485 ( .IN1(n3953), .IN2(n3954), .IN3(n3955), .IN4(n3956), .QN(
        n2042) );
  NOR4X0 U3486 ( .IN1(n75), .IN2(n161), .IN3(n627), .IN4(n3957), .QN(n3956) );
  NAND3X0 U3487 ( .IN1(n3958), .IN2(n2024), .IN3(n3959), .QN(n3941) );
  AOI222X1 U3488 ( .IN1(n2021), .IN2(n3880), .IN3(n3870), .IN4(n2028), .IN5(
        n255), .IN6(n3875), .QN(n3959) );
  AO22X1 U3489 ( .IN1(n1989), .IN2(n580), .IN3(n1993), .IN4(n581), .Q(n3875)
         );
  AO22X1 U3490 ( .IN1(n3951), .IN2(n23), .IN3(n3794), .IN4(n3884), .Q(n1993)
         );
  AO22X1 U3491 ( .IN1(n20), .IN2(n934), .IN3(n97), .IN4(n5), .Q(n3794) );
  AO222X1 U3492 ( .IN1(n3960), .IN2(n3884), .IN3(n3961), .IN4(n16), .IN5(n3951), .IN6(n678), .Q(n1989) );
  INVX0 U3493 ( .INP(n3953), .ZN(n3960) );
  OA22X1 U3494 ( .IN1(\fpu_add_frac_dp/n760 ), .IN2(\fpu_add_frac_dp/n528 ), 
        .IN3(\fpu_add_frac_dp/n572 ), .IN4(\fpu_add_frac_dp/n2517 ), .Q(n3953)
         );
  INVX0 U3495 ( .INP(n2016), .ZN(n2028) );
  AO22X1 U3496 ( .IN1(n3952), .IN2(n580), .IN3(n1991), .IN4(n581), .Q(n3870)
         );
  AO22X1 U3497 ( .IN1(n3951), .IN2(n271), .IN3(n3926), .IN4(n3884), .Q(n1991)
         );
  AND3X1 U3498 ( .IN1(n2031), .IN2(n3962), .IN3(n2030), .Q(n2024) );
  INVX0 U3499 ( .INP(n3566), .ZN(n3958) );
  AO22X1 U3500 ( .IN1(n1992), .IN2(n581), .IN3(n2027), .IN4(n580), .Q(n3566)
         );
  AO222X1 U3501 ( .IN1(n3963), .IN2(n3884), .IN3(n3961), .IN4(n156), .IN5(
        n3951), .IN6(n106), .Q(n2027) );
  INVX0 U3502 ( .INP(n3954), .ZN(n3963) );
  OA22X1 U3503 ( .IN1(\fpu_add_frac_dp/n762 ), .IN2(\fpu_add_frac_dp/n528 ), 
        .IN3(\fpu_add_frac_dp/n572 ), .IN4(\fpu_add_frac_dp/n2515 ), .Q(n3954)
         );
  AO22X1 U3504 ( .IN1(n3951), .IN2(n6), .IN3(n3793), .IN4(n3884), .Q(n1992) );
  AO22X1 U3505 ( .IN1(n314), .IN2(n20), .IN3(n5), .IN4(n95), .Q(n3793) );
  NAND2X0 U3506 ( .IN1(\fpu_add_frac_dp/n2448 ), .IN2(\fpu_add_frac_dp/n2308 ), 
        .QN(n2021) );
  OAI221X1 U3507 ( .IN1(n2016), .IN2(n3962), .IN3(n2030), .IN4(
        \fpu_add_frac_dp/n2308 ), .IN5(n2031), .QN(n3940) );
  AOI221X1 U3508 ( .IN1(\fpu_add_frac_dp/n2380 ), .IN2(n2638), .IN3(
        \fpu_add_frac_dp/n2306 ), .IN4(n3897), .IN5(n75), .QN(n2031) );
  AOI221X1 U3509 ( .IN1(n2638), .IN2(n70), .IN3(\fpu_add_frac_dp/n2306 ), 
        .IN4(n3891), .IN5(n161), .QN(n2030) );
  AO22X1 U3510 ( .IN1(n118), .IN2(n312), .IN3(n1857), .IN4(n47), .Q(n3891) );
  INVX0 U3511 ( .INP(\fpu_add_frac_dp/n2281 ), .ZN(n1857) );
  INVX0 U3512 ( .INP(\fpu_add_frac_dp/n579 ), .ZN(n2638) );
  OA221X1 U3513 ( .IN1(n624), .IN2(n3885), .IN3(\fpu_add_frac_dp/n2480 ), 
        .IN4(\fpu_add_frac_dp/n579 ), .IN5(\fpu_add_frac_dp/n763 ), .Q(n3962)
         );
  NAND2X0 U3514 ( .IN1(n962), .IN2(n255), .QN(n2016) );
  NAND3X0 U3515 ( .IN1(n3749), .IN2(n3752), .IN3(\fpu_add_frac_dp/n2385 ), 
        .QN(n3555) );
  AND2X1 U3516 ( .IN1(n3964), .IN2(n1314), .Q(n3752) );
  AO22X1 U3517 ( .IN1(n3753), .IN2(n1076), .IN3(n3754), .IN4(n569), .Q(n3964)
         );
  XOR2X1 U3518 ( .IN1(n694), .IN2(n3965), .Q(n3749) );
  OA22X1 U3519 ( .IN1(n3966), .IN2(n316), .IN3(n629), .IN4(n3967), .Q(n3965)
         );
  NOR2X0 U3520 ( .IN1(n3968), .IN2(\fpu_add_exp_dp/n111 ), .QN(n3966) );
  AOI221X1 U3521 ( .IN1(n3567), .IN2(n3572), .IN3(n3560), .IN4(n3573), .IN5(
        n3969), .QN(n3551) );
  AO22X1 U3522 ( .IN1(n3565), .IN2(n3880), .IN3(n3562), .IN4(n3575), .Q(n3969)
         );
  AO22X1 U3523 ( .IN1(n3882), .IN2(n581), .IN3(n1990), .IN4(n580), .Q(n3575)
         );
  OAI22X1 U3524 ( .IN1(\fpu_add_frac_dp/n575 ), .IN2(n3885), .IN3(
        \fpu_add_frac_dp/n2382 ), .IN4(n3970), .QN(n1990) );
  OA22X1 U3525 ( .IN1(\fpu_add_frac_dp/n572 ), .IN2(\fpu_add_frac_dp/n2480 ), 
        .IN3(\fpu_add_frac_dp/n763 ), .IN4(\fpu_add_frac_dp/n528 ), .Q(n3970)
         );
  OA22X1 U3526 ( .IN1(\fpu_add_frac_dp/n747 ), .IN2(\fpu_add_frac_dp/n545 ), 
        .IN3(\fpu_add_frac_dp/n573 ), .IN4(\fpu_add_frac_dp/n2269 ), .Q(n3885)
         );
  AO22X1 U3527 ( .IN1(n3951), .IN2(n205), .IN3(n3798), .IN4(n3884), .Q(n3882)
         );
  INVX0 U3528 ( .INP(n3923), .ZN(n3798) );
  OA22X1 U3529 ( .IN1(\fpu_add_frac_dp/n528 ), .IN2(\fpu_add_frac_dp/n755 ), 
        .IN3(\fpu_add_frac_dp/n2341 ), .IN4(\fpu_add_frac_dp/n572 ), .Q(n3923)
         );
  NOR2X0 U3530 ( .IN1(n311), .IN2(\fpu_add_frac_dp/n583 ), .QN(n3562) );
  AO22X1 U3531 ( .IN1(n1997), .IN2(n581), .IN3(n2026), .IN4(n580), .Q(n3880)
         );
  AO222X1 U3532 ( .IN1(n3971), .IN2(n3884), .IN3(n3961), .IN4(n3), .IN5(n3951), 
        .IN6(n679), .Q(n2026) );
  INVX0 U3533 ( .INP(n3955), .ZN(n3971) );
  OA22X1 U3534 ( .IN1(\fpu_add_frac_dp/n761 ), .IN2(\fpu_add_frac_dp/n528 ), 
        .IN3(\fpu_add_frac_dp/n572 ), .IN4(\fpu_add_frac_dp/n2516 ), .Q(n3955)
         );
  AO22X1 U3535 ( .IN1(n3951), .IN2(n162), .IN3(n3797), .IN4(n3884), .Q(n1997)
         );
  AO22X1 U3536 ( .IN1(n20), .IN2(n131), .IN3(n613), .IN4(n5), .Q(n3797) );
  NOR2X0 U3537 ( .IN1(\fpu_add_frac_dp/n583 ), .IN2(\fpu_add_frac_dp/n584 ), 
        .QN(n3565) );
  AO22X1 U3538 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n3952), .IN3(n1995), 
        .IN4(n580), .Q(n3573) );
  AO222X1 U3539 ( .IN1(n3789), .IN2(n901), .IN3(n3926), .IN4(n2653), .IN5(
        n3791), .IN6(n271), .Q(n1995) );
  AO22X1 U3540 ( .IN1(n20), .IN2(n931), .IN3(n98), .IN4(n5), .Q(n3926) );
  AO222X1 U3541 ( .IN1(n3951), .IN2(n696), .IN3(n3961), .IN4(n15), .IN5(n3957), 
        .IN6(n3884), .Q(n3952) );
  AO22X1 U3542 ( .IN1(n20), .IN2(n935), .IN3(n217), .IN4(n5), .Q(n3957) );
  NOR2X0 U3543 ( .IN1(\fpu_add_frac_dp/n573 ), .IN2(\fpu_add_frac_dp/n575 ), 
        .QN(n3961) );
  NOR2X0 U3544 ( .IN1(n653), .IN2(n311), .QN(n3560) );
  AO22X1 U3545 ( .IN1(\fpu_add_frac_dp/n2397 ), .IN2(n3896), .IN3(n1996), 
        .IN4(n580), .Q(n3572) );
  AO222X1 U3546 ( .IN1(n3789), .IN2(n75), .IN3(n3897), .IN4(n2653), .IN5(n3791), .IN6(\fpu_add_frac_dp/n2380 ), .Q(n1996) );
  NOR2X0 U3547 ( .IN1(\fpu_add_frac_dp/n2382 ), .IN2(\fpu_add_frac_dp/n571 ), 
        .QN(n3791) );
  INVX0 U3548 ( .INP(\fpu_add_frac_dp/n574 ), .ZN(n2653) );
  AO22X1 U3549 ( .IN1(n118), .IN2(n932), .IN3(n157), .IN4(n47), .Q(n3897) );
  NOR2X0 U3550 ( .IN1(\fpu_add_frac_dp/n2382 ), .IN2(\fpu_add_frac_dp/n513 ), 
        .QN(n3789) );
  AO22X1 U3551 ( .IN1(n3951), .IN2(n278), .IN3(n3799), .IN4(n3884), .Q(n3896)
         );
  INVX0 U3552 ( .INP(\fpu_add_frac_dp/n2382 ), .ZN(n3884) );
  INVX0 U3553 ( .INP(n2040), .ZN(n3799) );
  OA22X1 U3554 ( .IN1(\fpu_add_frac_dp/n757 ), .IN2(\fpu_add_frac_dp/n528 ), 
        .IN3(\fpu_add_frac_dp/n572 ), .IN4(\fpu_add_frac_dp/n2426 ), .Q(n2040)
         );
  NOR2X0 U3555 ( .IN1(\fpu_add_frac_dp/n545 ), .IN2(\fpu_add_frac_dp/n575 ), 
        .QN(n3951) );
  NOR2X0 U3556 ( .IN1(n653), .IN2(\fpu_add_frac_dp/n584 ), .QN(n3567) );
  NAND2X0 U3557 ( .IN1(\fpu_add_ctl/n313 ), .IN2(n1449), .QN(n1933) );
  INVX0 U3558 ( .INP(n1745), .ZN(n1746) );
  NAND2X0 U3559 ( .IN1(n3972), .IN2(n1311), .QN(n1745) );
  AO21X1 U3560 ( .IN1(n754), .IN2(n3972), .IN3(n1389), .Q(n3549) );
  NAND2X0 U3561 ( .IN1(n3973), .IN2(n3972), .QN(n2046) );
  NAND2X0 U3562 ( .IN1(fadd_clken_l), .IN2(n3972), .QN(
        \fpu_add_frac_dp/ckbuf_add_frac_dp/N1 ) );
  INVX0 U3563 ( .INP(se_add_frac), .ZN(n3972) );
  XOR3X1 U3564 ( .IN1(\fpu_add_frac_dp/n735 ), .IN2(\fpu_add_frac_dp/n598 ), 
        .IN3(n139), .Q(\fpu_add_frac_dp/a3stg_fracadd[0] ) );
  AO21X1 U3565 ( .IN1(n1455), .IN2(n1033), .IN3(n3974), .Q(
        \fpu_add_exp_dp/n722 ) );
  AO21X1 U3566 ( .IN1(n1451), .IN2(n1066), .IN3(n3975), .Q(
        \fpu_add_exp_dp/n721 ) );
  AO21X1 U3567 ( .IN1(n1451), .IN2(n1223), .IN3(n3976), .Q(
        \fpu_add_exp_dp/n720 ) );
  AO21X1 U3568 ( .IN1(n1451), .IN2(n60), .IN3(n3977), .Q(\fpu_add_exp_dp/n719 ) );
  AO21X1 U3569 ( .IN1(n1451), .IN2(n152), .IN3(n3978), .Q(
        \fpu_add_exp_dp/n718 ) );
  AO21X1 U3570 ( .IN1(n1451), .IN2(n1161), .IN3(n3979), .Q(
        \fpu_add_exp_dp/n717 ) );
  AO21X1 U3571 ( .IN1(n1451), .IN2(n1162), .IN3(n3980), .Q(
        \fpu_add_exp_dp/n716 ) );
  AO21X1 U3572 ( .IN1(n1451), .IN2(n1172), .IN3(n3981), .Q(
        \fpu_add_exp_dp/n715 ) );
  AO21X1 U3573 ( .IN1(n1451), .IN2(n1182), .IN3(n3982), .Q(
        \fpu_add_exp_dp/n714 ) );
  AO21X1 U3574 ( .IN1(n1452), .IN2(n1183), .IN3(n3983), .Q(
        \fpu_add_exp_dp/n713 ) );
  AO21X1 U3575 ( .IN1(n1451), .IN2(n1156), .IN3(n3984), .Q(
        \fpu_add_exp_dp/n712 ) );
  AO21X1 U3576 ( .IN1(n1452), .IN2(n509), .IN3(n3974), .Q(
        \fpu_add_exp_dp/n711 ) );
  AO21X1 U3577 ( .IN1(n1451), .IN2(n507), .IN3(n3975), .Q(
        \fpu_add_exp_dp/n710 ) );
  AO21X1 U3578 ( .IN1(n1452), .IN2(n508), .IN3(n3976), .Q(
        \fpu_add_exp_dp/n709 ) );
  AO21X1 U3579 ( .IN1(n1452), .IN2(n672), .IN3(n3977), .Q(
        \fpu_add_exp_dp/n708 ) );
  AO21X1 U3580 ( .IN1(n1452), .IN2(n674), .IN3(n3978), .Q(
        \fpu_add_exp_dp/n707 ) );
  AO21X1 U3581 ( .IN1(n1452), .IN2(n675), .IN3(n3979), .Q(
        \fpu_add_exp_dp/n706 ) );
  AO21X1 U3582 ( .IN1(n1452), .IN2(n668), .IN3(n3980), .Q(
        \fpu_add_exp_dp/n705 ) );
  AO21X1 U3583 ( .IN1(n1452), .IN2(n669), .IN3(n3981), .Q(
        \fpu_add_exp_dp/n704 ) );
  AO21X1 U3584 ( .IN1(n1452), .IN2(n658), .IN3(n3982), .Q(
        \fpu_add_exp_dp/n703 ) );
  AO21X1 U3585 ( .IN1(n1452), .IN2(n656), .IN3(n3983), .Q(
        \fpu_add_exp_dp/n702 ) );
  AO21X1 U3586 ( .IN1(n1452), .IN2(n657), .IN3(n3984), .Q(
        \fpu_add_exp_dp/n701 ) );
  AO22X1 U3587 ( .IN1(n1460), .IN2(n990), .IN3(n3985), .IN4(inq_in2[52]), .Q(
        \fpu_add_exp_dp/n700 ) );
  AO22X1 U3588 ( .IN1(n1460), .IN2(n991), .IN3(n3985), .IN4(inq_in2[53]), .Q(
        \fpu_add_exp_dp/n699 ) );
  AO22X1 U3589 ( .IN1(n1460), .IN2(n1005), .IN3(n3985), .IN4(inq_in2[54]), .Q(
        \fpu_add_exp_dp/n698 ) );
  AO22X1 U3590 ( .IN1(n1460), .IN2(n109), .IN3(n3985), .IN4(inq_in2[55]), .Q(
        \fpu_add_exp_dp/n697 ) );
  AO22X1 U3591 ( .IN1(n1460), .IN2(n110), .IN3(n3985), .IN4(inq_in2[56]), .Q(
        \fpu_add_exp_dp/n696 ) );
  AO22X1 U3592 ( .IN1(n1460), .IN2(n49), .IN3(n3985), .IN4(inq_in2[57]), .Q(
        \fpu_add_exp_dp/n695 ) );
  AO22X1 U3593 ( .IN1(n1460), .IN2(n42), .IN3(n3985), .IN4(inq_in2[58]), .Q(
        \fpu_add_exp_dp/n694 ) );
  AO22X1 U3594 ( .IN1(n1459), .IN2(n41), .IN3(n3985), .IN4(inq_in2[59]), .Q(
        \fpu_add_exp_dp/n693 ) );
  AO22X1 U3595 ( .IN1(n1460), .IN2(n126), .IN3(n3985), .IN4(inq_in2[60]), .Q(
        \fpu_add_exp_dp/n692 ) );
  AO22X1 U3596 ( .IN1(n1460), .IN2(n127), .IN3(n3985), .IN4(inq_in2[61]), .Q(
        \fpu_add_exp_dp/n691 ) );
  AO22X1 U3597 ( .IN1(n1460), .IN2(n105), .IN3(n3985), .IN4(inq_in2[62]), .Q(
        \fpu_add_exp_dp/n690 ) );
  OAI22X1 U3598 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n222 ), .IN3(n3987), .IN4(
        n3988), .QN(\fpu_add_exp_dp/n689 ) );
  OAI22X1 U3599 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n221 ), .IN3(n3987), .IN4(
        n3989), .QN(\fpu_add_exp_dp/n688 ) );
  OAI22X1 U3600 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n220 ), .IN3(n3987), .IN4(
        n3990), .QN(\fpu_add_exp_dp/n687 ) );
  OAI22X1 U3601 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n219 ), .IN3(n3987), .IN4(
        n3991), .QN(\fpu_add_exp_dp/n686 ) );
  OAI22X1 U3602 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n218 ), .IN3(n3987), .IN4(
        n3992), .QN(\fpu_add_exp_dp/n685 ) );
  OAI22X1 U3603 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n217 ), .IN3(n3987), .IN4(
        n3993), .QN(\fpu_add_exp_dp/n684 ) );
  OAI22X1 U3604 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n216 ), .IN3(n3987), .IN4(
        n3994), .QN(\fpu_add_exp_dp/n683 ) );
  OAI22X1 U3605 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n215 ), .IN3(n3987), .IN4(
        n3995), .QN(\fpu_add_exp_dp/n682 ) );
  AO22X1 U3606 ( .IN1(n1459), .IN2(n1180), .IN3(n3985), .IN4(inq_in2[60]), .Q(
        \fpu_add_exp_dp/n681 ) );
  AO22X1 U3607 ( .IN1(n1460), .IN2(n1075), .IN3(n3985), .IN4(inq_in2[61]), .Q(
        \fpu_add_exp_dp/n680 ) );
  AO22X1 U3608 ( .IN1(n1459), .IN2(n1181), .IN3(n3985), .IN4(inq_in2[62]), .Q(
        \fpu_add_exp_dp/n679 ) );
  AO21X1 U3609 ( .IN1(n1452), .IN2(n1159), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n678 ) );
  AO21X1 U3610 ( .IN1(n1452), .IN2(n1169), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n677 ) );
  AO21X1 U3611 ( .IN1(n1453), .IN2(n1160), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n676 ) );
  AO21X1 U3612 ( .IN1(n1453), .IN2(n958), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n675 ) );
  AO21X1 U3613 ( .IN1(n1453), .IN2(n959), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n674 ) );
  AO21X1 U3614 ( .IN1(n1453), .IN2(n960), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n673 ) );
  AO21X1 U3615 ( .IN1(n1453), .IN2(n937), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n672 ) );
  AO21X1 U3616 ( .IN1(n1453), .IN2(n936), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n671 ) );
  AO21X1 U3617 ( .IN1(n1453), .IN2(n510), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n670 ) );
  AO21X1 U3618 ( .IN1(n1453), .IN2(n61), .IN3(n3996), .Q(\fpu_add_exp_dp/n669 ) );
  AO21X1 U3619 ( .IN1(n1453), .IN2(n1174), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n668 ) );
  AO21X1 U3620 ( .IN1(n1453), .IN2(n1175), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n667 ) );
  AO21X1 U3621 ( .IN1(n1454), .IN2(n1176), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n666 ) );
  AO21X1 U3622 ( .IN1(n1453), .IN2(n1170), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n665 ) );
  AO21X1 U3623 ( .IN1(n1453), .IN2(n1177), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n664 ) );
  AO21X1 U3624 ( .IN1(n1454), .IN2(n1178), .IN3(n3996), .Q(
        \fpu_add_exp_dp/n663 ) );
  AND2X1 U3625 ( .IN1(inq_op[0]), .IN2(n3985), .Q(n3996) );
  AO21X1 U3626 ( .IN1(n1453), .IN2(n1164), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n662 ) );
  AO21X1 U3627 ( .IN1(n1454), .IN2(n1154), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n661 ) );
  AO21X1 U3628 ( .IN1(n1454), .IN2(n1165), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n660 ) );
  AO21X1 U3629 ( .IN1(n1454), .IN2(n514), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n659 ) );
  AO21X1 U3630 ( .IN1(n1454), .IN2(n515), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n658 ) );
  AO21X1 U3631 ( .IN1(n1454), .IN2(n516), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n657 ) );
  AO21X1 U3632 ( .IN1(n1454), .IN2(n546), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n656 ) );
  AO21X1 U3633 ( .IN1(n1454), .IN2(n545), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n655 ) );
  AO21X1 U3634 ( .IN1(n1454), .IN2(n1147), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n654 ) );
  AO21X1 U3635 ( .IN1(n1454), .IN2(n1150), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n653 ) );
  AO21X1 U3636 ( .IN1(n1454), .IN2(n928), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n652 ) );
  AO21X1 U3637 ( .IN1(n1454), .IN2(n151), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n651 ) );
  AO21X1 U3638 ( .IN1(n1455), .IN2(n558), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n650 ) );
  AO21X1 U3639 ( .IN1(n1455), .IN2(n1179), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n649 ) );
  AO21X1 U3640 ( .IN1(n1455), .IN2(n1166), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n648 ) );
  AO21X1 U3641 ( .IN1(n1455), .IN2(n1167), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n647 ) );
  AO21X1 U3642 ( .IN1(n1455), .IN2(n1155), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n646 ) );
  AO21X1 U3643 ( .IN1(n1455), .IN2(n1168), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n645 ) );
  AO21X1 U3644 ( .IN1(n1455), .IN2(n1171), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n644 ) );
  AO21X1 U3645 ( .IN1(n1455), .IN2(n1163), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n643 ) );
  AO21X1 U3646 ( .IN1(n1455), .IN2(n559), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n642 ) );
  AO21X1 U3647 ( .IN1(n1455), .IN2(n1148), .IN3(n3997), .Q(
        \fpu_add_exp_dp/n641 ) );
  AND2X1 U3648 ( .IN1(inq_op[1]), .IN2(n3985), .Q(n3997) );
  AO21X1 U3649 ( .IN1(n1455), .IN2(n13), .IN3(n3998), .Q(\fpu_add_exp_dp/n640 ) );
  AO21X1 U3650 ( .IN1(n1455), .IN2(n1239), .IN3(n3998), .Q(
        \fpu_add_exp_dp/n639 ) );
  AO21X1 U3651 ( .IN1(n1456), .IN2(n1240), .IN3(n3998), .Q(
        \fpu_add_exp_dp/n638 ) );
  AO21X1 U3652 ( .IN1(n1456), .IN2(n1241), .IN3(n3998), .Q(
        \fpu_add_exp_dp/n637 ) );
  AND2X1 U3653 ( .IN1(inq_op[7]), .IN2(n3985), .Q(n3998) );
  AO21X1 U3654 ( .IN1(n1456), .IN2(n992), .IN3(n3974), .Q(
        \fpu_add_exp_dp/n636 ) );
  AND2X1 U3655 ( .IN1(n3985), .IN2(inq_in1[52]), .Q(n3974) );
  AO21X1 U3656 ( .IN1(n1456), .IN2(n138), .IN3(n3975), .Q(
        \fpu_add_exp_dp/n635 ) );
  AND2X1 U3657 ( .IN1(n3985), .IN2(inq_in1[53]), .Q(n3975) );
  AO21X1 U3658 ( .IN1(n1456), .IN2(n993), .IN3(n3976), .Q(
        \fpu_add_exp_dp/n634 ) );
  AND2X1 U3659 ( .IN1(n3985), .IN2(inq_in1[54]), .Q(n3976) );
  AO21X1 U3660 ( .IN1(n1456), .IN2(n994), .IN3(n3977), .Q(
        \fpu_add_exp_dp/n633 ) );
  AND2X1 U3661 ( .IN1(n3985), .IN2(inq_in1[55]), .Q(n3977) );
  AO21X1 U3662 ( .IN1(n1456), .IN2(n995), .IN3(n3978), .Q(
        \fpu_add_exp_dp/n632 ) );
  AND2X1 U3663 ( .IN1(n3985), .IN2(inq_in1[56]), .Q(n3978) );
  AO21X1 U3664 ( .IN1(n1456), .IN2(n996), .IN3(n3979), .Q(
        \fpu_add_exp_dp/n631 ) );
  AND2X1 U3665 ( .IN1(n3985), .IN2(inq_in1[57]), .Q(n3979) );
  AO21X1 U3666 ( .IN1(n1456), .IN2(n997), .IN3(n3980), .Q(
        \fpu_add_exp_dp/n630 ) );
  AND2X1 U3667 ( .IN1(n3985), .IN2(inq_in1[58]), .Q(n3980) );
  AO21X1 U3668 ( .IN1(n1456), .IN2(n998), .IN3(n3981), .Q(
        \fpu_add_exp_dp/n629 ) );
  AND2X1 U3669 ( .IN1(n3985), .IN2(inq_in1[59]), .Q(n3981) );
  AO21X1 U3670 ( .IN1(n1456), .IN2(n999), .IN3(n3982), .Q(
        \fpu_add_exp_dp/n628 ) );
  AND2X1 U3671 ( .IN1(n3985), .IN2(inq_in1[60]), .Q(n3982) );
  AO21X1 U3672 ( .IN1(n1456), .IN2(n1000), .IN3(n3983), .Q(
        \fpu_add_exp_dp/n627 ) );
  AND2X1 U3673 ( .IN1(n3985), .IN2(inq_in1[61]), .Q(n3983) );
  AO21X1 U3674 ( .IN1(n1456), .IN2(n961), .IN3(n3984), .Q(
        \fpu_add_exp_dp/n626 ) );
  AND2X1 U3675 ( .IN1(n3985), .IN2(inq_in1[62]), .Q(n3984) );
  AO221X1 U3676 ( .IN1(n3985), .IN2(n3988), .IN3(n1451), .IN4(n491), .IN5(
        n3999), .Q(\fpu_add_exp_dp/n625 ) );
  INVX0 U3677 ( .INP(inq_in2[52]), .ZN(n3988) );
  AO221X1 U3678 ( .IN1(n3985), .IN2(n3989), .IN3(n1451), .IN4(n56), .IN5(n3999), .Q(\fpu_add_exp_dp/n624 ) );
  INVX0 U3679 ( .INP(inq_in2[53]), .ZN(n3989) );
  AO221X1 U3680 ( .IN1(n3985), .IN2(n3990), .IN3(n1451), .IN4(n309), .IN5(
        n3999), .Q(\fpu_add_exp_dp/n623 ) );
  NOR2X0 U3681 ( .IN1(n3987), .IN2(inq_op[1]), .QN(n3999) );
  INVX0 U3682 ( .INP(inq_in2[54]), .ZN(n3990) );
  AO22X1 U3683 ( .IN1(n1459), .IN2(n319), .IN3(n3985), .IN4(n3991), .Q(
        \fpu_add_exp_dp/n622 ) );
  INVX0 U3684 ( .INP(inq_in2[55]), .ZN(n3991) );
  AO22X1 U3685 ( .IN1(n1460), .IN2(n320), .IN3(n3985), .IN4(n3992), .Q(
        \fpu_add_exp_dp/n621 ) );
  INVX0 U3686 ( .INP(inq_in2[56]), .ZN(n3992) );
  AO22X1 U3687 ( .IN1(n1459), .IN2(n321), .IN3(n3985), .IN4(n3993), .Q(
        \fpu_add_exp_dp/n620 ) );
  INVX0 U3688 ( .INP(inq_in2[57]), .ZN(n3993) );
  AO22X1 U3689 ( .IN1(n1460), .IN2(n322), .IN3(n3985), .IN4(n3994), .Q(
        \fpu_add_exp_dp/n619 ) );
  INVX0 U3690 ( .INP(inq_in2[58]), .ZN(n3994) );
  AO22X1 U3691 ( .IN1(n1459), .IN2(n323), .IN3(n3985), .IN4(n3995), .Q(
        \fpu_add_exp_dp/n618 ) );
  INVX0 U3692 ( .INP(inq_in2[59]), .ZN(n3995) );
  INVX0 U3693 ( .INP(n3987), .ZN(n3985) );
  OAI22X1 U3694 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n150 ), .IN3(n3987), .IN4(
        inq_in2[60]), .QN(\fpu_add_exp_dp/n617 ) );
  OAI22X1 U3695 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n149 ), .IN3(n3987), .IN4(
        inq_in2[61]), .QN(\fpu_add_exp_dp/n616 ) );
  OAI22X1 U3696 ( .IN1(n3986), .IN2(\fpu_add_exp_dp/n47 ), .IN3(n3987), .IN4(
        inq_in2[62]), .QN(\fpu_add_exp_dp/n615 ) );
  NAND2X0 U3697 ( .IN1(a1stg_step), .IN2(\fpu_add_ctl/n470 ), .QN(n3987) );
  AO21X1 U3698 ( .IN1(n1467), .IN2(n645), .IN3(n4001), .Q(
        \fpu_add_exp_dp/n614 ) );
  AO21X1 U3699 ( .IN1(n1465), .IN2(n73), .IN3(n4002), .Q(\fpu_add_exp_dp/n613 ) );
  AO21X1 U3700 ( .IN1(n1464), .IN2(n287), .IN3(n4003), .Q(
        \fpu_add_exp_dp/n612 ) );
  AO21X1 U3701 ( .IN1(n1464), .IN2(n290), .IN3(n4004), .Q(
        \fpu_add_exp_dp/n611 ) );
  AO21X1 U3702 ( .IN1(n1465), .IN2(n648), .IN3(n4005), .Q(
        \fpu_add_exp_dp/n610 ) );
  AO21X1 U3703 ( .IN1(n1464), .IN2(n646), .IN3(n4006), .Q(
        \fpu_add_exp_dp/n609 ) );
  AO21X1 U3704 ( .IN1(n1467), .IN2(n711), .IN3(n4007), .Q(
        \fpu_add_exp_dp/n608 ) );
  AO21X1 U3705 ( .IN1(n1466), .IN2(n221), .IN3(n4008), .Q(
        \fpu_add_exp_dp/n607 ) );
  AO21X1 U3706 ( .IN1(n1464), .IN2(n35), .IN3(n4009), .Q(\fpu_add_exp_dp/n606 ) );
  AO21X1 U3707 ( .IN1(n1464), .IN2(n88), .IN3(n4010), .Q(\fpu_add_exp_dp/n605 ) );
  AO21X1 U3708 ( .IN1(n1467), .IN2(n289), .IN3(n4011), .Q(
        \fpu_add_exp_dp/n604 ) );
  AO21X1 U3709 ( .IN1(n1464), .IN2(n725), .IN3(n4012), .Q(
        \fpu_add_exp_dp/n603 ) );
  AO21X1 U3710 ( .IN1(n1464), .IN2(n315), .IN3(n4001), .Q(
        \fpu_add_exp_dp/n602 ) );
  AO22X1 U3711 ( .IN1(n4013), .IN2(n2622), .IN3(n1339), .IN4(n4014), .Q(n4001)
         );
  AO221X1 U3712 ( .IN1(n4015), .IN2(n672), .IN3(n4016), .IN4(n109), .IN5(n4017), .Q(n4014) );
  AO22X1 U3713 ( .IN1(n4018), .IN2(n990), .IN3(n4019), .IN4(n509), .Q(n4017)
         );
  AO21X1 U3714 ( .IN1(n1466), .IN2(n676), .IN3(n4002), .Q(
        \fpu_add_exp_dp/n601 ) );
  AO22X1 U3715 ( .IN1(n1338), .IN2(n4020), .IN3(n4013), .IN4(n4021), .Q(n4002)
         );
  XOR2X1 U3716 ( .IN1(n2622), .IN2(n2619), .Q(n4021) );
  AO221X1 U3717 ( .IN1(n4015), .IN2(n674), .IN3(n4016), .IN4(n110), .IN5(n4022), .Q(n4020) );
  AO22X1 U3718 ( .IN1(n4018), .IN2(n991), .IN3(n4019), .IN4(n507), .Q(n4022)
         );
  AO21X1 U3719 ( .IN1(n1467), .IN2(n687), .IN3(n4003), .Q(
        \fpu_add_exp_dp/n600 ) );
  AO22X1 U3720 ( .IN1(n2629), .IN2(n4013), .IN3(n1340), .IN4(n4023), .Q(n4003)
         );
  AO221X1 U3721 ( .IN1(n4015), .IN2(n675), .IN3(n4016), .IN4(n49), .IN5(n4024), 
        .Q(n4023) );
  AO22X1 U3722 ( .IN1(n4018), .IN2(n1005), .IN3(n4019), .IN4(n508), .Q(n4024)
         );
  OA21X1 U3723 ( .IN1(n2631), .IN2(n2623), .IN3(n4025), .Q(n2629) );
  AO21X1 U3724 ( .IN1(n1464), .IN2(n686), .IN3(n4004), .Q(
        \fpu_add_exp_dp/n599 ) );
  AO22X1 U3725 ( .IN1(n1340), .IN2(n4026), .IN3(n4027), .IN4(n4013), .Q(n4004)
         );
  NOR2X0 U3726 ( .IN1(n2651), .IN2(n2652), .QN(n4027) );
  NOR2X0 U3727 ( .IN1(n2649), .IN2(n4028), .QN(n2652) );
  AO221X1 U3728 ( .IN1(n4019), .IN2(n672), .IN3(n4018), .IN4(n109), .IN5(n4029), .Q(n4026) );
  AO22X1 U3729 ( .IN1(n4016), .IN2(n42), .IN3(n4015), .IN4(n668), .Q(n4029) );
  AO21X1 U3730 ( .IN1(n1466), .IN2(n685), .IN3(n4005), .Q(
        \fpu_add_exp_dp/n598 ) );
  AO22X1 U3731 ( .IN1(n1337), .IN2(n4030), .IN3(n4031), .IN4(n4013), .Q(n4005)
         );
  NOR2X0 U3732 ( .IN1(n2665), .IN2(n2666), .QN(n4031) );
  NOR2X0 U3733 ( .IN1(n2662), .IN2(n2651), .QN(n2666) );
  AO221X1 U3734 ( .IN1(n4019), .IN2(n674), .IN3(n4018), .IN4(n110), .IN5(n4032), .Q(n4030) );
  AO22X1 U3735 ( .IN1(n4016), .IN2(n41), .IN3(n4015), .IN4(n669), .Q(n4032) );
  AO21X1 U3736 ( .IN1(n1464), .IN2(n684), .IN3(n4006), .Q(
        \fpu_add_exp_dp/n597 ) );
  AO22X1 U3737 ( .IN1(n1339), .IN2(n4033), .IN3(n4034), .IN4(n4013), .Q(n4006)
         );
  NOR2X0 U3738 ( .IN1(n2729), .IN2(n2730), .QN(n4034) );
  NOR2X0 U3739 ( .IN1(n2718), .IN2(n2665), .QN(n2730) );
  INVX0 U3740 ( .INP(n4035), .ZN(n2665) );
  INVX0 U3741 ( .INP(n4036), .ZN(n2718) );
  AO221X1 U3742 ( .IN1(n4019), .IN2(n675), .IN3(n4018), .IN4(n49), .IN5(n4037), 
        .Q(n4033) );
  AO22X1 U3743 ( .IN1(n4016), .IN2(n126), .IN3(n4015), .IN4(n658), .Q(n4037)
         );
  AO21X1 U3744 ( .IN1(n1466), .IN2(n661), .IN3(n4007), .Q(
        \fpu_add_exp_dp/n596 ) );
  AO22X1 U3745 ( .IN1(n1338), .IN2(n4038), .IN3(n4039), .IN4(n4013), .Q(n4007)
         );
  OA21X1 U3746 ( .IN1(n2729), .IN2(n2700), .IN3(n4040), .Q(n4039) );
  AO221X1 U3747 ( .IN1(n4019), .IN2(n668), .IN3(n4018), .IN4(n42), .IN5(n4041), 
        .Q(n4038) );
  AO22X1 U3748 ( .IN1(n4016), .IN2(n127), .IN3(n4015), .IN4(n656), .Q(n4041)
         );
  AO21X1 U3749 ( .IN1(n1466), .IN2(n683), .IN3(n4008), .Q(
        \fpu_add_exp_dp/n595 ) );
  AO22X1 U3750 ( .IN1(n1340), .IN2(n4042), .IN3(n4043), .IN4(n4013), .Q(n4008)
         );
  AOI21X1 U3751 ( .IN1(n4040), .IN2(n2703), .IN3(n4044), .QN(n4043) );
  AO221X1 U3752 ( .IN1(n4019), .IN2(n669), .IN3(n4018), .IN4(n41), .IN5(n4045), 
        .Q(n4042) );
  AO22X1 U3753 ( .IN1(n4016), .IN2(n105), .IN3(n4015), .IN4(n657), .Q(n4045)
         );
  NOR2X0 U3754 ( .IN1(n4046), .IN2(n4047), .QN(n4015) );
  AO21X1 U3755 ( .IN1(a1stg_faddsubs), .IN2(n4047), .IN3(n4048), .Q(n4016) );
  AO21X1 U3756 ( .IN1(n1464), .IN2(n682), .IN3(n4009), .Q(
        \fpu_add_exp_dp/n594 ) );
  AO222X1 U3757 ( .IN1(n4049), .IN2(n126), .IN3(n4050), .IN4(n4013), .IN5(
        n4051), .IN6(n658), .Q(n4009) );
  OA21X1 U3758 ( .IN1(n2713), .IN2(n4044), .IN3(n4052), .Q(n4050) );
  AO21X1 U3759 ( .IN1(n1465), .IN2(n681), .IN3(n4010), .Q(
        \fpu_add_exp_dp/n593 ) );
  AO222X1 U3760 ( .IN1(n4049), .IN2(n127), .IN3(n4053), .IN4(n4013), .IN5(
        n4051), .IN6(n656), .Q(n4010) );
  AOI21X1 U3761 ( .IN1(n2710), .IN2(n4052), .IN3(n4054), .QN(n4053) );
  AO21X1 U3762 ( .IN1(n1465), .IN2(n680), .IN3(n4011), .Q(
        \fpu_add_exp_dp/n592 ) );
  AO222X1 U3763 ( .IN1(n4049), .IN2(n105), .IN3(n4013), .IN4(n4055), .IN5(
        n4051), .IN6(n657), .Q(n4011) );
  AND2X1 U3764 ( .IN1(n1340), .IN2(n4019), .Q(n4051) );
  NOR2X0 U3765 ( .IN1(n4047), .IN2(n4056), .QN(n4019) );
  XOR2X1 U3766 ( .IN1(n2706), .IN2(n4054), .Q(n4055) );
  AND2X1 U3767 ( .IN1(n1337), .IN2(n4018), .Q(n4049) );
  AO21X1 U3768 ( .IN1(n1658), .IN2(n4047), .IN3(a1stg_fdtos), .Q(n4018) );
  INVX0 U3769 ( .INP(n2050), .ZN(n4047) );
  AO21X1 U3770 ( .IN1(n1465), .IN2(n316), .IN3(n4012), .Q(
        \fpu_add_exp_dp/n591 ) );
  AND3X1 U3771 ( .IN1(n4013), .IN2(n2706), .IN3(n4054), .Q(n4012) );
  NOR2X0 U3772 ( .IN1(n4052), .IN2(n2710), .QN(n4054) );
  NAND2X0 U3773 ( .IN1(n559), .IN2(n1075), .QN(n2710) );
  NAND2X0 U3774 ( .IN1(n4044), .IN2(n2713), .QN(n4052) );
  NOR2X0 U3775 ( .IN1(\fpu_add_exp_dp/n176 ), .IN2(\fpu_add_exp_dp/n214 ), 
        .QN(n2713) );
  NOR2X0 U3776 ( .IN1(n4040), .IN2(n2703), .QN(n4044) );
  OA22X1 U3777 ( .IN1(\fpu_add_exp_dp/n215 ), .IN2(\fpu_add_exp_dp/n177 ), 
        .IN3(\fpu_add_exp_dp/n212 ), .IN4(\fpu_add_exp_dp/n196 ), .Q(n2703) );
  NAND2X0 U3778 ( .IN1(n2729), .IN2(n2700), .QN(n4040) );
  OAI22X1 U3779 ( .IN1(\fpu_add_exp_dp/n197 ), .IN2(\fpu_add_exp_dp/n213 ), 
        .IN3(\fpu_add_exp_dp/n178 ), .IN4(\fpu_add_exp_dp/n216 ), .QN(n2700)
         );
  NOR2X0 U3780 ( .IN1(n4035), .IN2(n4036), .QN(n2729) );
  OA22X1 U3781 ( .IN1(\fpu_add_exp_dp/n217 ), .IN2(\fpu_add_exp_dp/n179 ), 
        .IN3(\fpu_add_exp_dp/n214 ), .IN4(\fpu_add_exp_dp/n198 ), .Q(n4036) );
  NAND2X0 U3782 ( .IN1(n2651), .IN2(n2662), .QN(n4035) );
  OAI22X1 U3783 ( .IN1(\fpu_add_exp_dp/n199 ), .IN2(\fpu_add_exp_dp/n215 ), 
        .IN3(\fpu_add_exp_dp/n180 ), .IN4(\fpu_add_exp_dp/n218 ), .QN(n2662)
         );
  AND2X1 U3784 ( .IN1(n4028), .IN2(n2649), .Q(n2651) );
  OAI22X1 U3785 ( .IN1(\fpu_add_exp_dp/n200 ), .IN2(\fpu_add_exp_dp/n216 ), 
        .IN3(\fpu_add_exp_dp/n181 ), .IN4(\fpu_add_exp_dp/n219 ), .QN(n2649)
         );
  INVX0 U3786 ( .INP(n4025), .ZN(n4028) );
  NAND2X0 U3787 ( .IN1(n2623), .IN2(n2631), .QN(n4025) );
  OAI22X1 U3788 ( .IN1(\fpu_add_exp_dp/n220 ), .IN2(\fpu_add_exp_dp/n182 ), 
        .IN3(\fpu_add_exp_dp/n217 ), .IN4(\fpu_add_exp_dp/n201 ), .QN(n2631)
         );
  NOR2X0 U3789 ( .IN1(n2619), .IN2(n2622), .QN(n2623) );
  OA22X1 U3790 ( .IN1(\fpu_add_exp_dp/n222 ), .IN2(\fpu_add_exp_dp/n184 ), 
        .IN3(\fpu_add_exp_dp/n219 ), .IN4(\fpu_add_exp_dp/n203 ), .Q(n2622) );
  OA22X1 U3791 ( .IN1(\fpu_add_exp_dp/n202 ), .IN2(\fpu_add_exp_dp/n218 ), 
        .IN3(\fpu_add_exp_dp/n183 ), .IN4(\fpu_add_exp_dp/n221 ), .Q(n2619) );
  NOR2X0 U3792 ( .IN1(\fpu_add_exp_dp/n174 ), .IN2(\fpu_add_exp_dp/n212 ), 
        .QN(n2706) );
  NOR2X0 U3793 ( .IN1(n4057), .IN2(n4058), .QN(n4013) );
  AO21X1 U3794 ( .IN1(n1466), .IN2(n830), .IN3(n4059), .Q(
        \fpu_add_exp_dp/n589 ) );
  AO21X1 U3795 ( .IN1(n1465), .IN2(n297), .IN3(n4059), .Q(
        \fpu_add_exp_dp/n588 ) );
  AO21X1 U3796 ( .IN1(n1465), .IN2(n305), .IN3(n4059), .Q(
        \fpu_add_exp_dp/n587 ) );
  AO21X1 U3797 ( .IN1(n1466), .IN2(n304), .IN3(n4059), .Q(
        \fpu_add_exp_dp/n586 ) );
  AO21X1 U3798 ( .IN1(n1465), .IN2(n303), .IN3(n4059), .Q(
        \fpu_add_exp_dp/n585 ) );
  AO221X1 U3799 ( .IN1(n1462), .IN2(n299), .IN3(n4060), .IN4(n1340), .IN5(
        n4061), .Q(\fpu_add_exp_dp/n584 ) );
  AO21X1 U3800 ( .IN1(n1466), .IN2(n302), .IN3(n4062), .Q(
        \fpu_add_exp_dp/n583 ) );
  AO22X1 U3801 ( .IN1(n1472), .IN2(n308), .IN3(n1338), .IN4(n4063), .Q(
        \fpu_add_exp_dp/n582 ) );
  NAND2X0 U3802 ( .IN1(n4064), .IN2(n4065), .QN(n4063) );
  AO21X1 U3803 ( .IN1(n1465), .IN2(n301), .IN3(n4066), .Q(
        \fpu_add_exp_dp/n581 ) );
  AO21X1 U3804 ( .IN1(n1465), .IN2(n300), .IN3(n4066), .Q(
        \fpu_add_exp_dp/n580 ) );
  OA21X1 U3805 ( .IN1(n4067), .IN2(n4048), .IN3(n1338), .Q(n4066) );
  AO221X1 U3806 ( .IN1(n1462), .IN2(n298), .IN3(n4068), .IN4(n1340), .IN5(
        n4061), .Q(\fpu_add_exp_dp/n579 ) );
  AO21X1 U3807 ( .IN1(n4069), .IN2(n1340), .IN3(n4059), .Q(n4061) );
  AO21X1 U3808 ( .IN1(n1465), .IN2(n629), .IN3(n4062), .Q(
        \fpu_add_exp_dp/n578 ) );
  AO21X1 U3809 ( .IN1(n1465), .IN2(n694), .IN3(n4062), .Q(
        \fpu_add_exp_dp/n577 ) );
  AO21X1 U3810 ( .IN1(n1338), .IN2(n4067), .IN3(n4059), .Q(n4062) );
  NOR2X0 U3811 ( .IN1(n4070), .IN2(n4057), .QN(n4059) );
  OR3X1 U3812 ( .IN1(n4068), .IN2(n4069), .IN3(n4071), .Q(n4067) );
  INVX0 U3813 ( .INP(n4064), .ZN(n4071) );
  NOR2X0 U3814 ( .IN1(n4060), .IN2(n4072), .QN(n4064) );
  AO221X1 U3815 ( .IN1(n4073), .IN2(n4074), .IN3(n4075), .IN4(n315), .IN5(
        n4076), .Q(\fpu_add_exp_dp/n576 ) );
  AO21X1 U3816 ( .IN1(n1466), .IN2(n583), .IN3(n4077), .Q(n4076) );
  AO221X1 U3817 ( .IN1(n4075), .IN2(n676), .IN3(n1462), .IN4(n72), .IN5(n4078), 
        .Q(\fpu_add_exp_dp/n575 ) );
  AO21X1 U3818 ( .IN1(n4079), .IN2(n4073), .IN3(n4080), .Q(n4078) );
  INVX0 U3819 ( .INP(n4081), .ZN(n4079) );
  AO221X1 U3820 ( .IN1(n4075), .IN2(n687), .IN3(n1463), .IN4(n159), .IN5(n4082), .Q(\fpu_add_exp_dp/n574 ) );
  AO21X1 U3821 ( .IN1(n4083), .IN2(n4073), .IN3(n4080), .Q(n4082) );
  AO221X1 U3822 ( .IN1(n4075), .IN2(n686), .IN3(n1462), .IN4(n178), .IN5(n4084), .Q(\fpu_add_exp_dp/n573 ) );
  AO21X1 U3823 ( .IN1(n4085), .IN2(n4073), .IN3(n4080), .Q(n4084) );
  AO221X1 U3824 ( .IN1(n4075), .IN2(n685), .IN3(n1463), .IN4(n67), .IN5(n4086), 
        .Q(\fpu_add_exp_dp/n572 ) );
  AO21X1 U3825 ( .IN1(n4087), .IN2(n4073), .IN3(n4080), .Q(n4086) );
  AND2X1 U3826 ( .IN1(n1339), .IN2(n4088), .Q(n4080) );
  OR3X1 U3827 ( .IN1(n421), .IN2(n4089), .IN3(n718), .Q(n4088) );
  AO221X1 U3828 ( .IN1(n4075), .IN2(n684), .IN3(n1463), .IN4(n69), .IN5(n4090), 
        .Q(\fpu_add_exp_dp/n571 ) );
  AO22X1 U3829 ( .IN1(n4091), .IN2(n4073), .IN3(n1337), .IN4(n4089), .Q(n4090)
         );
  NAND2X0 U3830 ( .IN1(\fpu_add_ctl/n207 ), .IN2(n4092), .QN(n4089) );
  AO221X1 U3831 ( .IN1(n4093), .IN2(n4073), .IN3(n4075), .IN4(n661), .IN5(
        n4094), .Q(\fpu_add_exp_dp/n570 ) );
  AO21X1 U3832 ( .IN1(n1465), .IN2(n160), .IN3(n4077), .Q(n4094) );
  NAND2X0 U3833 ( .IN1(n4095), .IN2(n4096), .QN(n4077) );
  NAND3X0 U3834 ( .IN1(n1339), .IN2(n91), .IN3(n4097), .QN(n4096) );
  AO221X1 U3835 ( .IN1(n4075), .IN2(n683), .IN3(n1462), .IN4(n256), .IN5(n4098), .Q(\fpu_add_exp_dp/n569 ) );
  AO22X1 U3836 ( .IN1(n4099), .IN2(n4073), .IN3(n1339), .IN4(n4100), .Q(n4098)
         );
  NAND2X0 U3837 ( .IN1(\fpu_add_ctl/n147 ), .IN2(n4092), .QN(n4100) );
  AOI221X1 U3838 ( .IN1(n4097), .IN2(n91), .IN3(n4101), .IN4(n258), .IN5(n757), 
        .QN(n4092) );
  INVX0 U3839 ( .INP(n4102), .ZN(n4097) );
  AO221X1 U3840 ( .IN1(n4075), .IN2(n682), .IN3(n1463), .IN4(n71), .IN5(n4103), 
        .Q(\fpu_add_exp_dp/n568 ) );
  AO21X1 U3841 ( .IN1(n4104), .IN2(n4073), .IN3(n4105), .Q(n4103) );
  AO221X1 U3842 ( .IN1(n4075), .IN2(n681), .IN3(n1463), .IN4(n17), .IN5(n4106), 
        .Q(\fpu_add_exp_dp/n567 ) );
  AO21X1 U3843 ( .IN1(n4107), .IN2(n4073), .IN3(n4105), .Q(n4106) );
  AO221X1 U3844 ( .IN1(n4075), .IN2(n680), .IN3(n1462), .IN4(n181), .IN5(n4108), .Q(\fpu_add_exp_dp/n566 ) );
  AO221X1 U3845 ( .IN1(n1338), .IN2(n4109), .IN3(n4110), .IN4(n4073), .IN5(
        n4105), .Q(n4108) );
  INVX0 U3846 ( .INP(n4095), .ZN(n4105) );
  NAND3X0 U3847 ( .IN1(n1338), .IN2(n258), .IN3(n4101), .QN(n4095) );
  AND3X1 U3848 ( .IN1(n4111), .IN2(n4112), .IN3(n1340), .Q(n4073) );
  AO21X1 U3849 ( .IN1(n4102), .IN2(n91), .IN3(n258), .Q(n4112) );
  NAND4X0 U3850 ( .IN1(n4101), .IN2(n289), .IN3(n88), .IN4(n35), .QN(n4102) );
  AND4X1 U3851 ( .IN1(n1901), .IN2(n221), .IN3(n1910), .IN4(n4113), .Q(n4101)
         );
  NOR3X0 U3852 ( .IN1(\fpu_add_exp_dp/n141 ), .IN2(\fpu_add_exp_dp/n146 ), 
        .IN3(\fpu_add_exp_dp/n143 ), .QN(n4113) );
  NOR2X0 U3853 ( .IN1(\fpu_add_exp_dp/n142 ), .IN2(\fpu_add_exp_dp/n144 ), 
        .QN(n1910) );
  NAND2X0 U3854 ( .IN1(\fpu_add_ctl/n150 ), .IN2(\fpu_add_ctl/n207 ), .QN(
        n4109) );
  AO22X1 U3855 ( .IN1(n4000), .IN2(n728), .IN3(n4075), .IN4(n316), .Q(
        \fpu_add_exp_dp/n565 ) );
  OAI22X1 U3856 ( .IN1(n4057), .IN2(\fpu_add_exp_dp/n444 ), .IN3(n4114), .IN4(
        \fpu_add_exp_dp/n57 ), .QN(\fpu_add_exp_dp/n563 ) );
  AO22X1 U3857 ( .IN1(n1337), .IN2(n72), .IN3(n1469), .IN4(n643), .Q(
        \fpu_add_exp_dp/n562 ) );
  OAI22X1 U3858 ( .IN1(n4057), .IN2(\fpu_add_exp_dp/n431 ), .IN3(n4114), .IN4(
        \fpu_add_exp_dp/n438 ), .QN(\fpu_add_exp_dp/n561 ) );
  OAI22X1 U3859 ( .IN1(n4057), .IN2(\fpu_add_exp_dp/n434 ), .IN3(n4114), .IN4(
        \fpu_add_exp_dp/n439 ), .QN(\fpu_add_exp_dp/n560 ) );
  OAI22X1 U3860 ( .IN1(n4057), .IN2(\fpu_add_exp_dp/n432 ), .IN3(n4114), .IN4(
        \fpu_add_exp_dp/n440 ), .QN(\fpu_add_exp_dp/n559 ) );
  AO22X1 U3861 ( .IN1(n1339), .IN2(n69), .IN3(n1470), .IN4(n761), .Q(
        \fpu_add_exp_dp/n558 ) );
  AO22X1 U3862 ( .IN1(n1338), .IN2(n160), .IN3(n1469), .IN4(n666), .Q(
        \fpu_add_exp_dp/n557 ) );
  OAI22X1 U3863 ( .IN1(n4057), .IN2(\fpu_add_exp_dp/n442 ), .IN3(n4114), .IN4(
        \fpu_add_exp_dp/n50 ), .QN(\fpu_add_exp_dp/n556 ) );
  OAI22X1 U3864 ( .IN1(n4057), .IN2(\fpu_add_exp_dp/n445 ), .IN3(n4114), .IN4(
        \fpu_add_exp_dp/n450 ), .QN(\fpu_add_exp_dp/n555 ) );
  OAI22X1 U3865 ( .IN1(n4057), .IN2(\fpu_add_exp_dp/n443 ), .IN3(n4114), .IN4(
        \fpu_add_exp_dp/n48 ), .QN(\fpu_add_exp_dp/n554 ) );
  AO22X1 U3866 ( .IN1(n1340), .IN2(n181), .IN3(n1470), .IN4(n663), .Q(
        \fpu_add_exp_dp/n553 ) );
  OAI22X1 U3867 ( .IN1(n4057), .IN2(\fpu_add_exp_dp/n447 ), .IN3(n4114), .IN4(
        \fpu_add_exp_dp/n46 ), .QN(\fpu_add_exp_dp/n552 ) );
  AO21X1 U3868 ( .IN1(n1465), .IN2(n454), .IN3(n4115), .Q(
        \fpu_add_exp_dp/n550 ) );
  OA222X1 U3869 ( .IN1(n2959), .IN2(n2957), .IN3(n4116), .IN4(n4117), .IN5(
        n4118), .IN6(n4119), .Q(n4115) );
  AND2X1 U3870 ( .IN1(n2962), .IN2(n1339), .Q(n4116) );
  XOR2X1 U3871 ( .IN1(\fpu_add_ctl/n307 ), .IN2(n4120), .Q(n2957) );
  NOR2X0 U3872 ( .IN1(\fpu_add_ctl/n337 ), .IN2(\fpu_add_ctl/n937 ), .QN(n4120) );
  AO221X1 U3873 ( .IN1(n4121), .IN2(n4122), .IN3(n1463), .IN4(n440), .IN5(
        n4123), .Q(\fpu_add_exp_dp/n549 ) );
  NAND2X0 U3874 ( .IN1(n4124), .IN2(n4125), .QN(n4123) );
  NAND3X0 U3875 ( .IN1(n4126), .IN2(n4127), .IN3(n4128), .QN(n4124) );
  NAND2X0 U3876 ( .IN1(n4129), .IN2(n4130), .QN(n4127) );
  AO221X1 U3877 ( .IN1(n4122), .IN2(n4131), .IN3(n1462), .IN4(n439), .IN5(
        n4132), .Q(\fpu_add_exp_dp/n548 ) );
  NAND2X0 U3878 ( .IN1(n4133), .IN2(n4125), .QN(n4132) );
  NAND3X0 U3879 ( .IN1(n4126), .IN2(n4134), .IN3(n4135), .QN(n4133) );
  INVX0 U3880 ( .INP(n4136), .ZN(n4135) );
  NAND2X0 U3881 ( .IN1(n4137), .IN2(n4129), .QN(n4134) );
  INVX0 U3882 ( .INP(n4137), .ZN(n4131) );
  AO221X1 U3883 ( .IN1(n4122), .IN2(n4138), .IN3(n1463), .IN4(n438), .IN5(
        n4139), .Q(\fpu_add_exp_dp/n547 ) );
  NAND2X0 U3884 ( .IN1(n4140), .IN2(n4125), .QN(n4139) );
  NAND3X0 U3885 ( .IN1(n4126), .IN2(n4141), .IN3(n4142), .QN(n4140) );
  NAND2X0 U3886 ( .IN1(n4143), .IN2(n4129), .QN(n4141) );
  INVX0 U3887 ( .INP(n4143), .ZN(n4138) );
  AO221X1 U3888 ( .IN1(n4122), .IN2(n4144), .IN3(n1462), .IN4(n437), .IN5(
        n4145), .Q(\fpu_add_exp_dp/n546 ) );
  NAND2X0 U3889 ( .IN1(n4146), .IN2(n4125), .QN(n4145) );
  NAND3X0 U3890 ( .IN1(n4126), .IN2(n4147), .IN3(n4148), .QN(n4146) );
  NAND2X0 U3891 ( .IN1(n4149), .IN2(n4129), .QN(n4147) );
  INVX0 U3892 ( .INP(n4149), .ZN(n4144) );
  AO221X1 U3893 ( .IN1(n4122), .IN2(n4150), .IN3(n1462), .IN4(n436), .IN5(
        n4151), .Q(\fpu_add_exp_dp/n545 ) );
  NAND2X0 U3894 ( .IN1(n4152), .IN2(n4125), .QN(n4151) );
  NAND3X0 U3895 ( .IN1(n4126), .IN2(n4153), .IN3(n4154), .QN(n4152) );
  NAND2X0 U3896 ( .IN1(n4155), .IN2(n4129), .QN(n4153) );
  AO221X1 U3897 ( .IN1(n4156), .IN2(n4122), .IN3(n1462), .IN4(n435), .IN5(
        n4157), .Q(\fpu_add_exp_dp/n544 ) );
  NAND2X0 U3898 ( .IN1(n4158), .IN2(n4125), .QN(n4157) );
  NAND3X0 U3899 ( .IN1(n4126), .IN2(n4159), .IN3(n4160), .QN(n4158) );
  NAND2X0 U3900 ( .IN1(n4129), .IN2(n4161), .QN(n4159) );
  INVX0 U3901 ( .INP(n4161), .ZN(n4156) );
  AO221X1 U3902 ( .IN1(n4162), .IN2(n4122), .IN3(n1463), .IN4(n434), .IN5(
        n4163), .Q(\fpu_add_exp_dp/n543 ) );
  NAND2X0 U3903 ( .IN1(n4164), .IN2(n4125), .QN(n4163) );
  NAND2X0 U3904 ( .IN1(n4122), .IN2(n4119), .QN(n4125) );
  NAND3X0 U3905 ( .IN1(n4126), .IN2(n4165), .IN3(n4166), .QN(n4164) );
  NAND2X0 U3906 ( .IN1(n4129), .IN2(n4167), .QN(n4165) );
  INVX0 U3907 ( .INP(n4119), .ZN(n4129) );
  AND2X1 U3908 ( .IN1(n4126), .IN2(n2962), .Q(n4122) );
  AO21X1 U3909 ( .IN1(n1467), .IN2(n759), .IN3(n4168), .Q(
        \fpu_add_exp_dp/n542 ) );
  OA221X1 U3910 ( .IN1(n2962), .IN2(n4169), .IN3(n4170), .IN4(n4119), .IN5(
        n4171), .Q(n4168) );
  INVX0 U3911 ( .INP(n4172), .ZN(n4169) );
  AO21X1 U3912 ( .IN1(n1466), .IN2(n758), .IN3(n4173), .Q(
        \fpu_add_exp_dp/n541 ) );
  OA221X1 U3913 ( .IN1(n2962), .IN2(n4174), .IN3(n4175), .IN4(n4119), .IN5(
        n4171), .Q(n4173) );
  AO21X1 U3914 ( .IN1(n1466), .IN2(n760), .IN3(n4176), .Q(
        \fpu_add_exp_dp/n540 ) );
  OA221X1 U3915 ( .IN1(n2962), .IN2(n4177), .IN3(n4178), .IN4(n4119), .IN5(
        n4171), .Q(n4176) );
  AO21X1 U3916 ( .IN1(\fpu_add_ctl/n65 ), .IN2(n1338), .IN3(n4126), .Q(n4171)
         );
  AND2X1 U3917 ( .IN1(n1338), .IN2(n2959), .Q(n4126) );
  AO21X1 U3918 ( .IN1(\fpu_add_ctl/n90 ), .IN2(n4179), .IN3(
        \fpu_add_frac_dp/n596 ), .Q(n4119) );
  NAND2X0 U3919 ( .IN1(n2959), .IN2(n2960), .QN(n4179) );
  INVX0 U3920 ( .INP(n4180), .ZN(n4178) );
  OA22X1 U3921 ( .IN1(n4181), .IN2(\fpu_add_ctl/n315 ), .IN3(n4182), .IN4(
        n4183), .Q(n2962) );
  AO221X1 U3922 ( .IN1(n1462), .IN2(n764), .IN3(n1339), .IN4(n4184), .IN5(
        n4185), .Q(\fpu_add_exp_dp/n539 ) );
  AO221X1 U3923 ( .IN1(n4186), .IN2(n1337), .IN3(n1463), .IN4(n738), .IN5(
        n4187), .Q(\fpu_add_exp_dp/n538 ) );
  AO21X1 U3924 ( .IN1(n4117), .IN2(n4128), .IN3(n4185), .Q(n4187) );
  INVX0 U3925 ( .INP(n4188), .ZN(n4117) );
  AO221X1 U3926 ( .IN1(n1337), .IN2(n4189), .IN3(n1463), .IN4(n737), .IN5(
        n4185), .Q(\fpu_add_exp_dp/n537 ) );
  OAI21X1 U3927 ( .IN1(n4136), .IN2(n4186), .IN3(n4190), .QN(n4189) );
  AO221X1 U3928 ( .IN1(n1340), .IN2(n4191), .IN3(n1463), .IN4(n736), .IN5(
        n4185), .Q(\fpu_add_exp_dp/n536 ) );
  AO21X1 U3929 ( .IN1(n4142), .IN2(n4190), .IN3(n4192), .Q(n4191) );
  AO221X1 U3930 ( .IN1(n1339), .IN2(n4193), .IN3(n1463), .IN4(n735), .IN5(
        n4185), .Q(\fpu_add_exp_dp/n535 ) );
  OAI21X1 U3931 ( .IN1(n4194), .IN2(n4192), .IN3(n4195), .QN(n4193) );
  AO221X1 U3932 ( .IN1(n1338), .IN2(n4196), .IN3(n1464), .IN4(n734), .IN5(
        n4185), .Q(\fpu_add_exp_dp/n534 ) );
  AO21X1 U3933 ( .IN1(n4154), .IN2(n4195), .IN3(n4197), .Q(n4196) );
  AO221X1 U3934 ( .IN1(n1337), .IN2(n4198), .IN3(n1463), .IN4(n733), .IN5(
        n4185), .Q(\fpu_add_exp_dp/n533 ) );
  OAI21X1 U3935 ( .IN1(n4199), .IN2(n4197), .IN3(n4200), .QN(n4198) );
  AO221X1 U3936 ( .IN1(n1340), .IN2(n4201), .IN3(n1464), .IN4(n732), .IN5(
        n4185), .Q(\fpu_add_exp_dp/n532 ) );
  AO21X1 U3937 ( .IN1(n4166), .IN2(n4200), .IN3(n4202), .Q(n4201) );
  AO221X1 U3938 ( .IN1(n1339), .IN2(n4203), .IN3(n1464), .IN4(n442), .IN5(
        n4185), .Q(\fpu_add_exp_dp/n531 ) );
  OAI21X1 U3939 ( .IN1(n4172), .IN2(n4202), .IN3(n4204), .QN(n4203) );
  AO221X1 U3940 ( .IN1(n1338), .IN2(n4205), .IN3(n1463), .IN4(n441), .IN5(
        n4185), .Q(\fpu_add_exp_dp/n530 ) );
  AO21X1 U3941 ( .IN1(n4174), .IN2(n4204), .IN3(n4206), .Q(n4205) );
  AO221X1 U3942 ( .IN1(n1337), .IN2(n4207), .IN3(n1464), .IN4(n443), .IN5(
        n4185), .Q(\fpu_add_exp_dp/n529 ) );
  AND2X1 U3943 ( .IN1(n1340), .IN2(n4208), .Q(n4185) );
  NAND3X0 U3944 ( .IN1(n2963), .IN2(n2956), .IN3(n2950), .QN(n4208) );
  AO22X1 U3945 ( .IN1(n4209), .IN2(n4182), .IN3(n4181), .IN4(n622), .Q(n2963)
         );
  AO22X1 U3946 ( .IN1(n4210), .IN2(n108), .IN3(n4211), .IN4(n552), .Q(n4181)
         );
  INVX0 U3947 ( .INP(n4183), .ZN(n4209) );
  XOR2X1 U3948 ( .IN1(n4177), .IN2(n4206), .Q(n4207) );
  NOR2X0 U3949 ( .IN1(n4204), .IN2(n4174), .QN(n4206) );
  INVX0 U3950 ( .INP(n4212), .ZN(n4174) );
  NAND2X0 U3951 ( .IN1(n4202), .IN2(n4172), .QN(n4204) );
  NOR2X0 U3952 ( .IN1(n4200), .IN2(n4166), .QN(n4202) );
  NAND2X0 U3953 ( .IN1(n4197), .IN2(n4199), .QN(n4200) );
  NOR2X0 U3954 ( .IN1(n4195), .IN2(n4154), .QN(n4197) );
  NAND2X0 U3955 ( .IN1(n4192), .IN2(n4194), .QN(n4195) );
  NOR2X0 U3956 ( .IN1(n4190), .IN2(n4142), .QN(n4192) );
  NAND2X0 U3957 ( .IN1(n4186), .IN2(n4136), .QN(n4190) );
  NOR2X0 U3958 ( .IN1(n4213), .IN2(n4128), .QN(n4186) );
  INVX0 U3959 ( .INP(n4214), .ZN(n4128) );
  INVX0 U3960 ( .INP(n4215), .ZN(n4177) );
  NAND3X0 U3961 ( .IN1(n4188), .IN2(n4216), .IN3(n4217), .QN(
        \fpu_add_exp_dp/n528 ) );
  OR2X1 U3962 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n22 ), .Q(n4217) );
  NAND2X0 U3963 ( .IN1(n4213), .IN2(n1337), .QN(n4188) );
  OAI221X1 U3964 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n21 ), .IN3(n4214), .IN4(
        n4057), .IN5(n4216), .QN(\fpu_add_exp_dp/n527 ) );
  OAI221X1 U3965 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n20 ), .IN3(n4136), .IN4(
        n4057), .IN5(n4216), .QN(\fpu_add_exp_dp/n526 ) );
  OAI221X1 U3966 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n19 ), .IN3(n4218), .IN4(
        n4057), .IN5(n4216), .QN(\fpu_add_exp_dp/n525 ) );
  OAI221X1 U3967 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n18 ), .IN3(n4194), .IN4(
        n4057), .IN5(n4216), .QN(\fpu_add_exp_dp/n524 ) );
  OAI221X1 U3968 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n17 ), .IN3(n4219), .IN4(
        n4057), .IN5(n4216), .QN(\fpu_add_exp_dp/n523 ) );
  OAI221X1 U3969 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n16 ), .IN3(n4199), .IN4(
        n4057), .IN5(n4216), .QN(\fpu_add_exp_dp/n522 ) );
  OAI221X1 U3970 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n15 ), .IN3(n4220), .IN4(
        n4057), .IN5(n4216), .QN(\fpu_add_exp_dp/n521 ) );
  OAI221X1 U3971 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n14 ), .IN3(n4057), .IN4(
        n4172), .IN5(n4216), .QN(\fpu_add_exp_dp/n520 ) );
  OAI221X1 U3972 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n13 ), .IN3(n4057), .IN4(
        n4212), .IN5(n4216), .QN(\fpu_add_exp_dp/n519 ) );
  OAI221X1 U3973 ( .IN1(n4114), .IN2(\fpu_add_exp_dp/n12 ), .IN3(n4057), .IN4(
        n4215), .IN5(n4216), .QN(\fpu_add_exp_dp/n518 ) );
  NAND3X0 U3974 ( .IN1(n1337), .IN2(n4183), .IN3(\fpu_add_ctl/n315 ), .QN(
        n4216) );
  NAND2X0 U3975 ( .IN1(n2959), .IN2(n4221), .QN(n4183) );
  AO21X1 U3976 ( .IN1(n296), .IN2(n927), .IN3(n55), .Q(n4221) );
  AO21X1 U3977 ( .IN1(n1466), .IN2(n1236), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n517 ) );
  AO21X1 U3978 ( .IN1(n1467), .IN2(n1237), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n516 ) );
  AO21X1 U3979 ( .IN1(n1466), .IN2(n1225), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n515 ) );
  AO21X1 U3980 ( .IN1(n1466), .IN2(n1226), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n514 ) );
  AO21X1 U3981 ( .IN1(n1467), .IN2(n1227), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n513 ) );
  AO21X1 U3982 ( .IN1(n1467), .IN2(n1228), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n512 ) );
  AO21X1 U3983 ( .IN1(n1467), .IN2(n1229), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n511 ) );
  AO21X1 U3984 ( .IN1(n1467), .IN2(n1230), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n510 ) );
  AO21X1 U3985 ( .IN1(n1467), .IN2(n1231), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n509 ) );
  AO21X1 U3986 ( .IN1(n1467), .IN2(n1232), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n508 ) );
  AO21X1 U3987 ( .IN1(n1467), .IN2(n1238), .IN3(n4222), .Q(
        \fpu_add_exp_dp/n507 ) );
  AND3X1 U3988 ( .IN1(n2950), .IN2(n2956), .IN3(n1339), .Q(n4222) );
  AND3X1 U3989 ( .IN1(n2952), .IN2(n2948), .IN3(n2944), .Q(n2950) );
  AND3X1 U3990 ( .IN1(n2946), .IN2(n2942), .IN3(n2937), .Q(n2944) );
  AND3X1 U3991 ( .IN1(n2985), .IN2(n2940), .IN3(n2930), .Q(n2937) );
  INVX0 U3992 ( .INP(n2934), .ZN(n2930) );
  NAND3X0 U3993 ( .IN1(n2932), .IN2(n2928), .IN3(n2924), .QN(n2934) );
  AND3X1 U3994 ( .IN1(n2926), .IN2(n2922), .IN3(n2918), .Q(n2924) );
  AND3X1 U3995 ( .IN1(n2920), .IN2(n2916), .IN3(n2912), .Q(n2918) );
  AND3X1 U3996 ( .IN1(n2914), .IN2(n2910), .IN3(n2906), .Q(n2912) );
  AND3X1 U3997 ( .IN1(n2908), .IN2(n2904), .IN3(n2900), .Q(n2906) );
  AND3X1 U3998 ( .IN1(n2902), .IN2(n2898), .IN3(n2894), .Q(n2900) );
  AND3X1 U3999 ( .IN1(n2896), .IN2(n2891), .IN3(n2892), .Q(n2894) );
  INVX0 U4000 ( .INP(n2889), .ZN(n2892) );
  NAND2X0 U4001 ( .IN1(n2887), .IN2(n2888), .QN(n2889) );
  AO22X1 U4002 ( .IN1(n2878), .IN2(n2984), .IN3(n4223), .IN4(n2884), .Q(n2887)
         );
  NAND2X0 U4003 ( .IN1(n2885), .IN2(n2883), .QN(n4223) );
  INVX0 U4004 ( .INP(n2984), .ZN(n2885) );
  INVX0 U4005 ( .INP(n2883), .ZN(n2878) );
  NAND3X0 U4006 ( .IN1(n2983), .IN2(n2881), .IN3(n2869), .QN(n2883) );
  INVX0 U4007 ( .INP(n2875), .ZN(n2869) );
  NAND3X0 U4008 ( .IN1(n2982), .IN2(n2867), .IN3(n2863), .QN(n2875) );
  INVX0 U4009 ( .INP(n2872), .ZN(n2863) );
  NAND3X0 U4010 ( .IN1(n2981), .IN2(n2980), .IN3(n2856), .QN(n2872) );
  INVX0 U4011 ( .INP(n2860), .ZN(n2856) );
  NAND3X0 U4012 ( .IN1(n2858), .IN2(n2854), .IN3(n2850), .QN(n2860) );
  AND3X1 U4013 ( .IN1(n2852), .IN2(n2848), .IN3(n2844), .Q(n2850) );
  AND3X1 U4014 ( .IN1(n2846), .IN2(n2842), .IN3(n2838), .Q(n2844) );
  AND3X1 U4015 ( .IN1(n2840), .IN2(n2836), .IN3(n2832), .Q(n2838) );
  AND3X1 U4016 ( .IN1(n2834), .IN2(n2830), .IN3(n2826), .Q(n2832) );
  AND3X1 U4017 ( .IN1(n2979), .IN2(n2978), .IN3(n2817), .Q(n2826) );
  INVX0 U4018 ( .INP(n2823), .ZN(n2817) );
  NAND3X0 U4019 ( .IN1(n2977), .IN2(n2815), .IN3(n2811), .QN(n2823) );
  INVX0 U4020 ( .INP(n2820), .ZN(n2811) );
  NAND3X0 U4021 ( .IN1(n2976), .IN2(n2975), .IN3(n2802), .QN(n2820) );
  INVX0 U4022 ( .INP(n2808), .ZN(n2802) );
  NAND3X0 U4023 ( .IN1(n2974), .IN2(n2800), .IN3(n2796), .QN(n2808) );
  INVX0 U4024 ( .INP(n2805), .ZN(n2796) );
  NAND3X0 U4025 ( .IN1(n2798), .IN2(n2794), .IN3(n2790), .QN(n2805) );
  AND3X1 U4026 ( .IN1(n2792), .IN2(n2788), .IN3(n2784), .Q(n2790) );
  OA21X1 U4027 ( .IN1(n108), .IN2(n21), .IN3(n2786), .Q(n2784) );
  NOR2X0 U4028 ( .IN1(\fpu_add_exp_dp/n256 ), .IN2(\fpu_add_frac_dp/n2189 ), 
        .QN(\fpu_add_exp_dp/n448 ) );
  INVX0 U4029 ( .INP(rclk), .ZN(\fpu_add_frac_dp/n2189 ) );
  NOR2X0 U4030 ( .IN1(\fpu_add_exp_dp/n435 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N9 ) );
  NOR2X0 U4031 ( .IN1(\fpu_add_exp_dp/n433 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N8 ) );
  NOR2X0 U4032 ( .IN1(\fpu_add_exp_dp/n432 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N7 ) );
  NOR2X0 U4033 ( .IN1(\fpu_add_exp_dp/n434 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N6 ) );
  NOR2X0 U4034 ( .IN1(\fpu_add_exp_dp/n431 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N5 ) );
  NOR2X0 U4035 ( .IN1(\fpu_add_exp_dp/n436 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N4 ) );
  NOR2X0 U4036 ( .IN1(\fpu_add_exp_dp/n444 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N3 ) );
  NOR2X0 U4037 ( .IN1(\fpu_add_exp_dp/n447 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N14 ) );
  NOR2X0 U4038 ( .IN1(\fpu_add_exp_dp/n446 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N13 ) );
  NOR2X0 U4039 ( .IN1(\fpu_add_exp_dp/n443 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N12 ) );
  NOR2X0 U4040 ( .IN1(\fpu_add_exp_dp/n445 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N11 ) );
  NOR2X0 U4041 ( .IN1(\fpu_add_exp_dp/n442 ), .IN2(n4224), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre4/N10 ) );
  NAND3X0 U4042 ( .IN1(n3143), .IN2(n4225), .IN3(n4226), .QN(n4224) );
  NAND2X0 U4043 ( .IN1(n3171), .IN2(n3144), .QN(n4225) );
  INVX0 U4044 ( .INP(n3545), .ZN(n3143) );
  NOR2X0 U4045 ( .IN1(n4227), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N9 ) );
  AOI21X1 U4046 ( .IN1(n160), .IN2(n4229), .IN3(n4230), .QN(n4227) );
  NOR2X0 U4047 ( .IN1(n4231), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N8 ) );
  OA21X1 U4048 ( .IN1(\fpu_add_exp_dp/n433 ), .IN2(n4232), .IN3(n4229), .Q(
        n4231) );
  NOR2X0 U4049 ( .IN1(n4233), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N7 ) );
  AOI21X1 U4050 ( .IN1(n67), .IN2(n4234), .IN3(n4232), .QN(n4233) );
  NOR2X0 U4051 ( .IN1(n4235), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N6 ) );
  OA21X1 U4052 ( .IN1(\fpu_add_exp_dp/n434 ), .IN2(n4236), .IN3(n4234), .Q(
        n4235) );
  NOR2X0 U4053 ( .IN1(n4237), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N5 ) );
  AOI21X1 U4054 ( .IN1(n159), .IN2(n4238), .IN3(n4236), .QN(n4237) );
  NOR2X0 U4055 ( .IN1(n4239), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N4 ) );
  OA21X1 U4056 ( .IN1(\fpu_add_exp_dp/n444 ), .IN2(\fpu_add_exp_dp/n436 ), 
        .IN3(n4238), .Q(n4239) );
  NOR2X0 U4057 ( .IN1(n583), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N3 ) );
  NOR2X0 U4058 ( .IN1(\fpu_add_exp_dp/n447 ), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N14 ) );
  NOR3X0 U4059 ( .IN1(n4228), .IN2(\fpu_add_exp_dp/n446 ), .IN3(n4240), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N13 ) );
  NOR2X0 U4060 ( .IN1(n4241), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N12 ) );
  AOI21X1 U4061 ( .IN1(n17), .IN2(n4242), .IN3(n4240), .QN(n4241) );
  NOR2X0 U4062 ( .IN1(n4242), .IN2(n17), .QN(n4240) );
  INVX0 U4063 ( .INP(n4243), .ZN(n4242) );
  NOR2X0 U4064 ( .IN1(n4244), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N11 ) );
  AOI21X1 U4065 ( .IN1(n71), .IN2(n4245), .IN3(n4243), .QN(n4244) );
  NOR2X0 U4066 ( .IN1(n4245), .IN2(n71), .QN(n4243) );
  NOR2X0 U4067 ( .IN1(n4246), .IN2(n4228), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre3/N10 ) );
  NAND4X0 U4068 ( .IN1(n3175), .IN2(n4226), .IN3(n2601), .IN4(n3144), .QN(
        n4228) );
  INVX0 U4069 ( .INP(n3547), .ZN(n3144) );
  NOR2X0 U4070 ( .IN1(n583), .IN2(n3146), .QN(n3547) );
  NAND4X0 U4071 ( .IN1(\fpu_add_exp_dp/n435 ), .IN2(\fpu_add_exp_dp/n434 ), 
        .IN3(n4247), .IN4(n4248), .QN(n3146) );
  NOR4X0 U4072 ( .IN1(n17), .IN2(n4249), .IN3(n71), .IN4(n181), .QN(n4248) );
  NAND2X0 U4073 ( .IN1(\fpu_add_exp_dp/n442 ), .IN2(\fpu_add_exp_dp/n436 ), 
        .QN(n4249) );
  AND3X1 U4074 ( .IN1(\fpu_add_exp_dp/n433 ), .IN2(\fpu_add_exp_dp/n432 ), 
        .IN3(\fpu_add_exp_dp/n431 ), .Q(n4247) );
  NOR2X0 U4075 ( .IN1(n3545), .IN2(n3141), .QN(n2601) );
  INVX0 U4076 ( .INP(n3171), .ZN(n3141) );
  XNOR3X1 U4077 ( .IN1(\fpu_add_frac_dp/n673 ), .IN2(\fpu_add_frac_dp/n568 ), 
        .IN3(n4250), .Q(n3171) );
  INVX0 U4078 ( .INP(n2602), .ZN(n3175) );
  XNOR3X1 U4079 ( .IN1(\fpu_add_frac_dp/n674 ), .IN2(\fpu_add_frac_dp/n567 ), 
        .IN3(n4251), .Q(n2602) );
  OA21X1 U4080 ( .IN1(\fpu_add_exp_dp/n442 ), .IN2(n4230), .IN3(n4245), .Q(
        n4246) );
  NAND2X0 U4081 ( .IN1(n4230), .IN2(\fpu_add_exp_dp/n442 ), .QN(n4245) );
  NOR2X0 U4082 ( .IN1(n4229), .IN2(n160), .QN(n4230) );
  NAND2X0 U4083 ( .IN1(n4232), .IN2(\fpu_add_exp_dp/n433 ), .QN(n4229) );
  NOR2X0 U4084 ( .IN1(n4234), .IN2(n67), .QN(n4232) );
  NAND2X0 U4085 ( .IN1(n4236), .IN2(\fpu_add_exp_dp/n434 ), .QN(n4234) );
  NOR2X0 U4086 ( .IN1(n4238), .IN2(n159), .QN(n4236) );
  AO222X1 U4087 ( .IN1(n4252), .IN2(n160), .IN3(n4253), .IN4(n4161), .IN5(
        n1461), .IN6(n4199), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N9 ) );
  AO21X1 U4088 ( .IN1(n4254), .IN2(n666), .IN3(n4255), .Q(n4161) );
  AO222X1 U4089 ( .IN1(n4252), .IN2(n69), .IN3(n4253), .IN4(n4155), .IN5(n1461), .IN6(n4219), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N8 ) );
  INVX0 U4090 ( .INP(n4150), .ZN(n4155) );
  XNOR3X1 U4091 ( .IN1(\fpu_add_frac_dp/n593 ), .IN2(\fpu_add_exp_dp/n441 ), 
        .IN3(n4256), .Q(n4150) );
  AO222X1 U4092 ( .IN1(n4252), .IN2(n67), .IN3(n4253), .IN4(n4149), .IN5(n1462), .IN6(n4194), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N7 ) );
  XOR3X1 U4093 ( .IN1(\fpu_add_frac_dp/n594 ), .IN2(\fpu_add_exp_dp/n440 ), 
        .IN3(n4257), .Q(n4149) );
  AO222X1 U4094 ( .IN1(n4252), .IN2(n178), .IN3(n4253), .IN4(n4143), .IN5(
        n1462), .IN6(n4218), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N6 ) );
  XOR3X1 U4095 ( .IN1(\fpu_add_frac_dp/n2307 ), .IN2(\fpu_add_exp_dp/n439 ), 
        .IN3(n4258), .Q(n4143) );
  AO222X1 U4096 ( .IN1(n4252), .IN2(n159), .IN3(n4253), .IN4(n4137), .IN5(
        n1461), .IN6(n4136), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N5 ) );
  XOR3X1 U4097 ( .IN1(\fpu_add_frac_dp/n2471 ), .IN2(\fpu_add_exp_dp/n438 ), 
        .IN3(n4259), .Q(n4137) );
  AO222X1 U4098 ( .IN1(n4252), .IN2(n72), .IN3(n4253), .IN4(n4130), .IN5(n1462), .IN6(n4214), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N4 ) );
  INVX0 U4099 ( .INP(n4121), .ZN(n4130) );
  XOR3X1 U4100 ( .IN1(n4260), .IN2(\fpu_add_frac_dp/n2460 ), .IN3(n643), .Q(
        n4121) );
  AO222X1 U4101 ( .IN1(n4252), .IN2(n583), .IN3(n4253), .IN4(n4261), .IN5(
        n1461), .IN6(n4184), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N3 ) );
  INVX0 U4102 ( .INP(n4118), .ZN(n4261) );
  OA21X1 U4103 ( .IN1(n154), .IN2(\fpu_add_exp_dp/n57 ), .IN3(n4262), .Q(n4118) );
  AO222X1 U4104 ( .IN1(n4252), .IN2(n728), .IN3(n4263), .IN4(n4253), .IN5(
        n1461), .IN6(n4264), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N14 ) );
  XNOR2X1 U4105 ( .IN1(\fpu_add_exp_dp/n46 ), .IN2(n4265), .Q(n4263) );
  AO222X1 U4106 ( .IN1(n4252), .IN2(n181), .IN3(n4253), .IN4(n4180), .IN5(
        n1461), .IN6(n4215), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N13 ) );
  AO21X1 U4107 ( .IN1(n663), .IN2(n4266), .IN3(n4265), .Q(n4180) );
  NOR2X0 U4108 ( .IN1(n663), .IN2(n4266), .QN(n4265) );
  AO222X1 U4109 ( .IN1(n4252), .IN2(n17), .IN3(n4253), .IN4(n4267), .IN5(n1461), .IN6(n4212), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N12 ) );
  INVX0 U4110 ( .INP(n4175), .ZN(n4267) );
  OA21X1 U4111 ( .IN1(\fpu_add_exp_dp/n48 ), .IN2(n4268), .IN3(n4266), .Q(
        n4175) );
  NAND2X0 U4112 ( .IN1(\fpu_add_exp_dp/n48 ), .IN2(n4268), .QN(n4266) );
  INVX0 U4113 ( .INP(n4269), .ZN(n4268) );
  AO222X1 U4114 ( .IN1(n4252), .IN2(n71), .IN3(n4253), .IN4(n4270), .IN5(n1461), .IN6(n4172), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N11 ) );
  INVX0 U4115 ( .INP(n4170), .ZN(n4270) );
  OA21X1 U4116 ( .IN1(\fpu_add_exp_dp/n450 ), .IN2(n4271), .IN3(n4269), .Q(
        n4170) );
  NAND2X0 U4117 ( .IN1(\fpu_add_exp_dp/n450 ), .IN2(n4271), .QN(n4269) );
  INVX0 U4118 ( .INP(n4272), .ZN(n4271) );
  AO222X1 U4119 ( .IN1(n4253), .IN2(n4167), .IN3(n4252), .IN4(n256), .IN5(
        n1461), .IN6(n4220), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre2/N10 ) );
  AND2X1 U4120 ( .IN1(n1337), .IN2(\fpu_add_ctl/a3stg_opdec_9_0[3] ), .Q(n4252) );
  INVX0 U4121 ( .INP(n4162), .ZN(n4167) );
  OA21X1 U4122 ( .IN1(n4255), .IN2(\fpu_add_exp_dp/n50 ), .IN3(n4272), .Q(
        n4162) );
  NAND2X0 U4123 ( .IN1(\fpu_add_exp_dp/n50 ), .IN2(n4255), .QN(n4272) );
  NOR2X0 U4124 ( .IN1(n666), .IN2(n4254), .QN(n4255) );
  AO22X1 U4125 ( .IN1(n4273), .IN2(n761), .IN3(\fpu_add_frac_dp/n593 ), .IN4(
        n4274), .Q(n4254) );
  NAND2X0 U4126 ( .IN1(\fpu_add_exp_dp/n441 ), .IN2(n4256), .QN(n4274) );
  INVX0 U4127 ( .INP(n4256), .ZN(n4273) );
  AO22X1 U4128 ( .IN1(\fpu_add_exp_dp/n440 ), .IN2(n4257), .IN3(n4275), .IN4(
        n762), .Q(n4256) );
  OR2X1 U4129 ( .IN1(n4257), .IN2(\fpu_add_exp_dp/n440 ), .Q(n4275) );
  AO22X1 U4130 ( .IN1(\fpu_add_exp_dp/n439 ), .IN2(n4258), .IN3(n4276), .IN4(
        n584), .Q(n4257) );
  OR2X1 U4131 ( .IN1(n4258), .IN2(\fpu_add_exp_dp/n439 ), .Q(n4276) );
  AO22X1 U4132 ( .IN1(\fpu_add_exp_dp/n438 ), .IN2(n4259), .IN3(n4277), .IN4(
        n63), .Q(n4258) );
  OR2X1 U4133 ( .IN1(n4259), .IN2(\fpu_add_exp_dp/n438 ), .Q(n4277) );
  AO22X1 U4134 ( .IN1(n4260), .IN2(\fpu_add_exp_dp/n437 ), .IN3(n4278), .IN4(
        n582), .Q(n4259) );
  NAND2X0 U4135 ( .IN1(n643), .IN2(n4262), .QN(n4278) );
  INVX0 U4136 ( .INP(n4262), .ZN(n4260) );
  NAND2X0 U4137 ( .IN1(\fpu_add_exp_dp/n57 ), .IN2(n154), .QN(n4262) );
  NOR3X0 U4138 ( .IN1(n642), .IN2(\fpu_add_frac_dp/n596 ), .IN3(n4057), .QN(
        n4253) );
  NOR3X0 U4139 ( .IN1(n4279), .IN2(n4280), .IN3(n4281), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N9 ) );
  OA21X1 U4140 ( .IN1(\fpu_add_exp_dp/n433 ), .IN2(n4282), .IN3(
        \fpu_add_exp_dp/n435 ), .Q(n4281) );
  NOR2X0 U4141 ( .IN1(n4279), .IN2(n4283), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N8 ) );
  XOR2X1 U4142 ( .IN1(n69), .IN2(n4282), .Q(n4283) );
  NOR3X0 U4143 ( .IN1(n4279), .IN2(n4284), .IN3(n4285), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N7 ) );
  OA21X1 U4144 ( .IN1(\fpu_add_exp_dp/n434 ), .IN2(n4286), .IN3(
        \fpu_add_exp_dp/n432 ), .Q(n4285) );
  NOR2X0 U4145 ( .IN1(n4279), .IN2(n4287), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N6 ) );
  XOR2X1 U4146 ( .IN1(\fpu_add_exp_dp/n434 ), .IN2(n4288), .Q(n4287) );
  NOR3X0 U4147 ( .IN1(n4279), .IN2(n4288), .IN3(n4289), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N5 ) );
  OA21X1 U4148 ( .IN1(\fpu_add_exp_dp/n444 ), .IN2(\fpu_add_exp_dp/n436 ), 
        .IN3(\fpu_add_exp_dp/n431 ), .Q(n4289) );
  OA21X1 U4149 ( .IN1(n4290), .IN2(\fpu_add_exp_dp/i_a4stg_exp_pre1/N3 ), 
        .IN3(n4238), .Q(\fpu_add_exp_dp/i_a4stg_exp_pre1/N4 ) );
  NAND2X0 U4150 ( .IN1(\fpu_add_exp_dp/n444 ), .IN2(\fpu_add_exp_dp/n436 ), 
        .QN(n4238) );
  NOR2X0 U4151 ( .IN1(n72), .IN2(n4279), .QN(n4290) );
  NOR2X0 U4152 ( .IN1(n4279), .IN2(n583), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N3 ) );
  NOR2X0 U4153 ( .IN1(n4279), .IN2(n4291), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N14 ) );
  XOR2X1 U4154 ( .IN1(\fpu_add_exp_dp/n447 ), .IN2(n4292), .Q(n4291) );
  NOR3X0 U4155 ( .IN1(n4279), .IN2(n4292), .IN3(n4293), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N13 ) );
  OA21X1 U4156 ( .IN1(\fpu_add_exp_dp/n443 ), .IN2(n4294), .IN3(
        \fpu_add_exp_dp/n446 ), .Q(n4293) );
  NOR3X0 U4157 ( .IN1(\fpu_add_exp_dp/n443 ), .IN2(\fpu_add_exp_dp/n446 ), 
        .IN3(n4294), .QN(n4292) );
  NOR2X0 U4158 ( .IN1(n4279), .IN2(n4295), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N12 ) );
  XOR2X1 U4159 ( .IN1(n17), .IN2(n4294), .Q(n4295) );
  NOR3X0 U4160 ( .IN1(n4279), .IN2(n4296), .IN3(n4297), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N11 ) );
  OA21X1 U4161 ( .IN1(\fpu_add_exp_dp/n442 ), .IN2(n4298), .IN3(
        \fpu_add_exp_dp/n445 ), .Q(n4297) );
  INVX0 U4162 ( .INP(n4294), .ZN(n4296) );
  NAND3X0 U4163 ( .IN1(n256), .IN2(n71), .IN3(n4280), .QN(n4294) );
  NOR2X0 U4164 ( .IN1(n4279), .IN2(n4299), .QN(
        \fpu_add_exp_dp/i_a4stg_exp_pre1/N10 ) );
  XOR2X1 U4165 ( .IN1(\fpu_add_exp_dp/n442 ), .IN2(n4280), .Q(n4299) );
  INVX0 U4166 ( .INP(n4298), .ZN(n4280) );
  NAND3X0 U4167 ( .IN1(n69), .IN2(n160), .IN3(n4284), .QN(n4298) );
  INVX0 U4168 ( .INP(n4282), .ZN(n4284) );
  NAND3X0 U4169 ( .IN1(n67), .IN2(n178), .IN3(n4288), .QN(n4282) );
  INVX0 U4170 ( .INP(n4286), .ZN(n4288) );
  NAND3X0 U4171 ( .IN1(n72), .IN2(n583), .IN3(n159), .QN(n4286) );
  NAND2X0 U4172 ( .IN1(n4226), .IN2(n3545), .QN(n4279) );
  XNOR2X1 U4173 ( .IN1(\fpu_add_frac_dp/n569 ), .IN2(n4300), .Q(n3545) );
  OA22X1 U4174 ( .IN1(n4301), .IN2(n453), .IN3(n753), .IN4(n4250), .Q(n4300)
         );
  AND2X1 U4175 ( .IN1(n4250), .IN2(n753), .Q(n4301) );
  AO22X1 U4176 ( .IN1(n4251), .IN2(n359), .IN3(n4302), .IN4(n768), .Q(n4250)
         );
  OR2X1 U4177 ( .IN1(n359), .IN2(n4251), .Q(n4302) );
  AO22X1 U4178 ( .IN1(n3207), .IN2(n360), .IN3(n4303), .IN4(n769), .Q(n4251)
         );
  OR2X1 U4179 ( .IN1(n360), .IN2(n3207), .Q(n4303) );
  AO22X1 U4180 ( .IN1(n3209), .IN2(n361), .IN3(n4304), .IN4(n770), .Q(n3207)
         );
  OR2X1 U4181 ( .IN1(n361), .IN2(n3209), .Q(n4304) );
  AO22X1 U4182 ( .IN1(n3221), .IN2(n362), .IN3(n4305), .IN4(n771), .Q(n3209)
         );
  OR2X1 U4183 ( .IN1(n362), .IN2(n3221), .Q(n4305) );
  AO22X1 U4184 ( .IN1(n3241), .IN2(n363), .IN3(n4306), .IN4(n772), .Q(n3221)
         );
  OR2X1 U4185 ( .IN1(n363), .IN2(n3241), .Q(n4306) );
  AO22X1 U4186 ( .IN1(n3244), .IN2(n364), .IN3(n4307), .IN4(n773), .Q(n3241)
         );
  OR2X1 U4187 ( .IN1(n364), .IN2(n3244), .Q(n4307) );
  AO22X1 U4188 ( .IN1(n3265), .IN2(n365), .IN3(n4308), .IN4(n774), .Q(n3244)
         );
  OR2X1 U4189 ( .IN1(n365), .IN2(n3265), .Q(n4308) );
  AO22X1 U4190 ( .IN1(n3273), .IN2(n366), .IN3(n4309), .IN4(n775), .Q(n3265)
         );
  OR2X1 U4191 ( .IN1(n366), .IN2(n3273), .Q(n4309) );
  AO22X1 U4192 ( .IN1(n3281), .IN2(n367), .IN3(n4310), .IN4(n776), .Q(n3273)
         );
  OR2X1 U4193 ( .IN1(n367), .IN2(n3281), .Q(n4310) );
  AO22X1 U4194 ( .IN1(n3286), .IN2(n368), .IN3(n4311), .IN4(n777), .Q(n3281)
         );
  OR2X1 U4195 ( .IN1(n368), .IN2(n3286), .Q(n4311) );
  AO22X1 U4196 ( .IN1(n3291), .IN2(n369), .IN3(n4312), .IN4(n778), .Q(n3286)
         );
  OR2X1 U4197 ( .IN1(n369), .IN2(n3291), .Q(n4312) );
  AO22X1 U4198 ( .IN1(n3296), .IN2(n370), .IN3(n4313), .IN4(n779), .Q(n3291)
         );
  OR2X1 U4199 ( .IN1(n370), .IN2(n3296), .Q(n4313) );
  AO22X1 U4200 ( .IN1(n3309), .IN2(n371), .IN3(n4314), .IN4(n780), .Q(n3296)
         );
  OR2X1 U4201 ( .IN1(n371), .IN2(n3309), .Q(n4314) );
  AO22X1 U4202 ( .IN1(n3315), .IN2(n372), .IN3(n4315), .IN4(n781), .Q(n3309)
         );
  OR2X1 U4203 ( .IN1(n372), .IN2(n3315), .Q(n4315) );
  AO22X1 U4204 ( .IN1(n3323), .IN2(n373), .IN3(n4316), .IN4(n782), .Q(n3315)
         );
  OR2X1 U4205 ( .IN1(n373), .IN2(n3323), .Q(n4316) );
  AO22X1 U4206 ( .IN1(n3329), .IN2(n374), .IN3(n4317), .IN4(n783), .Q(n3323)
         );
  OR2X1 U4207 ( .IN1(n374), .IN2(n3329), .Q(n4317) );
  AO22X1 U4208 ( .IN1(n3335), .IN2(n375), .IN3(n4318), .IN4(n784), .Q(n3329)
         );
  OR2X1 U4209 ( .IN1(n375), .IN2(n3335), .Q(n4318) );
  AO22X1 U4210 ( .IN1(n3341), .IN2(n376), .IN3(n4319), .IN4(n785), .Q(n3335)
         );
  OR2X1 U4211 ( .IN1(n376), .IN2(n3341), .Q(n4319) );
  AO22X1 U4212 ( .IN1(n3347), .IN2(n377), .IN3(n4320), .IN4(n786), .Q(n3341)
         );
  OR2X1 U4213 ( .IN1(n377), .IN2(n3347), .Q(n4320) );
  AO22X1 U4214 ( .IN1(n3353), .IN2(n378), .IN3(n4321), .IN4(n787), .Q(n3347)
         );
  OR2X1 U4215 ( .IN1(n378), .IN2(n3353), .Q(n4321) );
  AO22X1 U4216 ( .IN1(n3359), .IN2(n379), .IN3(n4322), .IN4(n788), .Q(n3353)
         );
  OR2X1 U4217 ( .IN1(n379), .IN2(n3359), .Q(n4322) );
  AO22X1 U4218 ( .IN1(n3365), .IN2(n380), .IN3(n4323), .IN4(n789), .Q(n3359)
         );
  OR2X1 U4219 ( .IN1(n380), .IN2(n3365), .Q(n4323) );
  AO22X1 U4220 ( .IN1(n3371), .IN2(n381), .IN3(n4324), .IN4(n790), .Q(n3365)
         );
  OR2X1 U4221 ( .IN1(n381), .IN2(n3371), .Q(n4324) );
  AO22X1 U4222 ( .IN1(n3377), .IN2(n382), .IN3(n4325), .IN4(n791), .Q(n3371)
         );
  OR2X1 U4223 ( .IN1(n382), .IN2(n3377), .Q(n4325) );
  AO22X1 U4224 ( .IN1(n3383), .IN2(n383), .IN3(n4326), .IN4(n792), .Q(n3377)
         );
  OR2X1 U4225 ( .IN1(n383), .IN2(n3383), .Q(n4326) );
  AO22X1 U4226 ( .IN1(n3389), .IN2(n384), .IN3(n4327), .IN4(n793), .Q(n3383)
         );
  OR2X1 U4227 ( .IN1(n384), .IN2(n3389), .Q(n4327) );
  AO22X1 U4228 ( .IN1(n3395), .IN2(n385), .IN3(n4328), .IN4(n794), .Q(n3389)
         );
  OR2X1 U4229 ( .IN1(n385), .IN2(n3395), .Q(n4328) );
  AO22X1 U4230 ( .IN1(n3401), .IN2(n386), .IN3(n4329), .IN4(n795), .Q(n3395)
         );
  OR2X1 U4231 ( .IN1(n386), .IN2(n3401), .Q(n4329) );
  AO22X1 U4232 ( .IN1(n3407), .IN2(n387), .IN3(n4330), .IN4(n796), .Q(n3401)
         );
  OR2X1 U4233 ( .IN1(n387), .IN2(n3407), .Q(n4330) );
  AO22X1 U4234 ( .IN1(n3413), .IN2(n388), .IN3(n4331), .IN4(n797), .Q(n3407)
         );
  OR2X1 U4235 ( .IN1(n388), .IN2(n3413), .Q(n4331) );
  AO22X1 U4236 ( .IN1(n3419), .IN2(n389), .IN3(n4332), .IN4(n798), .Q(n3413)
         );
  OR2X1 U4237 ( .IN1(n389), .IN2(n3419), .Q(n4332) );
  AO22X1 U4238 ( .IN1(n3425), .IN2(n390), .IN3(n4333), .IN4(n799), .Q(n3419)
         );
  OR2X1 U4239 ( .IN1(n390), .IN2(n3425), .Q(n4333) );
  AO22X1 U4240 ( .IN1(n3431), .IN2(n391), .IN3(n4334), .IN4(n800), .Q(n3425)
         );
  OR2X1 U4241 ( .IN1(n391), .IN2(n3431), .Q(n4334) );
  AO22X1 U4242 ( .IN1(n3437), .IN2(n392), .IN3(n4335), .IN4(n801), .Q(n3431)
         );
  OR2X1 U4243 ( .IN1(n392), .IN2(n3437), .Q(n4335) );
  AO22X1 U4244 ( .IN1(n3443), .IN2(n393), .IN3(n4336), .IN4(n802), .Q(n3437)
         );
  OR2X1 U4245 ( .IN1(n393), .IN2(n3443), .Q(n4336) );
  AO22X1 U4246 ( .IN1(n3450), .IN2(n394), .IN3(n4337), .IN4(n803), .Q(n3443)
         );
  OR2X1 U4247 ( .IN1(n394), .IN2(n3450), .Q(n4337) );
  AO22X1 U4248 ( .IN1(n3456), .IN2(n395), .IN3(n4338), .IN4(n804), .Q(n3450)
         );
  OR2X1 U4249 ( .IN1(n395), .IN2(n3456), .Q(n4338) );
  AO22X1 U4250 ( .IN1(n3462), .IN2(n396), .IN3(n4339), .IN4(n805), .Q(n3456)
         );
  OR2X1 U4251 ( .IN1(n396), .IN2(n3462), .Q(n4339) );
  AO22X1 U4252 ( .IN1(n3468), .IN2(n397), .IN3(n4340), .IN4(n806), .Q(n3462)
         );
  OR2X1 U4253 ( .IN1(n397), .IN2(n3468), .Q(n4340) );
  AO22X1 U4254 ( .IN1(n3474), .IN2(n398), .IN3(n4341), .IN4(n807), .Q(n3468)
         );
  OR2X1 U4255 ( .IN1(n398), .IN2(n3474), .Q(n4341) );
  AO22X1 U4256 ( .IN1(n3480), .IN2(n399), .IN3(n4342), .IN4(n808), .Q(n3474)
         );
  OR2X1 U4257 ( .IN1(n399), .IN2(n3480), .Q(n4342) );
  AO22X1 U4258 ( .IN1(n3486), .IN2(n400), .IN3(n4343), .IN4(n809), .Q(n3480)
         );
  OR2X1 U4259 ( .IN1(n400), .IN2(n3486), .Q(n4343) );
  AO22X1 U4260 ( .IN1(n3492), .IN2(n401), .IN3(n4344), .IN4(n810), .Q(n3486)
         );
  OR2X1 U4261 ( .IN1(n401), .IN2(n3492), .Q(n4344) );
  AO22X1 U4262 ( .IN1(n3495), .IN2(n402), .IN3(n4345), .IN4(n811), .Q(n3492)
         );
  OR2X1 U4263 ( .IN1(n402), .IN2(n3495), .Q(n4345) );
  AO22X1 U4264 ( .IN1(n3497), .IN2(n403), .IN3(n4346), .IN4(n812), .Q(n3495)
         );
  OR2X1 U4265 ( .IN1(n403), .IN2(n3497), .Q(n4346) );
  AO22X1 U4266 ( .IN1(n3505), .IN2(n404), .IN3(n4347), .IN4(n813), .Q(n3497)
         );
  OR2X1 U4267 ( .IN1(n404), .IN2(n3505), .Q(n4347) );
  AO22X1 U4268 ( .IN1(n3515), .IN2(n405), .IN3(n4348), .IN4(n814), .Q(n3505)
         );
  OR2X1 U4269 ( .IN1(n405), .IN2(n3515), .Q(n4348) );
  AO22X1 U4270 ( .IN1(n3521), .IN2(n406), .IN3(n4349), .IN4(n815), .Q(n3515)
         );
  OR2X1 U4271 ( .IN1(n406), .IN2(n3521), .Q(n4349) );
  AO22X1 U4272 ( .IN1(n3525), .IN2(n407), .IN3(n4350), .IN4(n816), .Q(n3521)
         );
  OR2X1 U4273 ( .IN1(n407), .IN2(n3525), .Q(n4350) );
  AO22X1 U4274 ( .IN1(n3530), .IN2(n408), .IN3(n4351), .IN4(n817), .Q(n3525)
         );
  OR2X1 U4275 ( .IN1(n408), .IN2(n3530), .Q(n4351) );
  AO22X1 U4276 ( .IN1(n3537), .IN2(n409), .IN3(n4352), .IN4(n818), .Q(n3530)
         );
  OR2X1 U4277 ( .IN1(n409), .IN2(n3537), .Q(n4352) );
  AO22X1 U4278 ( .IN1(n3548), .IN2(n410), .IN3(n4353), .IN4(n819), .Q(n3537)
         );
  OR2X1 U4279 ( .IN1(n410), .IN2(n3548), .Q(n4353) );
  AO22X1 U4280 ( .IN1(n3544), .IN2(n411), .IN3(n4354), .IN4(n820), .Q(n3548)
         );
  OR2X1 U4281 ( .IN1(n411), .IN2(n3544), .Q(n4354) );
  AO22X1 U4282 ( .IN1(n3137), .IN2(n412), .IN3(n4355), .IN4(n821), .Q(n3544)
         );
  OR2X1 U4283 ( .IN1(n412), .IN2(n3137), .Q(n4355) );
  AO22X1 U4284 ( .IN1(n3138), .IN2(n413), .IN3(n4356), .IN4(n822), .Q(n3137)
         );
  OR2X1 U4285 ( .IN1(n413), .IN2(n3138), .Q(n4356) );
  AO22X1 U4286 ( .IN1(n3148), .IN2(n414), .IN3(n4357), .IN4(n823), .Q(n3138)
         );
  OR2X1 U4287 ( .IN1(n414), .IN2(n3148), .Q(n4357) );
  AO22X1 U4288 ( .IN1(n3151), .IN2(n415), .IN3(n4358), .IN4(n824), .Q(n3148)
         );
  OR2X1 U4289 ( .IN1(n415), .IN2(n3151), .Q(n4358) );
  AO22X1 U4290 ( .IN1(n3150), .IN2(n416), .IN3(n4359), .IN4(n825), .Q(n3151)
         );
  OR2X1 U4291 ( .IN1(n416), .IN2(n3150), .Q(n4359) );
  AO22X1 U4292 ( .IN1(n3080), .IN2(n417), .IN3(n4360), .IN4(n826), .Q(n3150)
         );
  OR2X1 U4293 ( .IN1(n417), .IN2(n3080), .Q(n4360) );
  AO22X1 U4294 ( .IN1(n3087), .IN2(n418), .IN3(n4361), .IN4(n827), .Q(n3080)
         );
  OR2X1 U4295 ( .IN1(n418), .IN2(n3087), .Q(n4361) );
  AO22X1 U4296 ( .IN1(n3098), .IN2(n419), .IN3(n4362), .IN4(n828), .Q(n3087)
         );
  OR2X1 U4297 ( .IN1(n419), .IN2(n3098), .Q(n4362) );
  AO22X1 U4298 ( .IN1(n139), .IN2(n852), .IN3(n4363), .IN4(n465), .Q(n3098) );
  NAND2X0 U4299 ( .IN1(\fpu_add_frac_dp/n598 ), .IN2(\fpu_add_frac_dp/n509 ), 
        .QN(n4363) );
  NOR2X0 U4300 ( .IN1(n4057), .IN2(\fpu_add_ctl/n142 ), .QN(n4226) );
  NAND2X0 U4301 ( .IN1(fadd_clken_l), .IN2(\fpu_add_ctl/n470 ), .QN(
        \fpu_add_exp_dp/ckbuf_add_exp_dp/N1 ) );
  AO22X1 U4302 ( .IN1(n4364), .IN2(inq_op[7]), .IN3(n4365), .IN4(
        \fpu_add_ctl/n314 ), .Q(\fpu_add_ctl/n752 ) );
  AO22X1 U4303 ( .IN1(inq_op[6]), .IN2(n4364), .IN3(n4365), .IN4(
        \fpu_add_ctl/n312 ), .Q(\fpu_add_ctl/n751 ) );
  AO22X1 U4304 ( .IN1(inq_op[5]), .IN2(n4364), .IN3(n4365), .IN4(n84), .Q(
        \fpu_add_ctl/n750 ) );
  AO22X1 U4305 ( .IN1(inq_op[4]), .IN2(n4364), .IN3(n4365), .IN4(n585), .Q(
        \fpu_add_ctl/n749 ) );
  AO22X1 U4306 ( .IN1(inq_op[3]), .IN2(n4364), .IN3(n4365), .IN4(n595), .Q(
        \fpu_add_ctl/n748 ) );
  AO22X1 U4307 ( .IN1(inq_op[2]), .IN2(n4364), .IN3(n4365), .IN4(n18), .Q(
        \fpu_add_ctl/n747 ) );
  AO22X1 U4308 ( .IN1(n4364), .IN2(inq_op[1]), .IN3(n4365), .IN4(n829), .Q(
        \fpu_add_ctl/n746 ) );
  AO22X1 U4309 ( .IN1(n4364), .IN2(inq_op[0]), .IN3(n4365), .IN4(
        \fpu_add_ctl/n320 ), .Q(\fpu_add_ctl/n745 ) );
  NOR2X0 U4310 ( .IN1(n3986), .IN2(\fpu_add_ctl/n210 ), .QN(n4365) );
  AND2X1 U4311 ( .IN1(inq_add), .IN2(\fpu_add_ctl/n47 ), .Q(n4364) );
  AO22X1 U4312 ( .IN1(inq_fcc[1]), .IN2(n4366), .IN3(n1458), .IN4(n1011), .Q(
        \fpu_add_ctl/n744 ) );
  AO22X1 U4313 ( .IN1(inq_fcc[0]), .IN2(n4366), .IN3(n1457), .IN4(n1010), .Q(
        \fpu_add_ctl/n743 ) );
  AO22X1 U4314 ( .IN1(n1337), .IN2(n1010), .IN3(n1468), .IN4(n563), .Q(
        \fpu_add_ctl/n742 ) );
  AO22X1 U4315 ( .IN1(n1339), .IN2(n1011), .IN3(n1468), .IN4(n564), .Q(
        \fpu_add_ctl/n741 ) );
  AO22X1 U4316 ( .IN1(n1338), .IN2(n563), .IN3(n1468), .IN4(n1012), .Q(
        \fpu_add_ctl/n740 ) );
  AO22X1 U4317 ( .IN1(n1340), .IN2(n564), .IN3(n1468), .IN4(n1013), .Q(
        \fpu_add_ctl/n739 ) );
  AO22X1 U4318 ( .IN1(n1337), .IN2(n1012), .IN3(n1468), .IN4(n554), .Q(
        \fpu_add_ctl/n738 ) );
  AO22X1 U4319 ( .IN1(n1339), .IN2(n1013), .IN3(n1468), .IN4(n555), .Q(
        \fpu_add_ctl/n737 ) );
  AO22X1 U4320 ( .IN1(inq_id[4]), .IN2(n4366), .IN3(n1458), .IN4(n566), .Q(
        \fpu_add_ctl/n736 ) );
  AO22X1 U4321 ( .IN1(inq_id[3]), .IN2(n4366), .IN3(n1457), .IN4(n565), .Q(
        \fpu_add_ctl/n735 ) );
  AO22X1 U4322 ( .IN1(inq_id[2]), .IN2(n4366), .IN3(n1458), .IN4(n1216), .Q(
        \fpu_add_ctl/n734 ) );
  AO22X1 U4323 ( .IN1(inq_id[1]), .IN2(n4366), .IN3(n1457), .IN4(n1015), .Q(
        \fpu_add_ctl/n733 ) );
  AO22X1 U4324 ( .IN1(inq_id[0]), .IN2(n4366), .IN3(n1458), .IN4(n1014), .Q(
        \fpu_add_ctl/n732 ) );
  AO22X1 U4325 ( .IN1(n1338), .IN2(n1014), .IN3(n1468), .IN4(n567), .Q(
        \fpu_add_ctl/n731 ) );
  AO22X1 U4326 ( .IN1(n1340), .IN2(n1015), .IN3(n1468), .IN4(n568), .Q(
        \fpu_add_ctl/n730 ) );
  OAI22X1 U4327 ( .IN1(n4057), .IN2(\fpu_add_ctl/n183 ), .IN3(n4114), .IN4(
        \fpu_add_ctl/n182 ), .QN(\fpu_add_ctl/n729 ) );
  AO22X1 U4328 ( .IN1(n1337), .IN2(n565), .IN3(n1468), .IN4(n1016), .Q(
        \fpu_add_ctl/n728 ) );
  AO22X1 U4329 ( .IN1(n1339), .IN2(n566), .IN3(n1468), .IN4(n1017), .Q(
        \fpu_add_ctl/n727 ) );
  AO22X1 U4330 ( .IN1(n1338), .IN2(n567), .IN3(n1468), .IN4(n1018), .Q(
        \fpu_add_ctl/n726 ) );
  AO22X1 U4331 ( .IN1(n1340), .IN2(n568), .IN3(n1468), .IN4(n1019), .Q(
        \fpu_add_ctl/n725 ) );
  OAI22X1 U4332 ( .IN1(n4057), .IN2(\fpu_add_ctl/n182 ), .IN3(n4114), .IN4(
        \fpu_add_ctl/n326 ), .QN(\fpu_add_ctl/n724 ) );
  AO22X1 U4333 ( .IN1(n1337), .IN2(n1016), .IN3(n1468), .IN4(n269), .Q(
        \fpu_add_ctl/n723 ) );
  AO22X1 U4334 ( .IN1(n1339), .IN2(n1017), .IN3(n1469), .IN4(n89), .Q(
        \fpu_add_ctl/n722 ) );
  AO22X1 U4335 ( .IN1(n1338), .IN2(n1018), .IN3(n1469), .IN4(n342), .Q(
        \fpu_add_ctl/n721 ) );
  AO22X1 U4336 ( .IN1(n1340), .IN2(n1019), .IN3(n1469), .IN4(n341), .Q(
        \fpu_add_ctl/n720 ) );
  AO22X1 U4337 ( .IN1(n1472), .IN2(n354), .IN3(n4367), .IN4(\fpu_add_ctl/n308 ), .Q(\fpu_add_ctl/n719 ) );
  NOR2X0 U4338 ( .IN1(n4368), .IN2(n89), .QN(n4367) );
  AO22X1 U4339 ( .IN1(n1472), .IN2(n353), .IN3(n4369), .IN4(n4370), .Q(
        \fpu_add_ctl/n718 ) );
  NOR2X0 U4340 ( .IN1(n89), .IN2(n269), .QN(n4369) );
  AO22X1 U4341 ( .IN1(n1472), .IN2(n352), .IN3(n4371), .IN4(\fpu_add_ctl/n177 ), .Q(\fpu_add_ctl/n717 ) );
  NOR2X0 U4342 ( .IN1(\fpu_add_ctl/n308 ), .IN2(n4368), .QN(n4371) );
  AO22X1 U4343 ( .IN1(n1472), .IN2(n351), .IN3(n4372), .IN4(n4370), .Q(
        \fpu_add_ctl/n716 ) );
  NOR2X0 U4344 ( .IN1(\fpu_add_ctl/n308 ), .IN2(n89), .QN(n4372) );
  AO22X1 U4345 ( .IN1(n1472), .IN2(n350), .IN3(n4373), .IN4(\fpu_add_ctl/n308 ), .Q(\fpu_add_ctl/n715 ) );
  NOR2X0 U4346 ( .IN1(\fpu_add_ctl/n177 ), .IN2(n4368), .QN(n4373) );
  AO22X1 U4347 ( .IN1(n1472), .IN2(n349), .IN3(n4374), .IN4(n4370), .Q(
        \fpu_add_ctl/n714 ) );
  NOR2X0 U4348 ( .IN1(\fpu_add_ctl/n177 ), .IN2(n269), .QN(n4374) );
  AO22X1 U4349 ( .IN1(n4000), .IN2(n348), .IN3(n4375), .IN4(n4376), .Q(
        \fpu_add_ctl/n713 ) );
  INVX0 U4350 ( .INP(n4368), .ZN(n4376) );
  NAND2X0 U4351 ( .IN1(\fpu_add_ctl/n326 ), .IN2(n1337), .QN(n4368) );
  AO22X1 U4352 ( .IN1(n1472), .IN2(n347), .IN3(n4375), .IN4(n4370), .Q(
        \fpu_add_ctl/n712 ) );
  NOR2X0 U4353 ( .IN1(n4057), .IN2(\fpu_add_ctl/n326 ), .QN(n4370) );
  NOR2X0 U4354 ( .IN1(\fpu_add_ctl/n308 ), .IN2(\fpu_add_ctl/n177 ), .QN(n4375) );
  AO22X1 U4355 ( .IN1(n1337), .IN2(n342), .IN3(n1469), .IN4(n894), .Q(
        \fpu_add_ctl/n711 ) );
  AO22X1 U4356 ( .IN1(n1339), .IN2(n341), .IN3(n1469), .IN4(n893), .Q(
        \fpu_add_ctl/n710 ) );
  AO22X1 U4357 ( .IN1(n1338), .IN2(n354), .IN3(n1469), .IN4(n892), .Q(
        \fpu_add_ctl/n709 ) );
  AO22X1 U4358 ( .IN1(n1340), .IN2(n353), .IN3(n1469), .IN4(n891), .Q(
        \fpu_add_ctl/n708 ) );
  AO22X1 U4359 ( .IN1(n1337), .IN2(n352), .IN3(n1469), .IN4(n890), .Q(
        \fpu_add_ctl/n707 ) );
  AO22X1 U4360 ( .IN1(n1339), .IN2(n351), .IN3(n1469), .IN4(n889), .Q(
        \fpu_add_ctl/n706 ) );
  AO22X1 U4361 ( .IN1(n1338), .IN2(n350), .IN3(n1469), .IN4(n888), .Q(
        \fpu_add_ctl/n705 ) );
  AO22X1 U4362 ( .IN1(n1340), .IN2(n349), .IN3(n1469), .IN4(n887), .Q(
        \fpu_add_ctl/n704 ) );
  AO22X1 U4363 ( .IN1(n1337), .IN2(n348), .IN3(n1470), .IN4(n886), .Q(
        \fpu_add_ctl/n703 ) );
  AO22X1 U4364 ( .IN1(n1339), .IN2(n347), .IN3(n1470), .IN4(n885), .Q(
        \fpu_add_ctl/n702 ) );
  AO22X1 U4365 ( .IN1(inq_rnd_mode[1]), .IN2(n4366), .IN3(n1458), .IN4(n1021), 
        .Q(\fpu_add_ctl/n701 ) );
  AO22X1 U4366 ( .IN1(inq_rnd_mode[0]), .IN2(n4366), .IN3(n1458), .IN4(n1020), 
        .Q(\fpu_add_ctl/n700 ) );
  AO22X1 U4367 ( .IN1(n1338), .IN2(n1020), .IN3(n1470), .IN4(n505), .Q(
        \fpu_add_ctl/n699 ) );
  AO22X1 U4368 ( .IN1(n1340), .IN2(n1021), .IN3(n1470), .IN4(n504), .Q(
        \fpu_add_ctl/n698 ) );
  AO22X1 U4369 ( .IN1(n1337), .IN2(n505), .IN3(n1470), .IN4(n146), .Q(
        \fpu_add_ctl/n697 ) );
  AO22X1 U4370 ( .IN1(n1339), .IN2(n504), .IN3(n1470), .IN4(n147), .Q(
        \fpu_add_ctl/n696 ) );
  AO22X1 U4371 ( .IN1(n1338), .IN2(n146), .IN3(n1470), .IN4(n882), .Q(
        \fpu_add_ctl/n695 ) );
  AO22X1 U4372 ( .IN1(n1340), .IN2(n147), .IN3(n1470), .IN4(n883), .Q(
        \fpu_add_ctl/n694 ) );
  AO21X1 U4373 ( .IN1(n1457), .IN2(n915), .IN3(n4377), .Q(\fpu_add_ctl/n693 )
         );
  AO21X1 U4374 ( .IN1(n1457), .IN2(n325), .IN3(n4377), .Q(\fpu_add_ctl/n692 )
         );
  AO21X1 U4375 ( .IN1(n1457), .IN2(n44), .IN3(n4377), .Q(\fpu_add_ctl/n691 )
         );
  AO21X1 U4376 ( .IN1(n1457), .IN2(n700), .IN3(n4377), .Q(\fpu_add_ctl/n690 )
         );
  AO21X1 U4377 ( .IN1(n1457), .IN2(n295), .IN3(n4377), .Q(\fpu_add_ctl/n689 )
         );
  AND2X1 U4378 ( .IN1(n4366), .IN2(inq_op[1]), .Q(n4377) );
  AO21X1 U4379 ( .IN1(n1333), .IN2(n849), .IN3(n4378), .Q(\fpu_add_ctl/n688 )
         );
  AO21X1 U4380 ( .IN1(n1334), .IN2(n1001), .IN3(n4379), .Q(\fpu_add_ctl/n687 )
         );
  AO21X1 U4381 ( .IN1(n1335), .IN2(n560), .IN3(n4380), .Q(\fpu_add_ctl/n686 )
         );
  AO22X1 U4382 ( .IN1(n1333), .IN2(n570), .IN3(\fpu_add_ctl/n47 ), .IN4(n1658), 
        .Q(\fpu_add_ctl/n685 ) );
  INVX0 U4383 ( .INP(n4056), .ZN(n1658) );
  AO22X1 U4384 ( .IN1(n1335), .IN2(n571), .IN3(\fpu_add_ctl/n47 ), .IN4(n4381), 
        .Q(\fpu_add_ctl/n684 ) );
  NAND2X0 U4385 ( .IN1(n4070), .IN2(n4046), .QN(n4381) );
  NAND3X0 U4386 ( .IN1(n4382), .IN2(n4383), .IN3(n4384), .QN(
        \fpu_add_ctl/n683 ) );
  NAND2X0 U4387 ( .IN1(n1335), .IN2(n355), .QN(n4384) );
  INVX0 U4388 ( .INP(n4378), .ZN(n4383) );
  NOR2X0 U4389 ( .IN1(n4385), .IN2(\fpu_add_ctl/n312 ), .QN(n4378) );
  AO221X1 U4390 ( .IN1(\fpu_add_ctl/n47 ), .IN2(n2719), .IN3(n1336), .IN4(n858), .IN5(n4380), .Q(\fpu_add_ctl/n682 ) );
  AO22X1 U4391 ( .IN1(n1336), .IN2(n511), .IN3(n4386), .IN4(\fpu_add_ctl/n47 ), 
        .Q(\fpu_add_ctl/n681 ) );
  AO22X1 U4392 ( .IN1(n1334), .IN2(n757), .IN3(n4379), .IN4(n254), .Q(
        \fpu_add_ctl/n680 ) );
  AO22X1 U4393 ( .IN1(n1333), .IN2(n718), .IN3(n4380), .IN4(n158), .Q(
        \fpu_add_ctl/n679 ) );
  INVX0 U4394 ( .INP(n4387), .ZN(n4380) );
  AO22X1 U4395 ( .IN1(n1335), .IN2(n421), .IN3(n4379), .IN4(\fpu_add_ctl/n312 ), .Q(\fpu_add_ctl/n678 ) );
  INVX0 U4396 ( .INP(n4382), .ZN(n4379) );
  AO22X1 U4397 ( .IN1(n1336), .IN2(n128), .IN3(\fpu_add_ctl/n47 ), .IN4(n4388), 
        .Q(\fpu_add_ctl/n677 ) );
  NAND2X0 U4398 ( .IN1(n4070), .IN2(n4058), .QN(n4388) );
  INVX0 U4399 ( .INP(a1stg_fsdtoix), .ZN(n4058) );
  AO22X1 U4400 ( .IN1(n1334), .IN2(n1076), .IN3(n4072), .IN4(\fpu_add_ctl/n47 ), .Q(\fpu_add_ctl/n676 ) );
  NOR2X0 U4401 ( .IN1(n4389), .IN2(n4390), .QN(n4072) );
  AO22X1 U4402 ( .IN1(n1333), .IN2(n553), .IN3(\fpu_add_ctl/n47 ), .IN4(n4060), 
        .Q(\fpu_add_ctl/n675 ) );
  NOR2X0 U4403 ( .IN1(n4391), .IN2(n4390), .QN(n4060) );
  AO22X1 U4404 ( .IN1(n1335), .IN2(n569), .IN3(\fpu_add_ctl/n47 ), .IN4(n4068), 
        .Q(\fpu_add_ctl/n674 ) );
  NOR2X0 U4405 ( .IN1(n4392), .IN2(n4389), .QN(n4068) );
  AO22X1 U4406 ( .IN1(n1336), .IN2(n1022), .IN3(\fpu_add_ctl/n47 ), .IN4(n4069), .Q(\fpu_add_ctl/n673 ) );
  NOR2X0 U4407 ( .IN1(n4391), .IN2(n4392), .QN(n4069) );
  AO22X1 U4408 ( .IN1(n1334), .IN2(n258), .IN3(n4048), .IN4(\fpu_add_ctl/n47 ), 
        .Q(\fpu_add_ctl/n672 ) );
  AO22X1 U4409 ( .IN1(n1333), .IN2(n547), .IN3(n4393), .IN4(\fpu_add_ctl/n47 ), 
        .Q(\fpu_add_ctl/n671 ) );
  NOR2X0 U4410 ( .IN1(n4394), .IN2(n4392), .QN(n4393) );
  AO22X1 U4411 ( .IN1(n1335), .IN2(n1008), .IN3(n4395), .IN4(\fpu_add_ctl/n47 ), .Q(\fpu_add_ctl/n670 ) );
  NOR2X0 U4412 ( .IN1(n4394), .IN2(n4390), .QN(n4395) );
  AO22X1 U4413 ( .IN1(n1336), .IN2(n356), .IN3(\fpu_add_ctl/n47 ), .IN4(n2719), 
        .Q(\fpu_add_ctl/n669 ) );
  AO22X1 U4414 ( .IN1(n1334), .IN2(n1187), .IN3(\fpu_add_ctl/n47 ), .IN4(n4396), .Q(\fpu_add_ctl/n668 ) );
  AO22X1 U4415 ( .IN1(n1333), .IN2(n640), .IN3(\fpu_add_ctl/n47 ), .IN4(n1737), 
        .Q(\fpu_add_ctl/n667 ) );
  AO21X1 U4416 ( .IN1(n1336), .IN2(n1233), .IN3(n4397), .Q(\fpu_add_ctl/n666 )
         );
  AO21X1 U4417 ( .IN1(n1333), .IN2(n1218), .IN3(n4397), .Q(\fpu_add_ctl/n665 )
         );
  OAI21X1 U4418 ( .IN1(\fpu_add_ctl/n144 ), .IN2(n586), .IN3(n4398), .QN(
        \fpu_add_ctl/n664 ) );
  NAND4X0 U4419 ( .IN1(n4399), .IN2(\fpu_add_ctl/n318 ), .IN3(n4400), .IN4(
        n585), .QN(n4398) );
  AO22X1 U4420 ( .IN1(n1335), .IN2(n506), .IN3(\fpu_add_ctl/n47 ), .IN4(n2668), 
        .Q(\fpu_add_ctl/n663 ) );
  NAND3X0 U4421 ( .IN1(n4401), .IN2(n4382), .IN3(n4402), .QN(
        \fpu_add_ctl/n662 ) );
  OA22X1 U4422 ( .IN1(n4046), .IN2(n4403), .IN3(\fpu_add_ctl/n138 ), .IN4(n586), .Q(n4402) );
  NAND4X0 U4423 ( .IN1(n4404), .IN2(\fpu_add_ctl/n47 ), .IN3(n4405), .IN4(n158), .QN(n4382) );
  NAND4X0 U4424 ( .IN1(n4399), .IN2(\fpu_add_ctl/n303 ), .IN3(n18), .IN4(n158), 
        .QN(n4401) );
  AND3X1 U4425 ( .IN1(n4406), .IN2(\fpu_add_ctl/n314 ), .IN3(\fpu_add_ctl/n47 ), .Q(n4399) );
  NAND3X0 U4426 ( .IN1(n4387), .IN2(n4385), .IN3(n4407), .QN(
        \fpu_add_ctl/n661 ) );
  OA22X1 U4427 ( .IN1(n4056), .IN2(n4403), .IN3(\fpu_add_ctl/n113 ), .IN4(n586), .Q(n4407) );
  NAND2X0 U4428 ( .IN1(n4408), .IN2(n4409), .QN(n4056) );
  NAND4X0 U4429 ( .IN1(\fpu_add_ctl/n47 ), .IN2(n4410), .IN3(n4405), .IN4(n158), .QN(n4385) );
  NAND4X0 U4430 ( .IN1(\fpu_add_ctl/n47 ), .IN2(n4410), .IN3(n4405), .IN4(
        \fpu_add_ctl/n312 ), .QN(n4387) );
  AO22X1 U4431 ( .IN1(n1336), .IN2(n651), .IN3(\fpu_add_ctl/n47 ), .IN4(n4411), 
        .Q(\fpu_add_ctl/n660 ) );
  AO22X1 U4432 ( .IN1(n1334), .IN2(n1023), .IN3(\fpu_add_ctl/n47 ), .IN4(n295), 
        .Q(\fpu_add_ctl/n659 ) );
  AO22X1 U4433 ( .IN1(n1333), .IN2(n572), .IN3(\fpu_add_ctl/n49 ), .IN4(n849), 
        .Q(\fpu_add_ctl/n658 ) );
  AO22X1 U4434 ( .IN1(n1335), .IN2(n573), .IN3(\fpu_add_ctl/n49 ), .IN4(n1001), 
        .Q(\fpu_add_ctl/n657 ) );
  AO22X1 U4435 ( .IN1(n1336), .IN2(n1024), .IN3(\fpu_add_ctl/n49 ), .IN4(n560), 
        .Q(\fpu_add_ctl/n656 ) );
  AO22X1 U4436 ( .IN1(\fpu_add_ctl/a3stg_opdec_9_0[3] ), .IN2(n1336), .IN3(
        \fpu_add_ctl/n49 ), .IN4(n91), .Q(\fpu_add_ctl/n655 ) );
  AO22X1 U4437 ( .IN1(n1334), .IN2(n1025), .IN3(\fpu_add_ctl/n49 ), .IN4(n570), 
        .Q(\fpu_add_ctl/n654 ) );
  AO22X1 U4438 ( .IN1(n1333), .IN2(n1026), .IN3(\fpu_add_ctl/n49 ), .IN4(n562), 
        .Q(\fpu_add_ctl/n653 ) );
  AO22X1 U4439 ( .IN1(n1335), .IN2(n1027), .IN3(\fpu_add_ctl/n49 ), .IN4(n571), 
        .Q(\fpu_add_ctl/n652 ) );
  AO22X1 U4440 ( .IN1(n1336), .IN2(n895), .IN3(\fpu_add_ctl/n49 ), .IN4(n355), 
        .Q(\fpu_add_ctl/n651 ) );
  AO22X1 U4441 ( .IN1(n1334), .IN2(n455), .IN3(\fpu_add_ctl/n49 ), .IN4(n858), 
        .Q(\fpu_add_ctl/n650 ) );
  AO222X1 U4442 ( .IN1(n4412), .IN2(n146), .IN3(n4413), .IN4(n882), .IN5(n1461), .IN6(\fpu_add_ctl/n307 ), .Q(\fpu_add_ctl/n649 ) );
  AO222X1 U4443 ( .IN1(n4412), .IN2(n147), .IN3(n4413), .IN4(n883), .IN5(n1461), .IN6(n291), .Q(\fpu_add_ctl/n648 ) );
  AO22X1 U4444 ( .IN1(n1333), .IN2(n1028), .IN3(\fpu_add_ctl/n49 ), .IN4(n511), 
        .Q(\fpu_add_ctl/n647 ) );
  AO22X1 U4445 ( .IN1(n1335), .IN2(n336), .IN3(\fpu_add_ctl/n49 ), .IN4(
        \fpu_add_ctl/n329 ), .Q(\fpu_add_ctl/n646 ) );
  AO22X1 U4446 ( .IN1(n1336), .IN2(n1029), .IN3(\fpu_add_ctl/n49 ), .IN4(n356), 
        .Q(\fpu_add_ctl/n645 ) );
  AO21X1 U4447 ( .IN1(n1333), .IN2(n133), .IN3(n4397), .Q(\fpu_add_ctl/n644 )
         );
  AND2X1 U4448 ( .IN1(\fpu_add_ctl/n49 ), .IN2(n640), .Q(n4397) );
  AO22X1 U4449 ( .IN1(n1334), .IN2(n549), .IN3(\fpu_add_ctl/n49 ), .IN4(n1214), 
        .Q(\fpu_add_ctl/n643 ) );
  AO22X1 U4450 ( .IN1(n1333), .IN2(n1030), .IN3(\fpu_add_ctl/n49 ), .IN4(n506), 
        .Q(\fpu_add_ctl/n642 ) );
  AO22X1 U4451 ( .IN1(n1335), .IN2(n574), .IN3(\fpu_add_ctl/n49 ), .IN4(n1200), 
        .Q(\fpu_add_ctl/n641 ) );
  AO22X1 U4452 ( .IN1(n1336), .IN2(n575), .IN3(\fpu_add_ctl/n49 ), .IN4(n1201), 
        .Q(\fpu_add_ctl/n640 ) );
  AO22X1 U4453 ( .IN1(\fpu_add_ctl/n325 ), .IN2(n1334), .IN3(\fpu_add_ctl/n49 ), .IN4(n651), .Q(\fpu_add_ctl/n639 ) );
  AO22X1 U4454 ( .IN1(n1334), .IN2(n576), .IN3(\fpu_add_ctl/n49 ), .IN4(n1023), 
        .Q(\fpu_add_ctl/n638 ) );
  AO22X1 U4455 ( .IN1(n1333), .IN2(n1031), .IN3(\fpu_add_ctl/n49 ), .IN4(n572), 
        .Q(\fpu_add_ctl/n637 ) );
  AO22X1 U4456 ( .IN1(n1335), .IN2(n1032), .IN3(\fpu_add_ctl/n49 ), .IN4(n573), 
        .Q(\fpu_add_ctl/n636 ) );
  AO22X1 U4457 ( .IN1(n1336), .IN2(n492), .IN3(\fpu_add_ctl/n49 ), .IN4(n1024), 
        .Q(\fpu_add_ctl/n635 ) );
  AO22X1 U4458 ( .IN1(n1334), .IN2(n55), .IN3(\fpu_add_ctl/n49 ), .IN4(
        \fpu_add_ctl/a3stg_opdec_9_0[3] ), .Q(\fpu_add_ctl/n634 ) );
  AO22X1 U4459 ( .IN1(n1333), .IN2(n21), .IN3(\fpu_add_ctl/n49 ), .IN4(n1025), 
        .Q(\fpu_add_ctl/n633 ) );
  AO22X1 U4460 ( .IN1(n1335), .IN2(n148), .IN3(\fpu_add_ctl/n49 ), .IN4(n1026), 
        .Q(\fpu_add_ctl/n632 ) );
  AO22X1 U4461 ( .IN1(n1336), .IN2(n420), .IN3(\fpu_add_ctl/n49 ), .IN4(n1027), 
        .Q(\fpu_add_ctl/n631 ) );
  AO22X1 U4462 ( .IN1(\fpu_add_ctl/n319 ), .IN2(n1333), .IN3(\fpu_add_ctl/n49 ), .IN4(n895), .Q(\fpu_add_ctl/n630 ) );
  AO22X1 U4463 ( .IN1(n1334), .IN2(n324), .IN3(\fpu_add_ctl/n49 ), .IN4(n1028), 
        .Q(\fpu_add_ctl/n629 ) );
  AO22X1 U4464 ( .IN1(n1333), .IN2(n1246), .IN3(\fpu_add_ctl/n49 ), .IN4(n336), 
        .Q(\fpu_add_ctl/n628 ) );
  AO22X1 U4465 ( .IN1(n1335), .IN2(n490), .IN3(\fpu_add_ctl/n49 ), .IN4(n1029), 
        .Q(\fpu_add_ctl/n627 ) );
  AO22X1 U4466 ( .IN1(n1336), .IN2(n927), .IN3(\fpu_add_ctl/n49 ), .IN4(n133), 
        .Q(\fpu_add_ctl/n626 ) );
  AO22X1 U4467 ( .IN1(n1334), .IN2(n134), .IN3(\fpu_add_ctl/n49 ), .IN4(n549), 
        .Q(\fpu_add_ctl/n625 ) );
  AO22X1 U4468 ( .IN1(n1333), .IN2(n333), .IN3(\fpu_add_ctl/n49 ), .IN4(n1030), 
        .Q(\fpu_add_ctl/n624 ) );
  AO22X1 U4469 ( .IN1(n1335), .IN2(n135), .IN3(\fpu_add_ctl/n49 ), .IN4(n574), 
        .Q(\fpu_add_ctl/n623 ) );
  AO22X1 U4470 ( .IN1(n1336), .IN2(n136), .IN3(\fpu_add_ctl/n49 ), .IN4(n575), 
        .Q(\fpu_add_ctl/n622 ) );
  AO22X1 U4471 ( .IN1(n1334), .IN2(n339), .IN3(\fpu_add_ctl/n325 ), .IN4(
        \fpu_add_ctl/n49 ), .Q(\fpu_add_ctl/n621 ) );
  AO22X1 U4472 ( .IN1(n1333), .IN2(n108), .IN3(\fpu_add_ctl/n49 ), .IN4(n1031), 
        .Q(\fpu_add_ctl/n620 ) );
  AO22X1 U4473 ( .IN1(n1335), .IN2(n552), .IN3(\fpu_add_ctl/n49 ), .IN4(n1032), 
        .Q(\fpu_add_ctl/n619 ) );
  AO22X1 U4474 ( .IN1(n1336), .IN2(n622), .IN3(\fpu_add_ctl/n49 ), .IN4(
        \fpu_add_ctl/n319 ), .Q(\fpu_add_ctl/n618 ) );
  AO22X1 U4475 ( .IN1(n1334), .IN2(n1069), .IN3(\fpu_add_ctl/n49 ), .IN4(n324), 
        .Q(\fpu_add_ctl/n617 ) );
  AO22X1 U4476 ( .IN1(n1333), .IN2(n1070), .IN3(\fpu_add_ctl/n49 ), .IN4(n134), 
        .Q(\fpu_add_ctl/n616 ) );
  AO22X1 U4477 ( .IN1(n1335), .IN2(n1071), .IN3(\fpu_add_ctl/n49 ), .IN4(n333), 
        .Q(\fpu_add_ctl/n615 ) );
  AO22X1 U4478 ( .IN1(n1336), .IN2(n1072), .IN3(\fpu_add_ctl/n49 ), .IN4(n135), 
        .Q(\fpu_add_ctl/n614 ) );
  AO22X1 U4479 ( .IN1(n1334), .IN2(n1073), .IN3(\fpu_add_ctl/n49 ), .IN4(n136), 
        .Q(\fpu_add_ctl/n613 ) );
  AO22X1 U4480 ( .IN1(n1335), .IN2(n1157), .IN3(\fpu_add_ctl/n49 ), .IN4(n339), 
        .Q(\fpu_add_ctl/n612 ) );
  AO222X1 U4481 ( .IN1(n4414), .IN2(n1069), .IN3(n4415), .IN4(n324), .IN5(
        n1334), .IN6(a6stg_fcmpop), .Q(\fpu_add_ctl/n611 ) );
  AO222X1 U4482 ( .IN1(n4414), .IN2(n1070), .IN3(n4415), .IN4(n134), .IN5(
        n1333), .IN6(a6stg_int_dst), .Q(\fpu_add_ctl/n610 ) );
  AO222X1 U4483 ( .IN1(n4414), .IN2(n1071), .IN3(n4415), .IN4(n333), .IN5(
        n1336), .IN6(a6stg_long_dst), .Q(\fpu_add_ctl/n609 ) );
  AO222X1 U4484 ( .IN1(n4414), .IN2(n1072), .IN3(n4415), .IN4(n135), .IN5(
        n1335), .IN6(a6stg_sng_dst), .Q(\fpu_add_ctl/n608 ) );
  AO222X1 U4485 ( .IN1(n4414), .IN2(n1073), .IN3(n4415), .IN4(n136), .IN5(
        n1334), .IN6(a6stg_dbl_dst), .Q(\fpu_add_ctl/n607 ) );
  AND3X1 U4486 ( .IN1(\fpu_add_ctl/n315 ), .IN2(n642), .IN3(\fpu_add_ctl/n49 ), 
        .Q(n4415) );
  AND2X1 U4487 ( .IN1(\fpu_add_ctl/n49 ), .IN2(n622), .Q(n4414) );
  AO22X1 U4488 ( .IN1(n1336), .IN2(n1242), .IN3(\fpu_add_ctl/n49 ), .IN4(n576), 
        .Q(\fpu_add_ctl/n606 ) );
  AO21X1 U4489 ( .IN1(n1457), .IN2(n129), .IN3(n4416), .Q(\fpu_add_ctl/n605 )
         );
  AO21X1 U4490 ( .IN1(n1457), .IN2(n692), .IN3(n4416), .Q(\fpu_add_ctl/n604 )
         );
  AO21X1 U4491 ( .IN1(n1457), .IN2(n102), .IN3(n4416), .Q(\fpu_add_ctl/n603 )
         );
  AO21X1 U4492 ( .IN1(n1457), .IN2(n701), .IN3(n4416), .Q(\fpu_add_ctl/n602 )
         );
  AO21X1 U4493 ( .IN1(n1457), .IN2(n662), .IN3(n4416), .Q(\fpu_add_ctl/n601 )
         );
  AND2X1 U4494 ( .IN1(n4366), .IN2(inq_op[0]), .Q(n4416) );
  AO22X1 U4495 ( .IN1(inq_in2_exp_neq_ffs), .IN2(n4366), .IN3(n1459), .IN4(
        \fpu_add_ctl/n317 ), .Q(\fpu_add_ctl/n600 ) );
  AO22X1 U4496 ( .IN1(inq_in2_exp_eq_0), .IN2(n4366), .IN3(n1458), .IN4(n1086), 
        .Q(\fpu_add_ctl/n599 ) );
  AO22X1 U4497 ( .IN1(inq_in2_53_32_neq_0), .IN2(n4366), .IN3(n1459), .IN4(
        n730), .Q(\fpu_add_ctl/n598 ) );
  AO22X1 U4498 ( .IN1(inq_in2_50_0_neq_0), .IN2(n4366), .IN3(n1458), .IN4(n731), .Q(\fpu_add_ctl/n597 ) );
  AO22X1 U4499 ( .IN1(n4366), .IN2(inq_in2[63]), .IN3(n1459), .IN4(n649), .Q(
        \fpu_add_ctl/n596 ) );
  AO22X1 U4500 ( .IN1(n4366), .IN2(inq_in2[54]), .IN3(n1458), .IN4(n847), .Q(
        \fpu_add_ctl/n595 ) );
  AO22X1 U4501 ( .IN1(n4366), .IN2(inq_in2[51]), .IN3(n1459), .IN4(n460), .Q(
        \fpu_add_ctl/n594 ) );
  AO22X1 U4502 ( .IN1(inq_in1_exp_neq_ffs), .IN2(n4366), .IN3(n1458), .IN4(
        n598), .Q(\fpu_add_ctl/n593 ) );
  AO22X1 U4503 ( .IN1(inq_in1_exp_eq_0), .IN2(n4366), .IN3(n1459), .IN4(n1085), 
        .Q(\fpu_add_ctl/n592 ) );
  AO22X1 U4504 ( .IN1(inq_in1_53_32_neq_0), .IN2(n4366), .IN3(n1458), .IN4(
        n743), .Q(\fpu_add_ctl/n591 ) );
  AO22X1 U4505 ( .IN1(inq_in1_50_0_neq_0), .IN2(n4366), .IN3(n1459), .IN4(n744), .Q(\fpu_add_ctl/n590 ) );
  AO22X1 U4506 ( .IN1(inq_in1[63]), .IN2(n4366), .IN3(n1458), .IN4(n897), .Q(
        \fpu_add_ctl/n589 ) );
  AO22X1 U4507 ( .IN1(n4366), .IN2(inq_in1[54]), .IN3(n1459), .IN4(n1120), .Q(
        \fpu_add_ctl/n588 ) );
  AO22X1 U4508 ( .IN1(n4366), .IN2(inq_in1[51]), .IN3(n1458), .IN4(n1119), .Q(
        \fpu_add_ctl/n587 ) );
  NAND2X0 U4509 ( .IN1(n4417), .IN2(\fpu_add_ctl/n470 ), .QN(n3986) );
  AND2X1 U4510 ( .IN1(n1338), .IN2(n4418), .Q(n4366) );
  AO22X1 U4511 ( .IN1(n1472), .IN2(add_fcc_out[0]), .IN3(n4419), .IN4(n554), 
        .Q(\fpu_add_ctl/n586 ) );
  AO22X1 U4512 ( .IN1(n4000), .IN2(add_fcc_out[1]), .IN3(n4419), .IN4(n555), 
        .Q(\fpu_add_ctl/n585 ) );
  AO22X1 U4513 ( .IN1(n1337), .IN2(n897), .IN3(n1471), .IN4(n433), .Q(
        \fpu_add_ctl/n584 ) );
  AO22X1 U4514 ( .IN1(n1339), .IN2(n649), .IN3(n1471), .IN4(n270), .Q(
        \fpu_add_ctl/n583 ) );
  AO22X1 U4515 ( .IN1(n1338), .IN2(n1656), .IN3(n1470), .IN4(
        \fpu_add_ctl/n313 ), .Q(\fpu_add_ctl/n582 ) );
  AO22X1 U4516 ( .IN1(n1340), .IN2(n4420), .IN3(n1470), .IN4(n1210), .Q(
        \fpu_add_ctl/n581 ) );
  NAND4X0 U4517 ( .IN1(n4421), .IN2(n4422), .IN3(n4423), .IN4(n4424), .QN(
        n4420) );
  NOR4X0 U4518 ( .IN1(n4425), .IN2(n4426), .IN3(n4427), .IN4(n4428), .QN(n4424) );
  XOR2X1 U4519 ( .IN1(\fpu_add_frac_dp/n2493 ), .IN2(n702), .Q(n4427) );
  NOR2X0 U4520 ( .IN1(n4429), .IN2(n4430), .QN(n4423) );
  AO22X1 U4521 ( .IN1(n1337), .IN2(n1881), .IN3(n1469), .IN4(n1212), .Q(
        \fpu_add_ctl/n580 ) );
  OAI21X1 U4522 ( .IN1(n4425), .IN2(n4431), .IN3(n4432), .QN(n1881) );
  NAND4X0 U4523 ( .IN1(n4433), .IN2(n4434), .IN3(n4435), .IN4(n662), .QN(n4432) );
  OR3X1 U4524 ( .IN1(n4436), .IN2(\fpu_add_frac_dp/n900 ), .IN3(n650), .Q(
        n4434) );
  NAND2X0 U4525 ( .IN1(\fpu_add_frac_dp/n2364 ), .IN2(n283), .QN(n4433) );
  MUX21X1 U4526 ( .IN1(n4437), .IN2(n4438), .S(n4421), .Q(n4431) );
  AND4X1 U4527 ( .IN1(n4439), .IN2(n4440), .IN3(n4441), .IN4(n4442), .Q(n4421)
         );
  NOR4X0 U4528 ( .IN1(n4443), .IN2(n4444), .IN3(n4445), .IN4(n4446), .QN(n4442) );
  INVX0 U4529 ( .INP(n4447), .ZN(n4444) );
  OR3X1 U4530 ( .IN1(n4448), .IN2(n4449), .IN3(n4450), .Q(n4443) );
  OA221X1 U4531 ( .IN1(n428), .IN2(n54), .IN3(n989), .IN4(n132), .IN5(n4451), 
        .Q(n4441) );
  OA21X1 U4532 ( .IN1(n1067), .IN2(n326), .IN3(n4452), .Q(n4451) );
  NOR2X0 U4533 ( .IN1(n4453), .IN2(n4454), .QN(n4439) );
  XOR2X1 U4534 ( .IN1(n647), .IN2(\fpu_add_frac_dp/n5608 ), .Q(n4453) );
  MUX21X1 U4535 ( .IN1(n4455), .IN2(n4456), .S(n4422), .Q(n4438) );
  AND4X1 U4536 ( .IN1(n4457), .IN2(n4458), .IN3(n4459), .IN4(n4460), .Q(n4422)
         );
  NOR4X0 U4537 ( .IN1(n4461), .IN2(n4462), .IN3(n4463), .IN4(n4464), .QN(n4460) );
  XOR2X1 U4538 ( .IN1(\fpu_add_frac_dp/n846 ), .IN2(\fpu_add_frac_dp/n2439 ), 
        .Q(n4464) );
  INVX0 U4539 ( .INP(n4465), .ZN(n4461) );
  AOI221X1 U4540 ( .IN1(\fpu_add_frac_dp/n2487 ), .IN2(\fpu_add_frac_dp/n921 ), 
        .IN3(\fpu_add_frac_dp/n2444 ), .IN4(\fpu_add_frac_dp/n845 ), .IN5(
        n4466), .QN(n4459) );
  MUX21X1 U4541 ( .IN1(n4467), .IN2(n4468), .S(n4430), .Q(n4456) );
  NAND4X0 U4542 ( .IN1(n4469), .IN2(n4470), .IN3(n4471), .IN4(n4472), .QN(
        n4430) );
  NAND2X0 U4543 ( .IN1(\fpu_add_frac_dp/n928 ), .IN2(\fpu_add_frac_dp/n2483 ), 
        .QN(n4472) );
  INVX0 U4544 ( .INP(n4473), .ZN(n4471) );
  XOR2X1 U4545 ( .IN1(n697), .IN2(\fpu_add_frac_dp/n2544 ), .Q(n4469) );
  OA221X1 U4546 ( .IN1(n4474), .IN2(n4475), .IN3(n4476), .IN4(n4477), .IN5(
        n4478), .Q(n4468) );
  OA22X1 U4547 ( .IN1(n4479), .IN2(n4480), .IN3(\fpu_add_frac_dp/n2536 ), 
        .IN4(n853), .Q(n4478) );
  NOR2X0 U4548 ( .IN1(n4481), .IN2(n4482), .QN(n4476) );
  NOR3X0 U4549 ( .IN1(n4483), .IN2(\fpu_add_frac_dp/n848 ), .IN3(
        \fpu_add_frac_dp/n2484 ), .QN(n4481) );
  INVX0 U4550 ( .INP(n4470), .ZN(n4475) );
  NOR4X0 U4551 ( .IN1(n4477), .IN2(n4482), .IN3(n4484), .IN4(n4483), .QN(n4470) );
  NOR2X0 U4552 ( .IN1(n330), .IN2(\fpu_add_frac_dp/n2368 ), .QN(n4483) );
  XOR2X1 U4553 ( .IN1(n670), .IN2(\fpu_add_frac_dp/n2484 ), .Q(n4484) );
  AO22X1 U4554 ( .IN1(\fpu_add_frac_dp/n2454 ), .IN2(n1007), .IN3(
        \fpu_add_frac_dp/n2368 ), .IN4(n330), .Q(n4482) );
  NAND3X0 U4555 ( .IN1(n4485), .IN2(n4479), .IN3(n4486), .QN(n4477) );
  AOI22X1 U4556 ( .IN1(\fpu_add_frac_dp/n2453 ), .IN2(\fpu_add_frac_dp/n847 ), 
        .IN3(n988), .IN4(\fpu_add_frac_dp/n5627 ), .QN(n4486) );
  OA22X1 U4557 ( .IN1(\fpu_add_frac_dp/n2453 ), .IN2(\fpu_add_frac_dp/n847 ), 
        .IN3(n703), .IN4(\fpu_add_frac_dp/n5629 ), .Q(n4479) );
  INVX0 U4558 ( .INP(n4480), .ZN(n4485) );
  AO21X1 U4559 ( .IN1(\fpu_add_frac_dp/n5629 ), .IN2(n703), .IN3(n4487), .Q(
        n4480) );
  XOR2X1 U4560 ( .IN1(\fpu_add_frac_dp/n2536 ), .IN2(\fpu_add_frac_dp/n2372 ), 
        .Q(n4487) );
  OA22X1 U4561 ( .IN1(n4488), .IN2(n4473), .IN3(n357), .IN4(n854), .Q(n4474)
         );
  AO21X1 U4562 ( .IN1(n1088), .IN2(n145), .IN3(n4489), .Q(n4473) );
  XOR2X1 U4563 ( .IN1(n357), .IN2(\fpu_add_frac_dp/n927 ), .Q(n4489) );
  OA21X1 U4564 ( .IN1(n1088), .IN2(n145), .IN3(n577), .Q(n4488) );
  NOR4X0 U4565 ( .IN1(n4490), .IN2(n4491), .IN3(n4492), .IN4(n4493), .QN(n4467) );
  AND2X1 U4566 ( .IN1(\fpu_add_frac_dp/n2472 ), .IN2(\fpu_add_frac_dp/n929 ), 
        .Q(n4493) );
  OA221X1 U4567 ( .IN1(\fpu_add_frac_dp/n932 ), .IN2(\fpu_add_frac_dp/n2459 ), 
        .IN3(n4494), .IN4(n4495), .IN5(n4496), .Q(n4492) );
  AOI21X1 U4568 ( .IN1(n695), .IN2(\fpu_add_frac_dp/n2366 ), .IN3(n4497), .QN(
        n4495) );
  OA21X1 U4569 ( .IN1(n4498), .IN2(n4499), .IN3(n4500), .Q(n4491) );
  INVX0 U4570 ( .INP(n4501), .ZN(n4499) );
  AND2X1 U4571 ( .IN1(\fpu_add_frac_dp/n2490 ), .IN2(\fpu_add_frac_dp/n931 ), 
        .Q(n4498) );
  OA221X1 U4572 ( .IN1(n4502), .IN2(n4428), .IN3(n4503), .IN4(n4504), .IN5(
        n4505), .Q(n4490) );
  INVX0 U4573 ( .INP(n4429), .ZN(n4505) );
  NAND4X0 U4574 ( .IN1(n4496), .IN2(n4506), .IN3(n4497), .IN4(n4507), .QN(
        n4429) );
  OA221X1 U4575 ( .IN1(\fpu_add_frac_dp/n934 ), .IN2(n337), .IN3(
        \fpu_add_frac_dp/n933 ), .IN4(n900), .IN5(n4508), .Q(n4507) );
  AOI21X1 U4576 ( .IN1(\fpu_add_frac_dp/n2296 ), .IN2(\fpu_add_frac_dp/n2533 ), 
        .IN3(n4494), .QN(n4508) );
  AND2X1 U4577 ( .IN1(\fpu_add_frac_dp/n932 ), .IN2(\fpu_add_frac_dp/n2459 ), 
        .Q(n4494) );
  OA22X1 U4578 ( .IN1(n695), .IN2(\fpu_add_frac_dp/n2366 ), .IN3(
        \fpu_add_frac_dp/n2533 ), .IN4(\fpu_add_frac_dp/n2296 ), .Q(n4497) );
  OR2X1 U4579 ( .IN1(\fpu_add_frac_dp/n2459 ), .IN2(\fpu_add_frac_dp/n932 ), 
        .Q(n4506) );
  AND4X1 U4580 ( .IN1(n4500), .IN2(n4509), .IN3(n4510), .IN4(n4501), .Q(n4496)
         );
  NAND2X0 U4581 ( .IN1(\fpu_add_frac_dp/n930 ), .IN2(\fpu_add_frac_dp/n2489 ), 
        .QN(n4501) );
  NAND2X0 U4582 ( .IN1(\fpu_add_frac_dp/n929 ), .IN2(\fpu_add_frac_dp/n2472 ), 
        .QN(n4510) );
  XOR2X1 U4583 ( .IN1(\fpu_add_frac_dp/n931 ), .IN2(\fpu_add_frac_dp/n2490 ), 
        .Q(n4509) );
  OA22X1 U4584 ( .IN1(\fpu_add_frac_dp/n2489 ), .IN2(\fpu_add_frac_dp/n930 ), 
        .IN3(\fpu_add_frac_dp/n2472 ), .IN4(\fpu_add_frac_dp/n929 ), .Q(n4500)
         );
  INVX0 U4585 ( .INP(n4426), .ZN(n4504) );
  NOR2X0 U4586 ( .IN1(\fpu_add_frac_dp/n2455 ), .IN2(\fpu_add_frac_dp/n935 ), 
        .QN(n4426) );
  NOR2X0 U4587 ( .IN1(\fpu_add_frac_dp/n2436 ), .IN2(n745), .QN(n4503) );
  AO22X1 U4588 ( .IN1(\fpu_add_frac_dp/n935 ), .IN2(\fpu_add_frac_dp/n2455 ), 
        .IN3(\fpu_add_frac_dp/n934 ), .IN4(n337), .Q(n4428) );
  NOR2X0 U4589 ( .IN1(\fpu_add_frac_dp/n2493 ), .IN2(\fpu_add_frac_dp/n851 ), 
        .QN(n4502) );
  OA21X1 U4590 ( .IN1(n1303), .IN2(n550), .IN3(n4511), .Q(n4455) );
  NAND3X0 U4591 ( .IN1(n4512), .IN2(n4513), .IN3(n4458), .QN(n4511) );
  OA21X1 U4592 ( .IN1(\fpu_add_frac_dp/n2486 ), .IN2(\fpu_add_frac_dp/n918 ), 
        .IN3(n4514), .Q(n4458) );
  XOR2X1 U4593 ( .IN1(\fpu_add_frac_dp/n2482 ), .IN2(\fpu_add_frac_dp/n917 ), 
        .Q(n4514) );
  NAND3X0 U4594 ( .IN1(n4515), .IN2(n4516), .IN3(n4517), .QN(n4513) );
  INVX0 U4595 ( .INP(n4462), .ZN(n4517) );
  NAND2X0 U4596 ( .IN1(n4518), .IN2(n4519), .QN(n4462) );
  XOR2X1 U4597 ( .IN1(\fpu_add_frac_dp/n844 ), .IN2(\fpu_add_frac_dp/n2488 ), 
        .Q(n4518) );
  OAI21X1 U4598 ( .IN1(n4520), .IN2(n4463), .IN3(n4457), .QN(n4515) );
  OA221X1 U4599 ( .IN1(\fpu_add_frac_dp/n2458 ), .IN2(\fpu_add_frac_dp/n919 ), 
        .IN3(\fpu_add_frac_dp/n2492 ), .IN4(\fpu_add_frac_dp/n920 ), .IN5(
        n4516), .Q(n4457) );
  NAND2X0 U4600 ( .IN1(\fpu_add_frac_dp/n919 ), .IN2(\fpu_add_frac_dp/n2458 ), 
        .QN(n4516) );
  AO22X1 U4601 ( .IN1(\fpu_add_frac_dp/n920 ), .IN2(\fpu_add_frac_dp/n2492 ), 
        .IN3(n335), .IN4(n1078), .Q(n4463) );
  OA22X1 U4602 ( .IN1(n4521), .IN2(n4522), .IN3(n1078), .IN4(n335), .Q(n4520)
         );
  AND2X1 U4603 ( .IN1(\fpu_add_frac_dp/n2487 ), .IN2(\fpu_add_frac_dp/n921 ), 
        .Q(n4522) );
  OA21X1 U4604 ( .IN1(\fpu_add_frac_dp/n2439 ), .IN2(n4466), .IN3(n4465), .Q(
        n4521) );
  OA22X1 U4605 ( .IN1(\fpu_add_frac_dp/n2487 ), .IN2(\fpu_add_frac_dp/n921 ), 
        .IN3(\fpu_add_frac_dp/n2485 ), .IN4(\fpu_add_frac_dp/n922 ), .Q(n4465)
         );
  AND2X1 U4606 ( .IN1(\fpu_add_frac_dp/n922 ), .IN2(\fpu_add_frac_dp/n2485 ), 
        .Q(n4466) );
  NAND3X0 U4607 ( .IN1(\fpu_add_frac_dp/n2488 ), .IN2(n4519), .IN3(
        \fpu_add_frac_dp/n844 ), .QN(n4512) );
  NAND2X0 U4608 ( .IN1(\fpu_add_frac_dp/n918 ), .IN2(\fpu_add_frac_dp/n2486 ), 
        .QN(n4519) );
  OA221X1 U4609 ( .IN1(n1089), .IN2(n340), .IN3(n4448), .IN4(n4523), .IN5(
        n4524), .Q(n4437) );
  NAND3X0 U4610 ( .IN1(n1158), .IN2(n427), .IN3(n4525), .QN(n4524) );
  MUX21X1 U4611 ( .IN1(n4526), .IN2(n4527), .S(n4450), .Q(n4523) );
  NAND4X0 U4612 ( .IN1(n4528), .IN2(n4529), .IN3(n4530), .IN4(n4531), .QN(
        n4450) );
  NOR2X0 U4613 ( .IN1(n4532), .IN2(n4533), .QN(n4530) );
  XOR2X1 U4614 ( .IN1(n677), .IN2(\fpu_add_frac_dp/n2538 ), .Q(n4528) );
  AO22X1 U4615 ( .IN1(n4533), .IN2(n4534), .IN3(n4535), .IN4(n4531), .Q(n4527)
         );
  OA21X1 U4616 ( .IN1(\fpu_add_frac_dp/n5626 ), .IN2(\fpu_add_frac_dp/n2476 ), 
        .IN3(n4534), .Q(n4531) );
  OA21X1 U4617 ( .IN1(n4536), .IN2(n4537), .IN3(n4538), .Q(n4535) );
  INVX0 U4618 ( .INP(n4529), .ZN(n4537) );
  OA221X1 U4619 ( .IN1(\fpu_add_frac_dp/n904 ), .IN2(\fpu_add_frac_dp/n5611 ), 
        .IN3(\fpu_add_frac_dp/n903 ), .IN4(\fpu_add_frac_dp/n5624 ), .IN5(
        n4538), .Q(n4529) );
  NAND2X0 U4620 ( .IN1(\fpu_add_frac_dp/n903 ), .IN2(\fpu_add_frac_dp/n5624 ), 
        .QN(n4538) );
  NOR2X0 U4621 ( .IN1(\fpu_add_frac_dp/n2373 ), .IN2(n4532), .QN(n4536) );
  AND2X1 U4622 ( .IN1(\fpu_add_frac_dp/n904 ), .IN2(\fpu_add_frac_dp/n5611 ), 
        .Q(n4532) );
  NAND2X0 U4623 ( .IN1(\fpu_add_frac_dp/n2415 ), .IN2(n1065), .QN(n4534) );
  AO22X1 U4624 ( .IN1(\fpu_add_frac_dp/n5626 ), .IN2(\fpu_add_frac_dp/n2476 ), 
        .IN3(\fpu_add_frac_dp/n5625 ), .IN4(n917), .Q(n4533) );
  MUX21X1 U4625 ( .IN1(n4539), .IN2(n4540), .S(n4445), .Q(n4526) );
  NAND3X0 U4626 ( .IN1(n4541), .IN2(n4542), .IN3(n4543), .QN(n4445) );
  OA22X1 U4627 ( .IN1(n719), .IN2(n125), .IN3(n306), .IN4(n46), .Q(n4543) );
  INVX0 U4628 ( .INP(n4544), .ZN(n4542) );
  XOR2X1 U4629 ( .IN1(n292), .IN2(\fpu_add_frac_dp/n841 ), .Q(n4541) );
  AND3X1 U4630 ( .IN1(n4545), .IN2(n4546), .IN3(n4547), .Q(n4540) );
  OA22X1 U4631 ( .IN1(n4548), .IN2(n4544), .IN3(n578), .IN4(n57), .Q(n4547) );
  AO221X1 U4632 ( .IN1(n125), .IN2(n719), .IN3(n46), .IN4(n306), .IN5(n4549), 
        .Q(n4544) );
  OA21X1 U4633 ( .IN1(n719), .IN2(n125), .IN3(n292), .Q(n4548) );
  OR3X1 U4634 ( .IN1(n4550), .IN2(n4551), .IN3(n4552), .Q(n4546) );
  AND2X1 U4635 ( .IN1(n4553), .IN2(n4554), .Q(n4552) );
  NAND3X0 U4636 ( .IN1(n4555), .IN2(n4556), .IN3(n4557), .QN(n4554) );
  AO22X1 U4637 ( .IN1(\fpu_add_frac_dp/n907 ), .IN2(\fpu_add_frac_dp/n5620 ), 
        .IN3(n4558), .IN4(n4559), .Q(n4557) );
  INVX0 U4638 ( .INP(n4560), .ZN(n4559) );
  NAND2X0 U4639 ( .IN1(\fpu_add_frac_dp/n2438 ), .IN2(n709), .QN(n4558) );
  OR3X1 U4640 ( .IN1(n4549), .IN2(n306), .IN3(n46), .Q(n4545) );
  NAND4X0 U4641 ( .IN1(n4561), .IN2(n4553), .IN3(n4562), .IN4(n4563), .QN(
        n4549) );
  NOR4X0 U4642 ( .IN1(n4564), .IN2(n4560), .IN3(n4551), .IN4(n4565), .QN(n4563) );
  INVX0 U4643 ( .INP(n4555), .ZN(n4565) );
  NAND2X0 U4644 ( .IN1(\fpu_add_frac_dp/n839 ), .IN2(\fpu_add_frac_dp/n2462 ), 
        .QN(n4555) );
  NOR2X0 U4645 ( .IN1(\fpu_add_frac_dp/n905 ), .IN2(\fpu_add_frac_dp/n5621 ), 
        .QN(n4551) );
  NOR2X0 U4646 ( .IN1(\fpu_add_frac_dp/n907 ), .IN2(\fpu_add_frac_dp/n5620 ), 
        .QN(n4560) );
  AO21X1 U4647 ( .IN1(\fpu_add_frac_dp/n2438 ), .IN2(n709), .IN3(n4550), .Q(
        n4564) );
  NOR2X0 U4648 ( .IN1(n763), .IN2(\fpu_add_frac_dp/n2540 ), .QN(n4550) );
  OA22X1 U4649 ( .IN1(n1079), .IN2(n141), .IN3(n578), .IN4(n57), .Q(n4562) );
  OA22X1 U4650 ( .IN1(n848), .IN2(\fpu_add_frac_dp/n2543 ), .IN3(
        \fpu_add_frac_dp/n2462 ), .IN4(\fpu_add_frac_dp/n839 ), .Q(n4553) );
  INVX0 U4651 ( .INP(n4556), .ZN(n4561) );
  AO222X1 U4652 ( .IN1(n1079), .IN2(n141), .IN3(\fpu_add_frac_dp/n908 ), .IN4(
        n463), .IN5(\fpu_add_frac_dp/n907 ), .IN6(\fpu_add_frac_dp/n5620 ), 
        .Q(n4556) );
  OA21X1 U4653 ( .IN1(n4566), .IN2(n4454), .IN3(n4452), .Q(n4539) );
  NAND2X0 U4654 ( .IN1(\fpu_add_frac_dp/n911 ), .IN2(\fpu_add_frac_dp/n5623 ), 
        .QN(n4452) );
  OAI22X1 U4655 ( .IN1(\fpu_add_frac_dp/n5623 ), .IN2(\fpu_add_frac_dp/n911 ), 
        .IN3(n916), .IN4(\fpu_add_frac_dp/n912 ), .QN(n4454) );
  OA21X1 U4656 ( .IN1(n4567), .IN2(n4568), .IN3(n4447), .Q(n4566) );
  OA22X1 U4657 ( .IN1(n857), .IN2(\fpu_add_frac_dp/n2365 ), .IN3(
        \fpu_add_frac_dp/n2295 ), .IN4(\fpu_add_frac_dp/n2532 ), .Q(n4447) );
  NOR2X0 U4658 ( .IN1(n1067), .IN2(n326), .QN(n4568) );
  OA22X1 U4659 ( .IN1(n4569), .IN2(n4446), .IN3(n358), .IN4(n855), .Q(n4567)
         );
  AO21X1 U4660 ( .IN1(\fpu_add_frac_dp/n2441 ), .IN2(n704), .IN3(n4570), .Q(
        n4446) );
  XOR2X1 U4661 ( .IN1(n358), .IN2(\fpu_add_frac_dp/n913 ), .Q(n4570) );
  OA21X1 U4662 ( .IN1(n4571), .IN2(n4572), .IN3(n4440), .Q(n4569) );
  OA22X1 U4663 ( .IN1(\fpu_add_frac_dp/n2445 ), .IN2(\fpu_add_frac_dp/n843 ), 
        .IN3(n704), .IN4(\fpu_add_frac_dp/n2441 ), .Q(n4440) );
  NOR2X0 U4664 ( .IN1(n989), .IN2(n132), .QN(n4572) );
  OA22X1 U4665 ( .IN1(n4573), .IN2(n4449), .IN3(\fpu_add_frac_dp/n2514 ), 
        .IN4(n856), .Q(n4571) );
  AO21X1 U4666 ( .IN1(n428), .IN2(n54), .IN3(n4574), .Q(n4449) );
  XOR2X1 U4667 ( .IN1(\fpu_add_frac_dp/n2514 ), .IN2(\fpu_add_frac_dp/n2367 ), 
        .Q(n4574) );
  OA21X1 U4668 ( .IN1(n428), .IN2(n54), .IN3(n647), .Q(n4573) );
  NAND3X0 U4669 ( .IN1(n4575), .IN2(n4525), .IN3(n4576), .QN(n4448) );
  XOR2X1 U4670 ( .IN1(\fpu_add_frac_dp/n2535 ), .IN2(\fpu_add_frac_dp/n2350 ), 
        .Q(n4576) );
  NAND2X0 U4671 ( .IN1(n340), .IN2(n1089), .QN(n4525) );
  NAND2X0 U4672 ( .IN1(\fpu_add_frac_dp/n901 ), .IN2(\fpu_add_frac_dp/n2491 ), 
        .QN(n4575) );
  AND2X1 U4673 ( .IN1(n4577), .IN2(n662), .Q(n4425) );
  AO221X1 U4674 ( .IN1(\fpu_add_frac_dp/n2364 ), .IN2(n283), .IN3(
        \fpu_add_frac_dp/n2442 ), .IN4(n747), .IN5(n4578), .Q(n4577) );
  AO21X1 U4675 ( .IN1(n548), .IN2(n1304), .IN3(n4435), .Q(n4578) );
  AO221X1 U4676 ( .IN1(\fpu_add_frac_dp/n900 ), .IN2(n650), .IN3(
        \fpu_add_frac_dp/n5643 ), .IN4(\fpu_add_frac_dp/n5644 ), .IN5(n4436), 
        .Q(n4435) );
  NOR2X0 U4677 ( .IN1(n283), .IN2(\fpu_add_frac_dp/n2364 ), .QN(n4436) );
  AO22X1 U4678 ( .IN1(n1339), .IN2(n1880), .IN3(n1470), .IN4(n1004), .Q(
        \fpu_add_ctl/n579 ) );
  AND4X1 U4679 ( .IN1(n4579), .IN2(n4580), .IN3(n4581), .IN4(n4582), .Q(n1880)
         );
  NOR4X0 U4680 ( .IN1(n4583), .IN2(n4584), .IN3(n4585), .IN4(n4586), .QN(n4582) );
  XOR2X1 U4681 ( .IN1(\fpu_add_frac_dp/n2475 ), .IN2(n712), .Q(n4586) );
  XOR2X1 U4682 ( .IN1(\fpu_add_frac_dp/n2467 ), .IN2(n713), .Q(n4585) );
  XOR2X1 U4683 ( .IN1(\fpu_add_frac_dp/n2466 ), .IN2(n714), .Q(n4584) );
  XOR2X1 U4684 ( .IN1(\fpu_add_frac_dp/n2469 ), .IN2(n715), .Q(n4583) );
  AND3X1 U4685 ( .IN1(n4587), .IN2(n4588), .IN3(n4589), .Q(n4581) );
  XOR2X1 U4686 ( .IN1(\fpu_add_frac_dp/n940 ), .IN2(\fpu_add_frac_dp/n2474 ), 
        .Q(n4589) );
  NAND2X0 U4687 ( .IN1(\fpu_add_ctl/n116 ), .IN2(n4590), .QN(n4588) );
  NAND3X0 U4688 ( .IN1(n4591), .IN2(n4592), .IN3(n4593), .QN(n4590) );
  XOR2X1 U4689 ( .IN1(n591), .IN2(\fpu_add_frac_dp/n2521 ), .Q(n4593) );
  XOR2X1 U4690 ( .IN1(n593), .IN2(\fpu_add_frac_dp/n2534 ), .Q(n4592) );
  XOR2X1 U4691 ( .IN1(n592), .IN2(\fpu_add_frac_dp/n945 ), .Q(n4591) );
  XOR2X1 U4692 ( .IN1(\fpu_add_frac_dp/n942 ), .IN2(\fpu_add_frac_dp/n2473 ), 
        .Q(n4587) );
  XOR2X1 U4693 ( .IN1(\fpu_add_frac_dp/n937 ), .IN2(\fpu_add_frac_dp/n2468 ), 
        .Q(n4580) );
  XOR2X1 U4694 ( .IN1(\fpu_add_frac_dp/n943 ), .IN2(\fpu_add_frac_dp/n2446 ), 
        .Q(n4579) );
  OAI22X1 U4695 ( .IN1(n4057), .IN2(n2050), .IN3(n4114), .IN4(
        \fpu_add_ctl/n38 ), .QN(\fpu_add_ctl/n578 ) );
  OA22X1 U4696 ( .IN1(n2685), .IN2(n2687), .IN3(n2686), .IN4(n4594), .Q(n2050)
         );
  AND2X1 U4697 ( .IN1(n2687), .IN2(n2685), .Q(n4594) );
  NAND2X0 U4698 ( .IN1(n928), .IN2(n105), .QN(n2686) );
  NOR2X0 U4699 ( .IN1(\fpu_add_exp_dp/n245 ), .IN2(\fpu_add_exp_dp/n174 ), 
        .QN(n2687) );
  AOI22X1 U4700 ( .IN1(n2680), .IN2(n2681), .IN3(n2679), .IN4(n4595), .QN(
        n2685) );
  OR2X1 U4701 ( .IN1(n2681), .IN2(n2680), .Q(n4595) );
  OA21X1 U4702 ( .IN1(\fpu_add_exp_dp/n246 ), .IN2(\fpu_add_exp_dp/n175 ), 
        .IN3(\fpu_add_exp_dp/n170 ), .Q(n2679) );
  AO22X1 U4703 ( .IN1(n2682), .IN2(n2684), .IN3(n2683), .IN4(n4596), .Q(n2681)
         );
  OR2X1 U4704 ( .IN1(n2684), .IN2(n2682), .Q(n4596) );
  OA21X1 U4705 ( .IN1(\fpu_add_exp_dp/n247 ), .IN2(\fpu_add_exp_dp/n176 ), 
        .IN3(\fpu_add_exp_dp/n171 ), .Q(n2683) );
  AO22X1 U4706 ( .IN1(n2688), .IN2(n2690), .IN3(n4597), .IN4(n2689), .Q(n2684)
         );
  AO22X1 U4707 ( .IN1(n936), .IN2(n105), .IN3(n545), .IN4(n41), .Q(n2689) );
  OR2X1 U4708 ( .IN1(n2690), .IN2(n2688), .Q(n4597) );
  AO22X1 U4709 ( .IN1(n2692), .IN2(n2693), .IN3(n2691), .IN4(n4598), .Q(n2690)
         );
  OR2X1 U4710 ( .IN1(n2693), .IN2(n2692), .Q(n4598) );
  OA22X1 U4711 ( .IN1(\fpu_add_exp_dp/n249 ), .IN2(\fpu_add_exp_dp/n178 ), 
        .IN3(\fpu_add_exp_dp/n246 ), .IN4(\fpu_add_exp_dp/n197 ), .Q(n2691) );
  AO22X1 U4712 ( .IN1(n2720), .IN2(n2722), .IN3(n2721), .IN4(n4599), .Q(n2693)
         );
  OR2X1 U4713 ( .IN1(n2722), .IN2(n2720), .Q(n4599) );
  OA22X1 U4714 ( .IN1(\fpu_add_exp_dp/n250 ), .IN2(\fpu_add_exp_dp/n179 ), 
        .IN3(\fpu_add_exp_dp/n247 ), .IN4(\fpu_add_exp_dp/n198 ), .Q(n2721) );
  AO22X1 U4715 ( .IN1(n2659), .IN2(n2661), .IN3(n2660), .IN4(n4600), .Q(n2722)
         );
  OR2X1 U4716 ( .IN1(n2661), .IN2(n2659), .Q(n4600) );
  OA22X1 U4717 ( .IN1(\fpu_add_exp_dp/n251 ), .IN2(\fpu_add_exp_dp/n180 ), 
        .IN3(\fpu_add_exp_dp/n248 ), .IN4(\fpu_add_exp_dp/n199 ), .Q(n2660) );
  AO22X1 U4718 ( .IN1(n2645), .IN2(n2647), .IN3(n2646), .IN4(n4601), .Q(n2661)
         );
  OR2X1 U4719 ( .IN1(n2647), .IN2(n2645), .Q(n4601) );
  OA22X1 U4720 ( .IN1(\fpu_add_exp_dp/n252 ), .IN2(\fpu_add_exp_dp/n181 ), 
        .IN3(\fpu_add_exp_dp/n249 ), .IN4(\fpu_add_exp_dp/n200 ), .Q(n2646) );
  AO22X1 U4721 ( .IN1(n4602), .IN2(n2635), .IN3(n2634), .IN4(n4603), .Q(n2647)
         );
  NAND2X0 U4722 ( .IN1(n4604), .IN2(n2633), .QN(n4603) );
  OA22X1 U4723 ( .IN1(\fpu_add_exp_dp/n253 ), .IN2(\fpu_add_exp_dp/n182 ), 
        .IN3(\fpu_add_exp_dp/n250 ), .IN4(\fpu_add_exp_dp/n201 ), .Q(n2634) );
  INVX0 U4724 ( .INP(n4604), .ZN(n2635) );
  OA22X1 U4725 ( .IN1(n2052), .IN2(n2621), .IN3(n2620), .IN4(n4605), .Q(n4604)
         );
  AND2X1 U4726 ( .IN1(n2621), .IN2(n2052), .Q(n4605) );
  AO22X1 U4727 ( .IN1(n1066), .IN2(n558), .IN3(n152), .IN4(n61), .Q(n2620) );
  OA22X1 U4728 ( .IN1(\fpu_add_exp_dp/n232 ), .IN2(\fpu_add_exp_dp/n194 ), 
        .IN3(\fpu_add_exp_dp/n229 ), .IN4(\fpu_add_exp_dp/n210 ), .Q(n2621) );
  OR2X1 U4729 ( .IN1(n2612), .IN2(n2611), .Q(n2052) );
  OA22X1 U4730 ( .IN1(\fpu_add_exp_dp/n233 ), .IN2(\fpu_add_exp_dp/n195 ), 
        .IN3(\fpu_add_exp_dp/n230 ), .IN4(\fpu_add_exp_dp/n211 ), .Q(n2611) );
  AO221X1 U4731 ( .IN1(n151), .IN2(n1033), .IN3(n510), .IN4(n60), .IN5(n13), 
        .Q(n2612) );
  INVX0 U4732 ( .INP(n2633), .ZN(n4602) );
  OA22X1 U4733 ( .IN1(\fpu_add_exp_dp/n209 ), .IN2(\fpu_add_exp_dp/n228 ), 
        .IN3(\fpu_add_exp_dp/n193 ), .IN4(\fpu_add_exp_dp/n231 ), .Q(n2633) );
  AO22X1 U4734 ( .IN1(n958), .IN2(n42), .IN3(n514), .IN4(n109), .Q(n2645) );
  AO22X1 U4735 ( .IN1(n959), .IN2(n41), .IN3(n515), .IN4(n110), .Q(n2659) );
  AO22X1 U4736 ( .IN1(n960), .IN2(n126), .IN3(n516), .IN4(n49), .Q(n2720) );
  AO22X1 U4737 ( .IN1(n937), .IN2(n127), .IN3(n546), .IN4(n42), .Q(n2692) );
  OA221X1 U4738 ( .IN1(\fpu_add_exp_dp/n248 ), .IN2(\fpu_add_exp_dp/n177 ), 
        .IN3(\fpu_add_exp_dp/n245 ), .IN4(\fpu_add_exp_dp/n196 ), .IN5(
        \fpu_add_exp_dp/n172 ), .Q(n2688) );
  NOR2X0 U4739 ( .IN1(\fpu_add_exp_dp/n187 ), .IN2(\fpu_add_exp_dp/n225 ), 
        .QN(n2682) );
  NOR2X0 U4740 ( .IN1(\fpu_add_exp_dp/n186 ), .IN2(\fpu_add_exp_dp/n224 ), 
        .QN(n2680) );
  AO22X1 U4741 ( .IN1(n1472), .IN2(n851), .IN3(n1340), .IN4(n1741), .Q(
        \fpu_add_ctl/n577 ) );
  OAI22X1 U4742 ( .IN1(n4057), .IN2(n1752), .IN3(n4114), .IN4(
        \fpu_add_ctl/n338 ), .QN(\fpu_add_ctl/n576 ) );
  AO22X1 U4743 ( .IN1(n1338), .IN2(n1751), .IN3(n1470), .IN4(n1173), .Q(
        \fpu_add_ctl/n575 ) );
  AO22X1 U4744 ( .IN1(n1340), .IN2(n1749), .IN3(n1471), .IN4(n1213), .Q(
        \fpu_add_ctl/n574 ) );
  AND2X1 U4745 ( .IN1(n4606), .IN2(n338), .Q(n1749) );
  AO22X1 U4746 ( .IN1(n102), .IN2(n847), .IN3(n460), .IN4(n44), .Q(n4606) );
  AO22X1 U4747 ( .IN1(n4607), .IN2(n1339), .IN3(n1471), .IN4(n422), .Q(
        \fpu_add_ctl/n573 ) );
  AO22X1 U4748 ( .IN1(n4000), .IN2(n1068), .IN3(n4608), .IN4(n1340), .Q(
        \fpu_add_ctl/n572 ) );
  NOR2X0 U4749 ( .IN1(n4609), .IN2(n598), .QN(n4608) );
  OA22X1 U4750 ( .IN1(\fpu_add_ctl/n203 ), .IN2(\fpu_add_ctl/n127 ), .IN3(
        \fpu_add_ctl/n332 ), .IN4(\fpu_add_ctl/n205 ), .Q(n4609) );
  AO21X1 U4751 ( .IN1(n1467), .IN2(n1217), .IN3(n4610), .Q(\fpu_add_ctl/n571 )
         );
  NOR4X0 U4752 ( .IN1(n4611), .IN2(n4612), .IN3(\fpu_add_ctl/n122 ), .IN4(
        \fpu_add_ctl/n117 ), .QN(n4610) );
  OA21X1 U4753 ( .IN1(n4613), .IN2(n4614), .IN3(\fpu_add_ctl/n202 ), .Q(n4612)
         );
  OR3X1 U4754 ( .IN1(n4615), .IN2(n4616), .IN3(n4057), .Q(n4611) );
  AO22X1 U4755 ( .IN1(n1337), .IN2(n1657), .IN3(n1471), .IN4(n957), .Q(
        \fpu_add_ctl/n570 ) );
  AO22X1 U4756 ( .IN1(n4000), .IN2(n149), .IN3(n4617), .IN4(n4618), .Q(
        \fpu_add_ctl/n569 ) );
  NAND4X0 U4757 ( .IN1(n4619), .IN2(n640), .IN3(n4620), .IN4(n4621), .QN(n4618) );
  OA22X1 U4758 ( .IN1(\fpu_add_ctl/n316 ), .IN2(n4622), .IN3(\fpu_add_ctl/n41 ), .IN4(n4623), .Q(n4621) );
  AOI22X1 U4759 ( .IN1(n422), .IN2(\fpu_add_ctl/n310 ), .IN3(n1068), .IN4(
        \fpu_add_ctl/n338 ), .QN(n4623) );
  OA21X1 U4760 ( .IN1(\fpu_add_ctl/n34 ), .IN2(n422), .IN3(\fpu_add_ctl/n310 ), 
        .Q(n4622) );
  NAND4X0 U4761 ( .IN1(n4624), .IN2(\fpu_add_ctl/n37 ), .IN3(\fpu_add_ctl/n31 ), .IN4(n4625), .QN(n4620) );
  NOR3X0 U4762 ( .IN1(n4626), .IN2(\fpu_add_ctl/n200 ), .IN3(
        \fpu_add_ctl/n196 ), .QN(n4625) );
  NOR2X0 U4763 ( .IN1(n4627), .IN2(n433), .QN(n4626) );
  NAND4X0 U4764 ( .IN1(\fpu_add_ctl/n37 ), .IN2(n4628), .IN3(n4629), .IN4(
        n4630), .QN(n4619) );
  AO21X1 U4765 ( .IN1(n4631), .IN2(n4632), .IN3(n4627), .Q(n4630) );
  XOR2X1 U4766 ( .IN1(\fpu_add_ctl/n139 ), .IN2(\fpu_add_ctl/n316 ), .Q(n4627)
         );
  OAI21X1 U4767 ( .IN1(n4624), .IN2(n4631), .IN3(\fpu_add_ctl/n41 ), .QN(n4629) );
  NAND2X0 U4768 ( .IN1(\fpu_add_ctl/n313 ), .IN2(n957), .QN(n4628) );
  AO21X1 U4769 ( .IN1(n1337), .IN2(n270), .IN3(n4075), .Q(n4617) );
  NOR2X0 U4770 ( .IN1(n4057), .IN2(\fpu_add_ctl/n938 ), .QN(n4075) );
  NAND3X0 U4771 ( .IN1(n4633), .IN2(n4634), .IN3(n4635), .QN(
        \fpu_add_ctl/n568 ) );
  MUX21X1 U4772 ( .IN1(n4636), .IN2(n4637), .S(\fpu_add_ctl/n316 ), .Q(n4635)
         );
  NAND2X0 U4773 ( .IN1(n4000), .IN2(n1082), .QN(n4633) );
  NAND3X0 U4774 ( .IN1(n4638), .IN2(n4634), .IN3(n4639), .QN(
        \fpu_add_ctl/n567 ) );
  MUX21X1 U4775 ( .IN1(n4637), .IN2(n4636), .S(\fpu_add_ctl/n316 ), .Q(n4639)
         );
  NAND4X0 U4776 ( .IN1(n4640), .IN2(n4631), .IN3(n4632), .IN4(n754), .QN(n4636) );
  NAND2X0 U4777 ( .IN1(n4641), .IN2(n4640), .QN(n4637) );
  MUX21X1 U4778 ( .IN1(n4642), .IN2(\fpu_add_ctl/n32 ), .S(\fpu_add_ctl/n313 ), 
        .Q(n4641) );
  NOR2X0 U4779 ( .IN1(n4624), .IN2(n4631), .QN(n4642) );
  OA21X1 U4780 ( .IN1(\fpu_add_ctl/n39 ), .IN2(\fpu_add_ctl/n335 ), .IN3(
        \fpu_add_ctl/n38 ), .Q(n4631) );
  INVX0 U4781 ( .INP(n4632), .ZN(n4624) );
  NAND2X0 U4782 ( .IN1(\fpu_add_ctl/n40 ), .IN2(n1004), .QN(n4632) );
  NAND2X0 U4783 ( .IN1(n4640), .IN2(n851), .QN(n4634) );
  NOR2X0 U4784 ( .IN1(n4057), .IN2(\fpu_add_ctl/n143 ), .QN(n4640) );
  NAND2X0 U4785 ( .IN1(n4000), .IN2(n1083), .QN(n4638) );
  AO22X1 U4786 ( .IN1(n1339), .IN2(n149), .IN3(n1471), .IN4(n884), .Q(
        \fpu_add_ctl/n566 ) );
  AO222X1 U4787 ( .IN1(n4412), .IN2(n149), .IN3(n4413), .IN4(n884), .IN5(n1461), .IN6(n444), .Q(\fpu_add_ctl/n565 ) );
  NOR2X0 U4788 ( .IN1(n455), .IN2(n4057), .QN(n4413) );
  NOR2X0 U4789 ( .IN1(n4057), .IN2(\fpu_add_ctl/n101 ), .QN(n4412) );
  AO22X1 U4790 ( .IN1(n1338), .IN2(n1082), .IN3(n1471), .IN4(n556), .Q(
        \fpu_add_ctl/n564 ) );
  AO22X1 U4791 ( .IN1(n1340), .IN2(n1083), .IN3(n1471), .IN4(n557), .Q(
        \fpu_add_ctl/n563 ) );
  AO22X1 U4792 ( .IN1(n1337), .IN2(n444), .IN3(n1471), .IN4(add_sign_out), .Q(
        \fpu_add_ctl/n562 ) );
  AO22X1 U4793 ( .IN1(n1472), .IN2(add_cc_out[0]), .IN3(n4419), .IN4(n556), 
        .Q(\fpu_add_ctl/n561 ) );
  AO22X1 U4794 ( .IN1(n4000), .IN2(add_cc_out[1]), .IN3(n4419), .IN4(n557), 
        .Q(\fpu_add_ctl/n560 ) );
  NOR2X0 U4795 ( .IN1(n4057), .IN2(\fpu_add_ctl/n86 ), .QN(n4419) );
  AO22X1 U4796 ( .IN1(n1339), .IN2(n4643), .IN3(n1471), .IN4(n903), .Q(
        \fpu_add_ctl/n559 ) );
  AO221X1 U4797 ( .IN1(n1751), .IN2(n4644), .IN3(n4607), .IN4(n4645), .IN5(
        n4646), .Q(n4643) );
  NAND2X0 U4798 ( .IN1(n4647), .IN2(n1740), .QN(n4646) );
  NAND3X0 U4799 ( .IN1(n1657), .IN2(n1737), .IN3(n1656), .QN(n1740) );
  INVX0 U4800 ( .INP(n4648), .ZN(n1656) );
  NOR4X0 U4801 ( .IN1(n4649), .IN2(n598), .IN3(\fpu_add_ctl/n317 ), .IN4(n4650), .QN(n1657) );
  OA22X1 U4802 ( .IN1(\fpu_add_ctl/n330 ), .IN2(n4613), .IN3(
        \fpu_add_ctl/n309 ), .IN4(n4616), .Q(n4650) );
  OA22X1 U4803 ( .IN1(\fpu_add_ctl/n330 ), .IN2(n4614), .IN3(
        \fpu_add_ctl/n309 ), .IN4(n4615), .Q(n4649) );
  NAND3X0 U4804 ( .IN1(n1741), .IN2(n18), .IN3(n4386), .QN(n4647) );
  INVX0 U4805 ( .INP(n1750), .ZN(n4607) );
  AO21X1 U4806 ( .IN1(n4651), .IN2(n4652), .IN3(n598), .Q(n1750) );
  NAND3X0 U4807 ( .IN1(n743), .IN2(n102), .IN3(\fpu_add_ctl/n332 ), .QN(n4652)
         );
  NAND3X0 U4808 ( .IN1(n744), .IN2(n44), .IN3(\fpu_add_ctl/n127 ), .QN(n4651)
         );
  OR3X1 U4809 ( .IN1(n4048), .IN2(a1stg_fdtos), .IN3(n4645), .Q(n4644) );
  AO21X1 U4810 ( .IN1(n4386), .IN2(\fpu_add_ctl/n318 ), .IN3(n1737), .Q(n4645)
         );
  AND4X1 U4811 ( .IN1(n4406), .IN2(n4400), .IN3(n585), .IN4(n172), .Q(n4386)
         );
  AOI21X1 U4812 ( .IN1(n4653), .IN2(n4654), .IN3(\fpu_add_ctl/n317 ), .QN(
        n1751) );
  NAND3X0 U4813 ( .IN1(n730), .IN2(n102), .IN3(\fpu_add_ctl/n333 ), .QN(n4654)
         );
  NAND3X0 U4814 ( .IN1(n731), .IN2(n44), .IN3(\fpu_add_ctl/n121 ), .QN(n4653)
         );
  AO22X1 U4815 ( .IN1(n4000), .IN2(n1077), .IN3(n1338), .IN4(n4655), .Q(
        \fpu_add_ctl/n558 ) );
  NAND2X0 U4816 ( .IN1(n1877), .IN2(n2719), .QN(n4655) );
  NAND2X0 U4817 ( .IN1(n4656), .IN2(n1867), .QN(n2719) );
  OA22X1 U4818 ( .IN1(n338), .IN2(\fpu_add_ctl/n324 ), .IN3(n915), .IN4(n129), 
        .Q(n1877) );
  AO22X1 U4819 ( .IN1(n4000), .IN2(n140), .IN3(n1337), .IN4(n4657), .Q(
        \fpu_add_ctl/n557 ) );
  AO21X1 U4820 ( .IN1(n1932), .IN2(n4658), .IN3(n903), .Q(n4657) );
  NAND4X0 U4821 ( .IN1(n4659), .IN2(n4660), .IN3(n4661), .IN4(n4662), .QN(
        n4658) );
  NOR4X0 U4822 ( .IN1(n4663), .IN2(n4087), .IN3(n4083), .IN4(n4085), .QN(n4662) );
  XOR3X1 U4823 ( .IN1(\fpu_add_exp_dp/n132 ), .IN2(\fpu_add_exp_dp/n119 ), 
        .IN3(n4664), .Q(n4085) );
  XOR3X1 U4824 ( .IN1(\fpu_add_exp_dp/n133 ), .IN2(\fpu_add_exp_dp/n120 ), 
        .IN3(n4665), .Q(n4083) );
  XOR3X1 U4825 ( .IN1(\fpu_add_exp_dp/n131 ), .IN2(\fpu_add_exp_dp/n118 ), 
        .IN3(n4666), .Q(n4087) );
  NAND4X0 U4826 ( .IN1(n4081), .IN2(n4667), .IN3(n4668), .IN4(n270), .QN(n4663) );
  OR2X1 U4827 ( .IN1(n4669), .IN2(\fpu_add_ctl/n130 ), .Q(n4668) );
  INVX0 U4828 ( .INP(n4074), .ZN(n4667) );
  XOR3X1 U4829 ( .IN1(\fpu_add_exp_dp/n135 ), .IN2(\fpu_add_exp_dp/n122 ), 
        .IN3(n128), .Q(n4074) );
  XNOR3X1 U4830 ( .IN1(\fpu_add_exp_dp/n134 ), .IN2(\fpu_add_exp_dp/n121 ), 
        .IN3(n4670), .Q(n4081) );
  NOR4X0 U4831 ( .IN1(n4091), .IN2(n4093), .IN3(n4099), .IN4(n4104), .QN(n4661) );
  XOR3X1 U4832 ( .IN1(\fpu_add_exp_dp/n127 ), .IN2(\fpu_add_exp_dp/n114 ), 
        .IN3(n4671), .Q(n4104) );
  XOR3X1 U4833 ( .IN1(\fpu_add_exp_dp/n128 ), .IN2(\fpu_add_exp_dp/n115 ), 
        .IN3(n4672), .Q(n4099) );
  XOR3X1 U4834 ( .IN1(\fpu_add_exp_dp/n129 ), .IN2(\fpu_add_exp_dp/n116 ), 
        .IN3(n4673), .Q(n4093) );
  XOR3X1 U4835 ( .IN1(\fpu_add_exp_dp/n130 ), .IN2(\fpu_add_exp_dp/n117 ), 
        .IN3(n4674), .Q(n4091) );
  NOR2X0 U4836 ( .IN1(n4107), .IN2(n4110), .QN(n4659) );
  XOR3X1 U4837 ( .IN1(\fpu_add_exp_dp/n125 ), .IN2(\fpu_add_exp_dp/n112 ), 
        .IN3(n4675), .Q(n4110) );
  XOR3X1 U4838 ( .IN1(\fpu_add_exp_dp/n126 ), .IN2(\fpu_add_exp_dp/n113 ), 
        .IN3(n4676), .Q(n4107) );
  AND2X1 U4839 ( .IN1(\fpu_add_ctl/n329 ), .IN2(n4111), .Q(n1932) );
  AO22X1 U4840 ( .IN1(n1338), .IN2(n1077), .IN3(n1471), .IN4(n137), .Q(
        \fpu_add_ctl/n556 ) );
  OAI22X1 U4841 ( .IN1(n4111), .IN2(n4057), .IN3(n4114), .IN4(
        \fpu_add_ctl/n16 ), .QN(\fpu_add_ctl/n555 ) );
  XNOR3X1 U4842 ( .IN1(\fpu_add_exp_dp/n124 ), .IN2(n629), .IN3(n3968), .Q(
        n4111) );
  INVX0 U4843 ( .INP(n3967), .ZN(n3968) );
  AO22X1 U4844 ( .IN1(n4675), .IN2(n298), .IN3(n4677), .IN4(n680), .Q(n3967)
         );
  OR2X1 U4845 ( .IN1(n298), .IN2(n4675), .Q(n4677) );
  AO22X1 U4846 ( .IN1(n4676), .IN2(n300), .IN3(n4678), .IN4(n681), .Q(n4675)
         );
  OR2X1 U4847 ( .IN1(n300), .IN2(n4676), .Q(n4678) );
  AO22X1 U4848 ( .IN1(n4671), .IN2(n301), .IN3(n4679), .IN4(n682), .Q(n4676)
         );
  OR2X1 U4849 ( .IN1(n301), .IN2(n4671), .Q(n4679) );
  AO22X1 U4850 ( .IN1(n4672), .IN2(n308), .IN3(n4680), .IN4(n683), .Q(n4671)
         );
  OR2X1 U4851 ( .IN1(n308), .IN2(n4672), .Q(n4680) );
  AO22X1 U4852 ( .IN1(n4673), .IN2(n302), .IN3(n4681), .IN4(n661), .Q(n4672)
         );
  OR2X1 U4853 ( .IN1(n302), .IN2(n4673), .Q(n4681) );
  AO22X1 U4854 ( .IN1(n4674), .IN2(n299), .IN3(n4682), .IN4(n684), .Q(n4673)
         );
  OR2X1 U4855 ( .IN1(n299), .IN2(n4674), .Q(n4682) );
  AO22X1 U4856 ( .IN1(n4666), .IN2(n303), .IN3(n4683), .IN4(n685), .Q(n4674)
         );
  OR2X1 U4857 ( .IN1(n303), .IN2(n4666), .Q(n4683) );
  AO22X1 U4858 ( .IN1(n4664), .IN2(n304), .IN3(n4684), .IN4(n686), .Q(n4666)
         );
  OR2X1 U4859 ( .IN1(n304), .IN2(n4664), .Q(n4684) );
  AO22X1 U4860 ( .IN1(n4665), .IN2(n305), .IN3(n4685), .IN4(n687), .Q(n4664)
         );
  OR2X1 U4861 ( .IN1(n305), .IN2(n4665), .Q(n4685) );
  AO22X1 U4862 ( .IN1(n4670), .IN2(n297), .IN3(n4686), .IN4(n676), .Q(n4665)
         );
  OR2X1 U4863 ( .IN1(n297), .IN2(n4670), .Q(n4686) );
  AO22X1 U4864 ( .IN1(n128), .IN2(n830), .IN3(n4687), .IN4(n315), .Q(n4670) );
  NAND2X0 U4865 ( .IN1(\fpu_add_exp_dp/n122 ), .IN2(\fpu_add_ctl/n129 ), .QN(
        n4687) );
  AO22X1 U4866 ( .IN1(n4000), .IN2(n1249), .IN3(n1339), .IN4(n4688), .Q(
        \fpu_add_ctl/n554 ) );
  AO22X1 U4867 ( .IN1(n3753), .IN2(n1008), .IN3(n3754), .IN4(n547), .Q(n4688)
         );
  AO22X1 U4868 ( .IN1(n4000), .IN2(n1272), .IN3(n4689), .IN4(n1339), .Q(
        \fpu_add_ctl/n553 ) );
  OA21X1 U4869 ( .IN1(n4690), .IN2(n4691), .IN3(n4692), .Q(n4689) );
  OAI22X1 U4870 ( .IN1(n3753), .IN2(\fpu_add_ctl/n110 ), .IN3(n3754), .IN4(
        \fpu_add_ctl/n109 ), .QN(n4692) );
  OR4X1 U4871 ( .IN1(n3753), .IN2(n221), .IN3(n35), .IN4(n88), .Q(n3754) );
  NAND2X0 U4872 ( .IN1(\fpu_add_exp_dp/n136 ), .IN2(\fpu_add_exp_dp/n137 ), 
        .QN(n3753) );
  NAND4X0 U4873 ( .IN1(n4669), .IN2(n4660), .IN3(\fpu_add_frac_dp/n2498 ), 
        .IN4(n1924), .QN(n4691) );
  NOR2X0 U4874 ( .IN1(n646), .IN2(n290), .QN(n1924) );
  INVX0 U4875 ( .INP(n4693), .ZN(n4660) );
  NAND4X0 U4876 ( .IN1(\fpu_add_exp_dp/n143 ), .IN2(\fpu_add_exp_dp/n145 ), 
        .IN3(\fpu_add_exp_dp/n146 ), .IN4(n1929), .QN(n4690) );
  AO22X1 U4877 ( .IN1(n4000), .IN2(n1265), .IN3(n4694), .IN4(n4695), .Q(
        \fpu_add_ctl/n552 ) );
  NOR4X0 U4878 ( .IN1(n4696), .IN2(n4669), .IN3(\fpu_add_ctl/n316 ), .IN4(
        \fpu_add_ctl/n133 ), .QN(n4695) );
  NOR4X0 U4879 ( .IN1(n4697), .IN2(n4698), .IN3(n4699), .IN4(n4700), .QN(n4669) );
  NAND4X0 U4880 ( .IN1(\fpu_add_frac_dp/n2434 ), .IN2(\fpu_add_frac_dp/n2433 ), 
        .IN3(n4701), .IN4(\fpu_add_frac_dp/n2297 ), .QN(n4700) );
  NOR2X0 U4881 ( .IN1(n722), .IN2(n423), .QN(n4701) );
  NAND4X0 U4882 ( .IN1(\fpu_add_frac_dp/n2277 ), .IN2(n904), .IN3(
        \fpu_add_frac_dp/n2304 ), .IN4(n4702), .QN(n4699) );
  AND3X1 U4883 ( .IN1(\fpu_add_frac_dp/n2432 ), .IN2(\fpu_add_frac_dp/n2362 ), 
        .IN3(\fpu_add_frac_dp/n2359 ), .Q(n4702) );
  NAND4X0 U4884 ( .IN1(\fpu_add_frac_dp/n2510 ), .IN2(\fpu_add_frac_dp/n2503 ), 
        .IN3(n4703), .IN4(\fpu_add_frac_dp/n2499 ), .QN(n4698) );
  NOR2X0 U4885 ( .IN1(n723), .IN2(n424), .QN(n4703) );
  NAND4X0 U4886 ( .IN1(\fpu_add_frac_dp/n2299 ), .IN2(\fpu_add_frac_dp/n2420 ), 
        .IN3(n4704), .IN4(\fpu_add_frac_dp/n2273 ), .QN(n4697) );
  NOR2X0 U4887 ( .IN1(n724), .IN2(n426), .QN(n4704) );
  NAND3X0 U4888 ( .IN1(n648), .IN2(n73), .IN3(n289), .QN(n4696) );
  NOR4X0 U4889 ( .IN1(n4705), .IN2(n4693), .IN3(n725), .IN4(n4057), .QN(n4694)
         );
  NAND4X0 U4890 ( .IN1(n4706), .IN2(n4707), .IN3(n4708), .IN4(n4709), .QN(
        n4693) );
  NOR4X0 U4891 ( .IN1(n4710), .IN2(n4711), .IN3(n4712), .IN4(n4713), .QN(n4709) );
  NAND4X0 U4892 ( .IN1(\fpu_add_frac_dp/n2276 ), .IN2(\fpu_add_frac_dp/n2302 ), 
        .IN3(\fpu_add_frac_dp/n2422 ), .IN4(\fpu_add_frac_dp/n2355 ), .QN(
        n4713) );
  NAND4X0 U4893 ( .IN1(\fpu_add_frac_dp/n2275 ), .IN2(\fpu_add_frac_dp/n2301 ), 
        .IN3(\fpu_add_frac_dp/n2421 ), .IN4(\fpu_add_frac_dp/n2511 ), .QN(
        n4712) );
  NAND4X0 U4894 ( .IN1(\fpu_add_frac_dp/n2435 ), .IN2(\fpu_add_frac_dp/n2354 ), 
        .IN3(\fpu_add_frac_dp/n2274 ), .IN4(\fpu_add_frac_dp/n2300 ), .QN(
        n4711) );
  NAND4X0 U4895 ( .IN1(n1009), .IN2(n561), .IN3(n153), .IN4(n62), .QN(n4710)
         );
  NOR4X0 U4896 ( .IN1(n4714), .IN2(n142), .IN3(n343), .IN4(n706), .QN(n4708)
         );
  NAND4X0 U4897 ( .IN1(\fpu_add_frac_dp/n2431 ), .IN2(\fpu_add_frac_dp/n2418 ), 
        .IN3(\fpu_add_frac_dp/n2351 ), .IN4(\fpu_add_frac_dp/n2505 ), .QN(
        n4714) );
  NOR4X0 U4898 ( .IN1(n58), .IN2(n143), .IN3(n344), .IN4(n707), .QN(n4707) );
  NOR4X0 U4899 ( .IN1(n59), .IN2(n144), .IN3(n345), .IN4(n708), .QN(n4706) );
  NAND3X0 U4900 ( .IN1(n1901), .IN2(n1929), .IN3(n1920), .QN(n4705) );
  NOR2X0 U4901 ( .IN1(n646), .IN2(\fpu_add_exp_dp/n144 ), .QN(n1920) );
  NOR4X0 U4902 ( .IN1(n711), .IN2(n221), .IN3(n35), .IN4(n88), .QN(n1929) );
  NOR2X0 U4903 ( .IN1(\fpu_add_exp_dp/n147 ), .IN2(\fpu_add_exp_dp/n145 ), 
        .QN(n1901) );
  AO22X1 U4904 ( .IN1(n1340), .IN2(n140), .IN3(n1471), .IN4(n512), .Q(
        \fpu_add_ctl/n551 ) );
  AO222X1 U4905 ( .IN1(n1472), .IN2(n1074), .IN3(n4715), .IN4(n140), .IN5(
        n4716), .IN6(n512), .Q(\fpu_add_ctl/n550 ) );
  AO22X1 U4906 ( .IN1(n1337), .IN2(n137), .IN3(n1471), .IN4(n905), .Q(
        \fpu_add_ctl/n549 ) );
  AO222X1 U4907 ( .IN1(n1472), .IN2(n452), .IN3(n4715), .IN4(n137), .IN5(n4716), .IN6(n905), .Q(\fpu_add_ctl/n548 ) );
  AO22X1 U4908 ( .IN1(n1339), .IN2(n4717), .IN3(n1471), .IN4(n513), .Q(
        \fpu_add_ctl/n547 ) );
  AO222X1 U4909 ( .IN1(n1472), .IN2(n1245), .IN3(n4715), .IN4(n4717), .IN5(
        n4716), .IN6(n513), .Q(\fpu_add_ctl/n546 ) );
  AOI21X1 U4910 ( .IN1(\fpu_add_ctl/n102 ), .IN2(\fpu_add_ctl/n325 ), .IN3(
        n4057), .QN(n4716) );
  OAI21X1 U4911 ( .IN1(\fpu_add_ctl/n16 ), .IN2(n4718), .IN3(\fpu_add_ctl/n13 ), .QN(n4717) );
  OA21X1 U4912 ( .IN1(\fpu_add_ctl/n15 ), .IN2(n4719), .IN3(\fpu_add_ctl/n14 ), 
        .Q(n4718) );
  OA21X1 U4913 ( .IN1(\fpu_add_frac_dp/n510 ), .IN2(\fpu_add_ctl/n97 ), .IN3(
        \fpu_add_frac_dp/n515 ), .Q(n4719) );
  AND3X1 U4914 ( .IN1(\fpu_add_ctl/n325 ), .IN2(n1340), .IN3(
        \fpu_add_ctl/n102 ), .Q(n4715) );
  AO22X1 U4915 ( .IN1(n1338), .IN2(n1074), .IN3(n1472), .IN4(add_exc_out[4]), 
        .Q(\fpu_add_ctl/n545 ) );
  AO21X1 U4916 ( .IN1(n1468), .IN2(n1234), .IN3(n4720), .Q(\fpu_add_ctl/n544 )
         );
  NOR4X0 U4917 ( .IN1(n4721), .IN2(n4722), .IN3(n4723), .IN4(n4057), .QN(n4720) );
  OA22X1 U4918 ( .IN1(\fpu_add_frac_dp/n582 ), .IN2(n4724), .IN3(
        \fpu_add_ctl/n941 ), .IN4(\fpu_add_ctl/n89 ), .Q(n4722) );
  INVX0 U4919 ( .INP(n4182), .ZN(n4721) );
  AO22X1 U4920 ( .IN1(n4210), .IN2(n21), .IN3(n4725), .IN4(n4211), .Q(n4182)
         );
  AO21X1 U4921 ( .IN1(n4726), .IN2(n4727), .IN3(n4728), .Q(n4211) );
  NOR4X0 U4922 ( .IN1(\fpu_add_ctl/n307 ), .IN2(n2880), .IN3(n4729), .IN4(n291), .QN(n4728) );
  NOR2X0 U4923 ( .IN1(n2984), .IN2(n4730), .QN(n4729) );
  INVX0 U4924 ( .INP(n2983), .ZN(n2880) );
  AO21X1 U4925 ( .IN1(n55), .IN2(n452), .IN3(n148), .Q(n4725) );
  AO22X1 U4926 ( .IN1(n4726), .IN2(n4731), .IN3(n4732), .IN4(n2973), .Q(n4210)
         );
  NAND2X0 U4927 ( .IN1(n4733), .IN2(n4734), .QN(n4732) );
  NAND3X0 U4928 ( .IN1(n4735), .IN2(n1084), .IN3(\fpu_add_ctl/n937 ), .QN(
        n4734) );
  INVX0 U4929 ( .INP(n4733), .ZN(n4726) );
  NAND2X0 U4930 ( .IN1(n4736), .IN2(n291), .QN(n4733) );
  XOR2X1 U4931 ( .IN1(\fpu_add_ctl/n337 ), .IN2(\fpu_add_ctl/n307 ), .Q(n4736)
         );
  OAI22X1 U4932 ( .IN1(n4057), .IN2(n2959), .IN3(n4114), .IN4(\fpu_add_ctl/n4 ), .QN(\fpu_add_ctl/n543 ) );
  OA21X1 U4933 ( .IN1(\fpu_add_ctl/n9 ), .IN2(n4737), .IN3(n4738), .Q(n2959)
         );
  OR3X1 U4934 ( .IN1(n4213), .IN2(n4724), .IN3(n4723), .Q(n4738) );
  NAND4X0 U4935 ( .IN1(n4214), .IN2(n4136), .IN3(n4739), .IN4(n4740), .QN(
        n4723) );
  NOR4X0 U4936 ( .IN1(\fpu_add_ctl/n9 ), .IN2(n4154), .IN3(n4160), .IN4(n4148), 
        .QN(n4740) );
  INVX0 U4937 ( .INP(n4194), .ZN(n4148) );
  INVX0 U4938 ( .INP(n4219), .ZN(n4154) );
  NOR2X0 U4939 ( .IN1(n4166), .IN2(n4142), .QN(n4739) );
  INVX0 U4940 ( .INP(n4218), .ZN(n4142) );
  AND2X1 U4941 ( .IN1(\fpu_add_ctl/n941 ), .IN2(n4741), .Q(n4724) );
  NAND4X0 U4942 ( .IN1(n4215), .IN2(n4172), .IN3(n4212), .IN4(n21), .QN(n4741)
         );
  INVX0 U4943 ( .INP(n4184), .ZN(n4213) );
  OA22X1 U4944 ( .IN1(n4742), .IN2(n4743), .IN3(\fpu_add_ctl/n941 ), .IN4(
        n4744), .Q(n4737) );
  NOR2X0 U4945 ( .IN1(n21), .IN2(n420), .QN(n4743) );
  INVX0 U4946 ( .INP(n4264), .ZN(n4742) );
  NAND4X0 U4947 ( .IN1(\fpu_add_exp_dp/n98 ), .IN2(\fpu_add_exp_dp/n85 ), 
        .IN3(\fpu_add_exp_dp/n61 ), .IN4(\fpu_add_exp_dp/n60 ), .QN(n4264) );
  OAI22X1 U4948 ( .IN1(\fpu_add_ctl/n3 ), .IN2(n4114), .IN3(n4745), .IN4(n4057), .QN(\fpu_add_ctl/n542 ) );
  OA21X1 U4949 ( .IN1(n4746), .IN2(n4747), .IN3(n4748), .Q(n4745) );
  NAND4X0 U4950 ( .IN1(\fpu_add_frac_dp/n596 ), .IN2(\fpu_add_ctl/n89 ), .IN3(
        n2960), .IN4(n4749), .QN(n4748) );
  NAND4X0 U4951 ( .IN1(n4750), .IN2(n4751), .IN3(n4752), .IN4(n4753), .QN(
        n4749) );
  NOR4X0 U4952 ( .IN1(n4754), .IN2(n4755), .IN3(n4756), .IN4(n4757), .QN(n4753) );
  NAND4X0 U4953 ( .IN1(\fpu_add_frac_dp/n210 ), .IN2(\fpu_add_frac_dp/n208 ), 
        .IN3(\fpu_add_frac_dp/n206 ), .IN4(\fpu_add_frac_dp/n204 ), .QN(n4757)
         );
  NAND4X0 U4954 ( .IN1(\fpu_add_frac_dp/n202 ), .IN2(\fpu_add_frac_dp/n200 ), 
        .IN3(\fpu_add_frac_dp/n198 ), .IN4(\fpu_add_frac_dp/n196 ), .QN(n4756)
         );
  NAND4X0 U4955 ( .IN1(\fpu_add_frac_dp/n194 ), .IN2(\fpu_add_frac_dp/n192 ), 
        .IN3(\fpu_add_frac_dp/n190 ), .IN4(\fpu_add_frac_dp/n188 ), .QN(n4755)
         );
  NAND4X0 U4956 ( .IN1(\fpu_add_frac_dp/n2358 ), .IN2(\fpu_add_frac_dp/n2291 ), 
        .IN3(\fpu_add_frac_dp/n2360 ), .IN4(\fpu_add_frac_dp/n2292 ), .QN(
        n4754) );
  NOR4X0 U4957 ( .IN1(n4758), .IN2(n4759), .IN3(n4760), .IN4(n4761), .QN(n4752) );
  NAND4X0 U4958 ( .IN1(\fpu_add_frac_dp/n2347 ), .IN2(\fpu_add_frac_dp/n2346 ), 
        .IN3(\fpu_add_frac_dp/n234 ), .IN4(\fpu_add_frac_dp/n232 ), .QN(n4761)
         );
  NAND4X0 U4959 ( .IN1(\fpu_add_frac_dp/n230 ), .IN2(\fpu_add_frac_dp/n2294 ), 
        .IN3(\fpu_add_frac_dp/n2293 ), .IN4(\fpu_add_frac_dp/n228 ), .QN(n4760) );
  NAND4X0 U4960 ( .IN1(\fpu_add_frac_dp/n226 ), .IN2(\fpu_add_frac_dp/n224 ), 
        .IN3(\fpu_add_frac_dp/n222 ), .IN4(\fpu_add_frac_dp/n220 ), .QN(n4759)
         );
  NAND4X0 U4961 ( .IN1(\fpu_add_frac_dp/n218 ), .IN2(\fpu_add_frac_dp/n216 ), 
        .IN3(\fpu_add_frac_dp/n214 ), .IN4(\fpu_add_frac_dp/n212 ), .QN(n4758)
         );
  NOR4X0 U4962 ( .IN1(n4762), .IN2(n4763), .IN3(n4764), .IN4(n4765), .QN(n4751) );
  NAND4X0 U4963 ( .IN1(\fpu_add_frac_dp/n250 ), .IN2(\fpu_add_frac_dp/n248 ), 
        .IN3(\fpu_add_frac_dp/n246 ), .IN4(\fpu_add_frac_dp/n244 ), .QN(n4765)
         );
  NAND4X0 U4964 ( .IN1(\fpu_add_frac_dp/n242 ), .IN2(\fpu_add_frac_dp/n2417 ), 
        .IN3(\fpu_add_frac_dp/n2414 ), .IN4(\fpu_add_frac_dp/n2413 ), .QN(
        n4764) );
  NAND4X0 U4965 ( .IN1(\fpu_add_frac_dp/n2412 ), .IN2(\fpu_add_frac_dp/n2410 ), 
        .IN3(\fpu_add_frac_dp/n2401 ), .IN4(\fpu_add_frac_dp/n240 ), .QN(n4763) );
  NAND4X0 U4966 ( .IN1(\fpu_add_frac_dp/n238 ), .IN2(\fpu_add_frac_dp/n236 ), 
        .IN3(\fpu_add_frac_dp/n2349 ), .IN4(\fpu_add_frac_dp/n2348 ), .QN(
        n4762) );
  NOR4X0 U4967 ( .IN1(n4766), .IN2(n4767), .IN3(n4768), .IN4(n4769), .QN(n4750) );
  NAND4X0 U4968 ( .IN1(\fpu_add_frac_dp/n282 ), .IN2(\fpu_add_frac_dp/n280 ), 
        .IN3(\fpu_add_frac_dp/n278 ), .IN4(\fpu_add_frac_dp/n276 ), .QN(n4769)
         );
  NAND4X0 U4969 ( .IN1(\fpu_add_frac_dp/n274 ), .IN2(\fpu_add_frac_dp/n272 ), 
        .IN3(\fpu_add_frac_dp/n270 ), .IN4(\fpu_add_frac_dp/n268 ), .QN(n4768)
         );
  NAND4X0 U4970 ( .IN1(\fpu_add_frac_dp/n266 ), .IN2(\fpu_add_frac_dp/n264 ), 
        .IN3(\fpu_add_frac_dp/n262 ), .IN4(\fpu_add_frac_dp/n260 ), .QN(n4767)
         );
  NAND4X0 U4971 ( .IN1(\fpu_add_frac_dp/n258 ), .IN2(\fpu_add_frac_dp/n256 ), 
        .IN3(\fpu_add_frac_dp/n254 ), .IN4(\fpu_add_frac_dp/n252 ), .QN(n4766)
         );
  NOR2X0 U4972 ( .IN1(n296), .IN2(\fpu_add_ctl/n939 ), .QN(n2960) );
  NAND4X0 U4973 ( .IN1(n4166), .IN2(n4160), .IN3(n4744), .IN4(n4770), .QN(
        n4747) );
  NOR3X0 U4974 ( .IN1(n4219), .IN2(n4218), .IN3(n4194), .QN(n4770) );
  NAND4X0 U4975 ( .IN1(\fpu_add_exp_dp/n92 ), .IN2(\fpu_add_exp_dp/n75 ), 
        .IN3(\fpu_add_exp_dp/n74 ), .IN4(\fpu_add_exp_dp/n105 ), .QN(n4194) );
  NAND4X0 U4976 ( .IN1(\fpu_add_exp_dp/n93 ), .IN2(\fpu_add_exp_dp/n77 ), 
        .IN3(\fpu_add_exp_dp/n76 ), .IN4(\fpu_add_exp_dp/n106 ), .QN(n4218) );
  NAND4X0 U4977 ( .IN1(\fpu_add_exp_dp/n91 ), .IN2(\fpu_add_exp_dp/n73 ), 
        .IN3(\fpu_add_exp_dp/n72 ), .IN4(\fpu_add_exp_dp/n104 ), .QN(n4219) );
  NOR3X0 U4978 ( .IN1(n4172), .IN2(n4215), .IN3(n4212), .QN(n4744) );
  NAND4X0 U4979 ( .IN1(\fpu_add_exp_dp/n87 ), .IN2(\fpu_add_exp_dp/n65 ), 
        .IN3(\fpu_add_exp_dp/n64 ), .IN4(\fpu_add_exp_dp/n100 ), .QN(n4212) );
  NAND4X0 U4980 ( .IN1(\fpu_add_exp_dp/n99 ), .IN2(\fpu_add_exp_dp/n86 ), 
        .IN3(\fpu_add_exp_dp/n63 ), .IN4(\fpu_add_exp_dp/n62 ), .QN(n4215) );
  NAND4X0 U4981 ( .IN1(\fpu_add_exp_dp/n88 ), .IN2(\fpu_add_exp_dp/n67 ), 
        .IN3(\fpu_add_exp_dp/n66 ), .IN4(\fpu_add_exp_dp/n101 ), .QN(n4172) );
  INVX0 U4982 ( .INP(n4199), .ZN(n4160) );
  NAND4X0 U4983 ( .IN1(\fpu_add_exp_dp/n90 ), .IN2(\fpu_add_exp_dp/n71 ), 
        .IN3(\fpu_add_exp_dp/n70 ), .IN4(\fpu_add_exp_dp/n103 ), .QN(n4199) );
  INVX0 U4984 ( .INP(n4220), .ZN(n4166) );
  NAND4X0 U4985 ( .IN1(\fpu_add_exp_dp/n89 ), .IN2(\fpu_add_exp_dp/n69 ), 
        .IN3(\fpu_add_exp_dp/n68 ), .IN4(\fpu_add_exp_dp/n102 ), .QN(n4220) );
  NAND4X0 U4986 ( .IN1(n4771), .IN2(n490), .IN3(n4772), .IN4(n4773), .QN(n4746) );
  NOR3X0 U4987 ( .IN1(n4136), .IN2(n4184), .IN3(n4214), .QN(n4773) );
  NAND4X0 U4988 ( .IN1(\fpu_add_exp_dp/n95 ), .IN2(\fpu_add_exp_dp/n81 ), 
        .IN3(\fpu_add_exp_dp/n80 ), .IN4(\fpu_add_exp_dp/n108 ), .QN(n4214) );
  NAND4X0 U4989 ( .IN1(\fpu_add_exp_dp/n96 ), .IN2(\fpu_add_exp_dp/n83 ), 
        .IN3(\fpu_add_exp_dp/n82 ), .IN4(\fpu_add_exp_dp/n109 ), .QN(n4184) );
  NAND4X0 U4990 ( .IN1(\fpu_add_exp_dp/n94 ), .IN2(\fpu_add_exp_dp/n79 ), 
        .IN3(\fpu_add_exp_dp/n78 ), .IN4(\fpu_add_exp_dp/n107 ), .QN(n4136) );
  NAND2X0 U4991 ( .IN1(\fpu_add_ctl/n89 ), .IN2(\fpu_add_frac_dp/n582 ), .QN(
        n4772) );
  NAND4X0 U4992 ( .IN1(n4774), .IN2(n4775), .IN3(n4776), .IN4(n4777), .QN(
        n4771) );
  NOR4X0 U4993 ( .IN1(n4778), .IN2(n2904), .IN3(n2898), .IN4(n2902), .QN(n4777) );
  NAND3X0 U4994 ( .IN1(\fpu_add_frac_dp/n333 ), .IN2(\fpu_add_frac_dp/n223 ), 
        .IN3(\fpu_add_frac_dp/n414 ), .QN(n2902) );
  NAND3X0 U4995 ( .IN1(\fpu_add_frac_dp/n334 ), .IN2(\fpu_add_frac_dp/n225 ), 
        .IN3(\fpu_add_frac_dp/n416 ), .QN(n2898) );
  NAND3X0 U4996 ( .IN1(\fpu_add_frac_dp/n332 ), .IN2(\fpu_add_frac_dp/n221 ), 
        .IN3(\fpu_add_frac_dp/n412 ), .QN(n2904) );
  OR4X1 U4997 ( .IN1(n2896), .IN2(n2891), .IN3(n2888), .IN4(n2984), .Q(n4778)
         );
  NAND3X0 U4998 ( .IN1(\fpu_add_frac_dp/n338 ), .IN2(\fpu_add_frac_dp/n233 ), 
        .IN3(\fpu_add_frac_dp/n424 ), .QN(n2984) );
  NAND3X0 U4999 ( .IN1(\fpu_add_frac_dp/n337 ), .IN2(\fpu_add_frac_dp/n231 ), 
        .IN3(\fpu_add_frac_dp/n422 ), .QN(n2888) );
  NAND3X0 U5000 ( .IN1(\fpu_add_frac_dp/n336 ), .IN2(\fpu_add_frac_dp/n229 ), 
        .IN3(\fpu_add_frac_dp/n420 ), .QN(n2891) );
  NAND3X0 U5001 ( .IN1(\fpu_add_frac_dp/n335 ), .IN2(\fpu_add_frac_dp/n227 ), 
        .IN3(\fpu_add_frac_dp/n418 ), .QN(n2896) );
  NOR4X0 U5002 ( .IN1(n4779), .IN2(n2914), .IN3(n2908), .IN4(n2910), .QN(n4776) );
  NAND3X0 U5003 ( .IN1(\fpu_add_frac_dp/n330 ), .IN2(\fpu_add_frac_dp/n217 ), 
        .IN3(\fpu_add_frac_dp/n408 ), .QN(n2910) );
  NAND3X0 U5004 ( .IN1(\fpu_add_frac_dp/n331 ), .IN2(\fpu_add_frac_dp/n219 ), 
        .IN3(\fpu_add_frac_dp/n410 ), .QN(n2908) );
  NAND3X0 U5005 ( .IN1(\fpu_add_frac_dp/n329 ), .IN2(\fpu_add_frac_dp/n215 ), 
        .IN3(\fpu_add_frac_dp/n406 ), .QN(n2914) );
  OR3X1 U5006 ( .IN1(n2920), .IN2(n2916), .IN3(n2922), .Q(n4779) );
  NAND3X0 U5007 ( .IN1(\fpu_add_frac_dp/n326 ), .IN2(\fpu_add_frac_dp/n209 ), 
        .IN3(\fpu_add_frac_dp/n400 ), .QN(n2922) );
  NAND3X0 U5008 ( .IN1(\fpu_add_frac_dp/n328 ), .IN2(\fpu_add_frac_dp/n213 ), 
        .IN3(\fpu_add_frac_dp/n404 ), .QN(n2916) );
  NAND3X0 U5009 ( .IN1(\fpu_add_frac_dp/n327 ), .IN2(\fpu_add_frac_dp/n211 ), 
        .IN3(\fpu_add_frac_dp/n402 ), .QN(n2920) );
  NOR4X0 U5010 ( .IN1(n4780), .IN2(n2932), .IN3(n2926), .IN4(n2928), .QN(n4775) );
  NAND3X0 U5011 ( .IN1(\fpu_add_frac_dp/n324 ), .IN2(\fpu_add_frac_dp/n205 ), 
        .IN3(\fpu_add_frac_dp/n396 ), .QN(n2928) );
  NAND3X0 U5012 ( .IN1(\fpu_add_frac_dp/n325 ), .IN2(\fpu_add_frac_dp/n207 ), 
        .IN3(\fpu_add_frac_dp/n398 ), .QN(n2926) );
  NAND3X0 U5013 ( .IN1(\fpu_add_frac_dp/n323 ), .IN2(\fpu_add_frac_dp/n203 ), 
        .IN3(\fpu_add_frac_dp/n394 ), .QN(n2932) );
  OR3X1 U5014 ( .IN1(n2985), .IN2(n2940), .IN3(n2942), .Q(n4780) );
  NAND3X0 U5015 ( .IN1(\fpu_add_frac_dp/n320 ), .IN2(\fpu_add_frac_dp/n197 ), 
        .IN3(\fpu_add_frac_dp/n388 ), .QN(n2942) );
  NAND3X0 U5016 ( .IN1(\fpu_add_frac_dp/n322 ), .IN2(\fpu_add_frac_dp/n201 ), 
        .IN3(\fpu_add_frac_dp/n392 ), .QN(n2940) );
  NAND3X0 U5017 ( .IN1(\fpu_add_frac_dp/n321 ), .IN2(\fpu_add_frac_dp/n199 ), 
        .IN3(\fpu_add_frac_dp/n390 ), .QN(n2985) );
  NOR4X0 U5018 ( .IN1(n4781), .IN2(n2952), .IN3(n2946), .IN4(n2948), .QN(n4774) );
  NAND3X0 U5019 ( .IN1(\fpu_add_frac_dp/n318 ), .IN2(\fpu_add_frac_dp/n193 ), 
        .IN3(\fpu_add_frac_dp/n384 ), .QN(n2948) );
  NAND3X0 U5020 ( .IN1(\fpu_add_frac_dp/n319 ), .IN2(\fpu_add_frac_dp/n195 ), 
        .IN3(\fpu_add_frac_dp/n386 ), .QN(n2946) );
  NAND3X0 U5021 ( .IN1(\fpu_add_frac_dp/n317 ), .IN2(\fpu_add_frac_dp/n191 ), 
        .IN3(\fpu_add_frac_dp/n382 ), .QN(n2952) );
  NAND3X0 U5022 ( .IN1(n3174), .IN2(n2986), .IN3(n4782), .QN(n4781) );
  INVX0 U5023 ( .INP(n2956), .ZN(n2986) );
  NAND3X0 U5024 ( .IN1(\fpu_add_frac_dp/n316 ), .IN2(\fpu_add_frac_dp/n189 ), 
        .IN3(\fpu_add_frac_dp/n380 ), .QN(n2956) );
  INVX0 U5025 ( .INP(n2987), .ZN(n3174) );
  NAND3X0 U5026 ( .IN1(\fpu_add_frac_dp/n315 ), .IN2(\fpu_add_frac_dp/n187 ), 
        .IN3(\fpu_add_frac_dp/n378 ), .QN(n2987) );
  OAI22X1 U5027 ( .IN1(\fpu_add_ctl/n2 ), .IN2(n4114), .IN3(n4783), .IN4(n4057), .QN(\fpu_add_ctl/n541 ) );
  OA21X1 U5028 ( .IN1(\fpu_add_ctl/n9 ), .IN2(n4784), .IN3(\fpu_add_ctl/n7 ), 
        .Q(n4783) );
  OA21X1 U5029 ( .IN1(n4785), .IN2(n4786), .IN3(n4787), .Q(n4784) );
  NAND3X0 U5030 ( .IN1(n4727), .IN2(n2884), .IN3(n4788), .QN(n4787) );
  NAND2X0 U5031 ( .IN1(\fpu_add_frac_dp/n582 ), .IN2(n148), .QN(n4788) );
  NAND2X0 U5032 ( .IN1(\fpu_add_ctl/n941 ), .IN2(\fpu_add_ctl/n77 ), .QN(n2884) );
  INVX0 U5033 ( .INP(n4782), .ZN(n4727) );
  NOR2X0 U5034 ( .IN1(n4730), .IN2(n2983), .QN(n4782) );
  NAND3X0 U5035 ( .IN1(\fpu_add_frac_dp/n339 ), .IN2(\fpu_add_frac_dp/n235 ), 
        .IN3(\fpu_add_frac_dp/n426 ), .QN(n2983) );
  NAND4X0 U5036 ( .IN1(n4789), .IN2(n4790), .IN3(n4791), .IN4(n4792), .QN(
        n4730) );
  NOR2X0 U5037 ( .IN1(n4793), .IN2(n4794), .QN(n4792) );
  NAND4X0 U5038 ( .IN1(n2813), .IN2(n2809), .IN3(n2806), .IN4(n2804), .QN(
        n4794) );
  INVX0 U5039 ( .INP(n2800), .ZN(n2804) );
  NAND3X0 U5040 ( .IN1(\fpu_add_frac_dp/n362 ), .IN2(\fpu_add_frac_dp/n281 ), 
        .IN3(\fpu_add_frac_dp/n472 ), .QN(n2800) );
  INVX0 U5041 ( .INP(n2974), .ZN(n2806) );
  NAND3X0 U5042 ( .IN1(\fpu_add_frac_dp/n361 ), .IN2(\fpu_add_frac_dp/n279 ), 
        .IN3(\fpu_add_frac_dp/n470 ), .QN(n2974) );
  INVX0 U5043 ( .INP(n2975), .ZN(n2809) );
  NAND3X0 U5044 ( .IN1(\fpu_add_frac_dp/n360 ), .IN2(\fpu_add_frac_dp/n277 ), 
        .IN3(\fpu_add_frac_dp/n468 ), .QN(n2975) );
  INVX0 U5045 ( .INP(n2976), .ZN(n2813) );
  NAND3X0 U5046 ( .IN1(\fpu_add_frac_dp/n359 ), .IN2(\fpu_add_frac_dp/n275 ), 
        .IN3(\fpu_add_frac_dp/n466 ), .QN(n2976) );
  OR4X1 U5047 ( .IN1(n2798), .IN2(n2794), .IN3(n2792), .IN4(n2788), .Q(n4793)
         );
  NAND3X0 U5048 ( .IN1(\fpu_add_frac_dp/n366 ), .IN2(\fpu_add_frac_dp/n289 ), 
        .IN3(\fpu_add_frac_dp/n480 ), .QN(n2788) );
  NAND3X0 U5049 ( .IN1(\fpu_add_frac_dp/n365 ), .IN2(\fpu_add_frac_dp/n287 ), 
        .IN3(\fpu_add_frac_dp/n478 ), .QN(n2792) );
  NAND3X0 U5050 ( .IN1(\fpu_add_frac_dp/n364 ), .IN2(\fpu_add_frac_dp/n285 ), 
        .IN3(\fpu_add_frac_dp/n476 ), .QN(n2794) );
  NAND3X0 U5051 ( .IN1(\fpu_add_frac_dp/n363 ), .IN2(\fpu_add_frac_dp/n283 ), 
        .IN3(\fpu_add_frac_dp/n474 ), .QN(n2798) );
  NOR4X0 U5052 ( .IN1(n4795), .IN2(n2836), .IN3(n2830), .IN4(n2834), .QN(n4791) );
  NAND3X0 U5053 ( .IN1(\fpu_add_frac_dp/n353 ), .IN2(\fpu_add_frac_dp/n263 ), 
        .IN3(\fpu_add_frac_dp/n454 ), .QN(n2834) );
  NAND3X0 U5054 ( .IN1(\fpu_add_frac_dp/n354 ), .IN2(\fpu_add_frac_dp/n265 ), 
        .IN3(\fpu_add_frac_dp/n456 ), .QN(n2830) );
  NAND3X0 U5055 ( .IN1(\fpu_add_frac_dp/n352 ), .IN2(\fpu_add_frac_dp/n261 ), 
        .IN3(\fpu_add_frac_dp/n452 ), .QN(n2836) );
  NAND4X0 U5056 ( .IN1(n2828), .IN2(n2824), .IN3(n2821), .IN4(n2819), .QN(
        n4795) );
  INVX0 U5057 ( .INP(n2815), .ZN(n2819) );
  NAND3X0 U5058 ( .IN1(\fpu_add_frac_dp/n358 ), .IN2(\fpu_add_frac_dp/n273 ), 
        .IN3(\fpu_add_frac_dp/n464 ), .QN(n2815) );
  INVX0 U5059 ( .INP(n2977), .ZN(n2821) );
  NAND3X0 U5060 ( .IN1(\fpu_add_frac_dp/n357 ), .IN2(\fpu_add_frac_dp/n271 ), 
        .IN3(\fpu_add_frac_dp/n462 ), .QN(n2977) );
  INVX0 U5061 ( .INP(n2978), .ZN(n2824) );
  NAND3X0 U5062 ( .IN1(\fpu_add_frac_dp/n356 ), .IN2(\fpu_add_frac_dp/n269 ), 
        .IN3(\fpu_add_frac_dp/n460 ), .QN(n2978) );
  INVX0 U5063 ( .INP(n2979), .ZN(n2828) );
  NAND3X0 U5064 ( .IN1(\fpu_add_frac_dp/n355 ), .IN2(\fpu_add_frac_dp/n267 ), 
        .IN3(\fpu_add_frac_dp/n458 ), .QN(n2979) );
  NOR4X0 U5065 ( .IN1(n4796), .IN2(n2858), .IN3(n2852), .IN4(n2854), .QN(n4790) );
  NAND3X0 U5066 ( .IN1(\fpu_add_frac_dp/n346 ), .IN2(\fpu_add_frac_dp/n249 ), 
        .IN3(\fpu_add_frac_dp/n440 ), .QN(n2854) );
  NAND3X0 U5067 ( .IN1(\fpu_add_frac_dp/n347 ), .IN2(\fpu_add_frac_dp/n251 ), 
        .IN3(\fpu_add_frac_dp/n442 ), .QN(n2852) );
  NAND3X0 U5068 ( .IN1(\fpu_add_frac_dp/n345 ), .IN2(\fpu_add_frac_dp/n247 ), 
        .IN3(\fpu_add_frac_dp/n438 ), .QN(n2858) );
  OR4X1 U5069 ( .IN1(n2848), .IN2(n2846), .IN3(n2842), .IN4(n2840), .Q(n4796)
         );
  NAND3X0 U5070 ( .IN1(\fpu_add_frac_dp/n351 ), .IN2(\fpu_add_frac_dp/n259 ), 
        .IN3(\fpu_add_frac_dp/n450 ), .QN(n2840) );
  NAND3X0 U5071 ( .IN1(\fpu_add_frac_dp/n350 ), .IN2(\fpu_add_frac_dp/n257 ), 
        .IN3(\fpu_add_frac_dp/n448 ), .QN(n2842) );
  NAND3X0 U5072 ( .IN1(\fpu_add_frac_dp/n349 ), .IN2(\fpu_add_frac_dp/n255 ), 
        .IN3(\fpu_add_frac_dp/n446 ), .QN(n2846) );
  NAND3X0 U5073 ( .IN1(\fpu_add_frac_dp/n348 ), .IN2(\fpu_add_frac_dp/n253 ), 
        .IN3(\fpu_add_frac_dp/n444 ), .QN(n2848) );
  NOR4X0 U5074 ( .IN1(n4797), .IN2(n2973), .IN3(n2881), .IN4(n4735), .QN(n4789) );
  OR2X1 U5075 ( .IN1(n4731), .IN2(n2786), .Q(n4735) );
  NAND3X0 U5076 ( .IN1(\fpu_add_frac_dp/n367 ), .IN2(\fpu_add_frac_dp/n291 ), 
        .IN3(\fpu_add_frac_dp/n482 ), .QN(n2786) );
  NAND3X0 U5077 ( .IN1(\fpu_add_frac_dp/n340 ), .IN2(\fpu_add_frac_dp/n237 ), 
        .IN3(\fpu_add_frac_dp/n428 ), .QN(n2881) );
  NAND4X0 U5078 ( .IN1(n2873), .IN2(n2871), .IN3(n2865), .IN4(n2861), .QN(
        n4797) );
  INVX0 U5079 ( .INP(n2980), .ZN(n2861) );
  NAND3X0 U5080 ( .IN1(\fpu_add_frac_dp/n344 ), .IN2(\fpu_add_frac_dp/n245 ), 
        .IN3(\fpu_add_frac_dp/n436 ), .QN(n2980) );
  INVX0 U5081 ( .INP(n2981), .ZN(n2865) );
  NAND3X0 U5082 ( .IN1(\fpu_add_frac_dp/n343 ), .IN2(\fpu_add_frac_dp/n243 ), 
        .IN3(\fpu_add_frac_dp/n434 ), .QN(n2981) );
  INVX0 U5083 ( .INP(n2867), .ZN(n2871) );
  NAND3X0 U5084 ( .IN1(\fpu_add_frac_dp/n342 ), .IN2(\fpu_add_frac_dp/n241 ), 
        .IN3(\fpu_add_frac_dp/n432 ), .QN(n2867) );
  INVX0 U5085 ( .INP(n2982), .ZN(n2873) );
  NAND3X0 U5086 ( .IN1(\fpu_add_frac_dp/n341 ), .IN2(\fpu_add_frac_dp/n239 ), 
        .IN3(\fpu_add_frac_dp/n430 ), .QN(n2982) );
  MUX21X1 U5087 ( .IN1(\fpu_add_frac_dp/n582 ), .IN2(\fpu_add_ctl/n78 ), .S(
        \fpu_add_ctl/n322 ), .Q(n4786) );
  NOR2X0 U5088 ( .IN1(n4731), .IN2(n2973), .QN(n4785) );
  NAND3X0 U5089 ( .IN1(\fpu_add_frac_dp/n368 ), .IN2(\fpu_add_frac_dp/n293 ), 
        .IN3(\fpu_add_frac_dp/n484 ), .QN(n2973) );
  NAND4X0 U5090 ( .IN1(\fpu_add_frac_dp/n313 ), .IN2(n3074), .IN3(n4798), 
        .IN4(n4799), .QN(n4731) );
  NOR4X0 U5091 ( .IN1(n4800), .IN2(n2967), .IN3(n2964), .IN4(n2966), .QN(n4799) );
  NAND3X0 U5092 ( .IN1(\fpu_add_frac_dp/n375 ), .IN2(\fpu_add_frac_dp/n307 ), 
        .IN3(\fpu_add_frac_dp/n498 ), .QN(n2966) );
  NAND2X0 U5093 ( .IN1(\fpu_add_frac_dp/n377 ), .IN2(\fpu_add_frac_dp/n311 ), 
        .QN(n2964) );
  NAND3X0 U5094 ( .IN1(\fpu_add_frac_dp/n374 ), .IN2(\fpu_add_frac_dp/n305 ), 
        .IN3(\fpu_add_frac_dp/n496 ), .QN(n2967) );
  OR2X1 U5095 ( .IN1(n2969), .IN2(n2968), .Q(n4800) );
  NAND3X0 U5096 ( .IN1(\fpu_add_frac_dp/n373 ), .IN2(\fpu_add_frac_dp/n303 ), 
        .IN3(\fpu_add_frac_dp/n494 ), .QN(n2968) );
  NAND3X0 U5097 ( .IN1(\fpu_add_frac_dp/n372 ), .IN2(\fpu_add_frac_dp/n301 ), 
        .IN3(\fpu_add_frac_dp/n492 ), .QN(n2969) );
  NOR3X0 U5098 ( .IN1(n2972), .IN2(n2971), .IN3(n2970), .QN(n4798) );
  NAND3X0 U5099 ( .IN1(\fpu_add_frac_dp/n371 ), .IN2(\fpu_add_frac_dp/n299 ), 
        .IN3(\fpu_add_frac_dp/n490 ), .QN(n2970) );
  NAND3X0 U5100 ( .IN1(\fpu_add_frac_dp/n370 ), .IN2(\fpu_add_frac_dp/n297 ), 
        .IN3(\fpu_add_frac_dp/n488 ), .QN(n2971) );
  NAND3X0 U5101 ( .IN1(\fpu_add_frac_dp/n369 ), .IN2(\fpu_add_frac_dp/n295 ), 
        .IN3(\fpu_add_frac_dp/n486 ), .QN(n2972) );
  INVX0 U5102 ( .INP(n2965), .ZN(n3074) );
  NAND3X0 U5103 ( .IN1(\fpu_add_frac_dp/n376 ), .IN2(\fpu_add_frac_dp/n309 ), 
        .IN3(\fpu_add_frac_dp/n500 ), .QN(n2965) );
  AO22X1 U5104 ( .IN1(n4000), .IN2(n1325), .IN3(n1340), .IN4(n4801), .Q(
        \fpu_add_ctl/n540 ) );
  AO221X1 U5105 ( .IN1(n1737), .IN2(n4648), .IN3(n2047), .IN4(
        \fpu_add_ctl/n940 ), .IN5(n4048), .Q(n4801) );
  INVX0 U5106 ( .INP(n4065), .ZN(n4048) );
  NAND4X0 U5107 ( .IN1(n4410), .IN2(n4802), .IN3(n4803), .IN4(
        \fpu_add_ctl/n312 ), .QN(n4065) );
  INVX0 U5108 ( .INP(n4804), .ZN(n2047) );
  NAND3X0 U5109 ( .IN1(n4805), .IN2(n4070), .IN3(n4806), .QN(n4648) );
  XOR3X1 U5110 ( .IN1(\fpu_add_ctl/n125 ), .IN2(\fpu_add_ctl/n940 ), .IN3(
        n4396), .Q(n4806) );
  NOR2X0 U5111 ( .IN1(n1867), .IN2(\fpu_add_ctl/n318 ), .QN(n4396) );
  NAND2X0 U5112 ( .IN1(n1737), .IN2(n1741), .QN(n4805) );
  NAND2X0 U5113 ( .IN1(n1752), .IN2(n1753), .QN(n1741) );
  NAND2X0 U5114 ( .IN1(\fpu_add_ctl/n324 ), .IN2(n4807), .QN(n1753) );
  AO22X1 U5115 ( .IN1(n692), .IN2(n4613), .IN3(n325), .IN4(n4616), .Q(n4807)
         );
  NAND2X0 U5116 ( .IN1(\fpu_add_ctl/n127 ), .IN2(\fpu_add_ctl/n124 ), .QN(
        n4616) );
  NAND2X0 U5117 ( .IN1(\fpu_add_ctl/n332 ), .IN2(\fpu_add_ctl/n123 ), .QN(
        n4613) );
  NAND2X0 U5118 ( .IN1(n338), .IN2(n4808), .QN(n1752) );
  AO22X1 U5119 ( .IN1(n692), .IN2(n4614), .IN3(n325), .IN4(n4615), .Q(n4808)
         );
  NAND2X0 U5120 ( .IN1(\fpu_add_ctl/n119 ), .IN2(\fpu_add_ctl/n121 ), .QN(
        n4615) );
  NAND2X0 U5121 ( .IN1(\fpu_add_ctl/n118 ), .IN2(\fpu_add_ctl/n333 ), .QN(
        n4614) );
  INVX0 U5122 ( .INP(n1867), .ZN(n1737) );
  NAND2X0 U5123 ( .IN1(n4409), .IN2(n4400), .QN(n1867) );
  INVX0 U5124 ( .INP(n4114), .ZN(n4000) );
  INVX0 U5125 ( .INP(n4403), .ZN(\fpu_add_ctl/n47 ) );
  NAND2X0 U5126 ( .IN1(\fpu_add_ctl/n49 ), .IN2(n4418), .QN(n4403) );
  NOR2X0 U5127 ( .IN1(n4057), .IN2(\fpu_add_ctl/n210 ), .QN(\fpu_add_ctl/n49 )
         );
  NAND2X0 U5128 ( .IN1(\fpu_add_ctl/n470 ), .IN2(n1312), .QN(n4057) );
  INVX0 U5129 ( .INP(n4809), .ZN(\fpu_add_ctl/n441 ) );
  NAND2X0 U5130 ( .IN1(n1336), .IN2(n91), .QN(\fpu_add_ctl/n426 ) );
  NAND2X0 U5131 ( .IN1(n1334), .IN2(n562), .QN(\fpu_add_ctl/n425 ) );
  NAND2X0 U5132 ( .IN1(\fpu_add_ctl/n329 ), .IN2(n1335), .QN(
        \fpu_add_ctl/n416 ) );
  NAND2X0 U5133 ( .IN1(n3973), .IN2(\fpu_add_ctl/n470 ), .QN(n4114) );
  NOR3X0 U5134 ( .IN1(n4810), .IN2(se_add_exp), .IN3(\fpu_add_ctl/n210 ), .QN(
        \fpu_add_ctl/i_add_pipe_active/N7 ) );
  NOR4X0 U5135 ( .IN1(n4811), .IN2(n651), .IN3(\fpu_add_ctl/n325 ), .IN4(n4411), .QN(n4810) );
  NAND4X0 U5136 ( .IN1(n4812), .IN2(n4813), .IN3(n4814), .IN4(n4804), .QN(
        n4411) );
  NAND3X0 U5137 ( .IN1(n4815), .IN2(n158), .IN3(n4405), .QN(n4804) );
  OR2X1 U5138 ( .IN1(n4404), .IN2(n4410), .Q(n4815) );
  NOR2X0 U5139 ( .IN1(n595), .IN2(\fpu_add_ctl/n318 ), .QN(n4404) );
  NOR2X0 U5140 ( .IN1(n4816), .IN2(n2668), .QN(n4814) );
  NOR2X0 U5141 ( .IN1(n4389), .IN2(n4817), .QN(n2668) );
  NAND3X0 U5142 ( .IN1(n4818), .IN2(n4400), .IN3(n4406), .QN(n4813) );
  INVX0 U5143 ( .INP(n4817), .ZN(n4400) );
  AO21X1 U5144 ( .IN1(\fpu_add_ctl/n318 ), .IN2(n585), .IN3(n172), .Q(n4818)
         );
  NAND3X0 U5145 ( .IN1(n4405), .IN2(\fpu_add_ctl/n312 ), .IN3(n4410), .QN(
        n4812) );
  NOR2X0 U5146 ( .IN1(n18), .IN2(\fpu_add_ctl/n321 ), .QN(n4410) );
  AND2X1 U5147 ( .IN1(n4803), .IN2(\fpu_add_ctl/n936 ), .Q(n4405) );
  NOR3X0 U5148 ( .IN1(n84), .IN2(n172), .IN3(n585), .QN(n4803) );
  NAND3X0 U5149 ( .IN1(\fpu_add_ctl/n66 ), .IN2(\fpu_add_ctl/n269 ), .IN3(
        \fpu_add_ctl/n79 ), .QN(n4811) );
  AND2X1 U5150 ( .IN1(grst_l), .IN2(\fpu_add_ctl/n470 ), .Q(
        \fpu_add_ctl/dffrl_add_ctl/N4 ) );
  INVX0 U5151 ( .INP(se_add_exp), .ZN(\fpu_add_ctl/n470 ) );
  AO222X1 U5152 ( .IN1(n4819), .IN2(n347), .IN3(n4820), .IN4(n885), .IN5(n3973), .IN6(\fpu_add_ctl/add_id_out[9] ), .Q(add_id_out_in[9]) );
  AO222X1 U5153 ( .IN1(n4819), .IN2(n348), .IN3(n4820), .IN4(n886), .IN5(n3973), .IN6(\fpu_add_ctl/add_id_out[8] ), .Q(add_id_out_in[8]) );
  AO222X1 U5154 ( .IN1(n4819), .IN2(n349), .IN3(n4820), .IN4(n887), .IN5(n3973), .IN6(\fpu_add_ctl/add_id_out[7] ), .Q(add_id_out_in[7]) );
  AO222X1 U5155 ( .IN1(n4819), .IN2(n350), .IN3(n4820), .IN4(n888), .IN5(n3973), .IN6(\fpu_add_ctl/add_id_out[6] ), .Q(add_id_out_in[6]) );
  AO222X1 U5156 ( .IN1(n4819), .IN2(n351), .IN3(n4820), .IN4(n889), .IN5(n3973), .IN6(\fpu_add_ctl/add_id_out[5] ), .Q(add_id_out_in[5]) );
  AO222X1 U5157 ( .IN1(n4819), .IN2(n352), .IN3(n4820), .IN4(n890), .IN5(n3973), .IN6(\fpu_add_ctl/add_id_out[4] ), .Q(add_id_out_in[4]) );
  AO222X1 U5158 ( .IN1(n4819), .IN2(n353), .IN3(n4820), .IN4(n891), .IN5(n3973), .IN6(\fpu_add_ctl/add_id_out[3] ), .Q(add_id_out_in[3]) );
  AO222X1 U5159 ( .IN1(n4819), .IN2(n354), .IN3(n4820), .IN4(n892), .IN5(n3973), .IN6(\fpu_add_ctl/add_id_out[2] ), .Q(add_id_out_in[2]) );
  AO222X1 U5160 ( .IN1(n4819), .IN2(n341), .IN3(n4820), .IN4(n893), .IN5(n3973), .IN6(\fpu_add_ctl/add_id_out[1] ), .Q(add_id_out_in[1]) );
  AO222X1 U5161 ( .IN1(n4819), .IN2(n342), .IN3(n4820), .IN4(n894), .IN5(n3973), .IN6(\fpu_add_ctl/add_id_out[0] ), .Q(add_id_out_in[0]) );
  NOR2X0 U5162 ( .IN1(n3973), .IN2(\fpu_add_ctl/n315 ), .QN(n4820) );
  NOR2X0 U5163 ( .IN1(n622), .IN2(n3973), .QN(n4819) );
  AO221X1 U5164 ( .IN1(n536), .IN2(n1306), .IN3(n1002), .IN4(n1308), .IN5(
        n1315), .Q(add_frac_out[9]) );
  AO221X1 U5165 ( .IN1(n537), .IN2(n1305), .IN3(n1003), .IN4(n65), .IN5(n1315), 
        .Q(add_frac_out[8]) );
  AO221X1 U5166 ( .IN1(n538), .IN2(n1307), .IN3(n1310), .IN4(n919), .IN5(n1315), .Q(add_frac_out[7]) );
  AO221X1 U5167 ( .IN1(n539), .IN2(n66), .IN3(n1309), .IN4(n920), .IN5(n1315), 
        .Q(add_frac_out[6]) );
  AO221X1 U5168 ( .IN1(n467), .IN2(n1308), .IN3(n1307), .IN4(n859), .IN5(n1315), .Q(add_frac_out[63]) );
  AO221X1 U5169 ( .IN1(n468), .IN2(n1310), .IN3(n66), .IN4(n907), .IN5(n4821), 
        .Q(add_frac_out[62]) );
  AO21X1 U5170 ( .IN1(n1006), .IN2(n579), .IN3(n1316), .Q(n4821) );
  AO221X1 U5171 ( .IN1(n963), .IN2(n65), .IN3(n1306), .IN4(n493), .IN5(n4822), 
        .Q(add_frac_out[61]) );
  AO21X1 U5172 ( .IN1(n1035), .IN2(n579), .IN3(n1317), .Q(n4822) );
  AO221X1 U5173 ( .IN1(n466), .IN2(n1309), .IN3(n1305), .IN4(n860), .IN5(n4823), .Q(add_frac_out[60]) );
  AO21X1 U5174 ( .IN1(n1036), .IN2(n579), .IN3(n1318), .Q(n4823) );
  AO221X1 U5175 ( .IN1(n540), .IN2(n1306), .IN3(n1308), .IN4(n921), .IN5(n1315), .Q(add_frac_out[5]) );
  AO221X1 U5176 ( .IN1(n933), .IN2(n1308), .IN3(n1307), .IN4(n494), .IN5(n4824), .Q(add_frac_out[59]) );
  AO21X1 U5177 ( .IN1(n1037), .IN2(n579), .IN3(n1316), .Q(n4824) );
  AO221X1 U5178 ( .IN1(n1309), .IN2(n1034), .IN3(n66), .IN4(n495), .IN5(n4825), 
        .Q(add_frac_out[58]) );
  AO21X1 U5179 ( .IN1(n1038), .IN2(n579), .IN3(n1317), .Q(n4825) );
  AO221X1 U5180 ( .IN1(n65), .IN2(n906), .IN3(n1306), .IN4(n496), .IN5(n4826), 
        .Q(add_frac_out[57]) );
  AO21X1 U5181 ( .IN1(n1039), .IN2(n579), .IN3(n1318), .Q(n4826) );
  AO221X1 U5182 ( .IN1(n1310), .IN2(n1064), .IN3(n1305), .IN4(n497), .IN5(
        n4827), .Q(add_frac_out[56]) );
  AO21X1 U5183 ( .IN1(n1040), .IN2(n579), .IN3(n1316), .Q(n4827) );
  AO221X1 U5184 ( .IN1(n1309), .IN2(n918), .IN3(n1307), .IN4(n498), .IN5(n4828), .Q(add_frac_out[55]) );
  AO21X1 U5185 ( .IN1(n1041), .IN2(n579), .IN3(n1317), .Q(n4828) );
  AO221X1 U5186 ( .IN1(n964), .IN2(n579), .IN3(n66), .IN4(n499), .IN5(n4829), 
        .Q(add_frac_out[54]) );
  AO21X1 U5187 ( .IN1(n909), .IN2(n1309), .IN3(n1318), .Q(n4829) );
  AO221X1 U5188 ( .IN1(n965), .IN2(n579), .IN3(n1306), .IN4(n500), .IN5(n4830), 
        .Q(add_frac_out[53]) );
  AO21X1 U5189 ( .IN1(n910), .IN2(n1308), .IN3(n1316), .Q(n4830) );
  AO221X1 U5190 ( .IN1(n966), .IN2(n579), .IN3(n1305), .IN4(n501), .IN5(n4831), 
        .Q(add_frac_out[52]) );
  AO21X1 U5191 ( .IN1(n911), .IN2(n1310), .IN3(n1317), .Q(n4831) );
  AO221X1 U5192 ( .IN1(n967), .IN2(n579), .IN3(n1307), .IN4(n502), .IN5(n4832), 
        .Q(add_frac_out[51]) );
  AO21X1 U5193 ( .IN1(n912), .IN2(n65), .IN3(n1318), .Q(n4832) );
  AO221X1 U5194 ( .IN1(n968), .IN2(n579), .IN3(n66), .IN4(n503), .IN5(n4833), 
        .Q(add_frac_out[50]) );
  AO21X1 U5195 ( .IN1(n913), .IN2(n1309), .IN3(n1316), .Q(n4833) );
  AO221X1 U5196 ( .IN1(n541), .IN2(n1305), .IN3(n65), .IN4(n922), .IN5(n1315), 
        .Q(add_frac_out[4]) );
  AO221X1 U5197 ( .IN1(n469), .IN2(n1310), .IN3(n1306), .IN4(n861), .IN5(n4834), .Q(add_frac_out[49]) );
  AO21X1 U5198 ( .IN1(n1042), .IN2(n579), .IN3(n1317), .Q(n4834) );
  AO221X1 U5199 ( .IN1(n470), .IN2(n65), .IN3(n1305), .IN4(n862), .IN5(n4835), 
        .Q(add_frac_out[48]) );
  AO21X1 U5200 ( .IN1(n1043), .IN2(n579), .IN3(n1318), .Q(n4835) );
  AO221X1 U5201 ( .IN1(n471), .IN2(n1309), .IN3(n1307), .IN4(n863), .IN5(n4836), .Q(add_frac_out[47]) );
  AO21X1 U5202 ( .IN1(n1044), .IN2(n579), .IN3(n1316), .Q(n4836) );
  AO221X1 U5203 ( .IN1(n472), .IN2(n1308), .IN3(n66), .IN4(n864), .IN5(n4837), 
        .Q(add_frac_out[46]) );
  AO21X1 U5204 ( .IN1(n1045), .IN2(n579), .IN3(n1317), .Q(n4837) );
  AO221X1 U5205 ( .IN1(n473), .IN2(n1310), .IN3(n1306), .IN4(n865), .IN5(n4838), .Q(add_frac_out[45]) );
  AO21X1 U5206 ( .IN1(n1046), .IN2(n579), .IN3(n1318), .Q(n4838) );
  AO221X1 U5207 ( .IN1(n474), .IN2(n65), .IN3(n1305), .IN4(n866), .IN5(n4839), 
        .Q(add_frac_out[44]) );
  AO21X1 U5208 ( .IN1(n1047), .IN2(n579), .IN3(n1316), .Q(n4839) );
  AO221X1 U5209 ( .IN1(n475), .IN2(n1309), .IN3(n1307), .IN4(n867), .IN5(n4840), .Q(add_frac_out[43]) );
  AO21X1 U5210 ( .IN1(n1048), .IN2(n579), .IN3(n1317), .Q(n4840) );
  AO221X1 U5211 ( .IN1(n476), .IN2(n1308), .IN3(n66), .IN4(n868), .IN5(n4841), 
        .Q(add_frac_out[42]) );
  AO21X1 U5212 ( .IN1(n1049), .IN2(n579), .IN3(n1318), .Q(n4841) );
  AO221X1 U5213 ( .IN1(n477), .IN2(n1310), .IN3(n1306), .IN4(n869), .IN5(n4842), .Q(add_frac_out[41]) );
  AO21X1 U5214 ( .IN1(n1050), .IN2(n579), .IN3(n1316), .Q(n4842) );
  AO221X1 U5215 ( .IN1(n478), .IN2(n65), .IN3(n1305), .IN4(n870), .IN5(n4843), 
        .Q(add_frac_out[40]) );
  AO21X1 U5216 ( .IN1(n1051), .IN2(n579), .IN3(n1317), .Q(n4843) );
  AO221X1 U5217 ( .IN1(n542), .IN2(n1307), .IN3(n1310), .IN4(n923), .IN5(n1315), .Q(add_frac_out[3]) );
  AO221X1 U5218 ( .IN1(n479), .IN2(n1309), .IN3(n1307), .IN4(n871), .IN5(n4844), .Q(add_frac_out[39]) );
  AO21X1 U5219 ( .IN1(n1052), .IN2(n579), .IN3(n1318), .Q(n4844) );
  AO221X1 U5220 ( .IN1(n480), .IN2(n1308), .IN3(n66), .IN4(n872), .IN5(n4845), 
        .Q(add_frac_out[38]) );
  AO21X1 U5221 ( .IN1(n1053), .IN2(n579), .IN3(n1316), .Q(n4845) );
  AO221X1 U5222 ( .IN1(n481), .IN2(n1310), .IN3(n1306), .IN4(n873), .IN5(n4846), .Q(add_frac_out[37]) );
  AO21X1 U5223 ( .IN1(n1054), .IN2(n579), .IN3(n1317), .Q(n4846) );
  AO221X1 U5224 ( .IN1(n482), .IN2(n65), .IN3(n1305), .IN4(n874), .IN5(n4847), 
        .Q(add_frac_out[36]) );
  AO21X1 U5225 ( .IN1(n1055), .IN2(n579), .IN3(n1318), .Q(n4847) );
  AO221X1 U5226 ( .IN1(n483), .IN2(n1309), .IN3(n1307), .IN4(n875), .IN5(n4848), .Q(add_frac_out[35]) );
  AO21X1 U5227 ( .IN1(n1056), .IN2(n579), .IN3(n1316), .Q(n4848) );
  AO221X1 U5228 ( .IN1(n484), .IN2(n1308), .IN3(n66), .IN4(n876), .IN5(n4849), 
        .Q(add_frac_out[34]) );
  AO21X1 U5229 ( .IN1(n1057), .IN2(n579), .IN3(n1317), .Q(n4849) );
  AO221X1 U5230 ( .IN1(n485), .IN2(n1310), .IN3(n1306), .IN4(n877), .IN5(n4850), .Q(add_frac_out[33]) );
  AO21X1 U5231 ( .IN1(n1058), .IN2(n579), .IN3(n1318), .Q(n4850) );
  AO221X1 U5232 ( .IN1(n486), .IN2(n65), .IN3(n1305), .IN4(n878), .IN5(n4851), 
        .Q(add_frac_out[32]) );
  AO21X1 U5233 ( .IN1(n1059), .IN2(n579), .IN3(n1316), .Q(n4851) );
  AO221X1 U5234 ( .IN1(n487), .IN2(n1309), .IN3(n1307), .IN4(n879), .IN5(n4852), .Q(add_frac_out[31]) );
  AO21X1 U5235 ( .IN1(n1060), .IN2(n579), .IN3(n1317), .Q(n4852) );
  AO221X1 U5236 ( .IN1(n488), .IN2(n1308), .IN3(n66), .IN4(n880), .IN5(n4853), 
        .Q(add_frac_out[30]) );
  AO21X1 U5237 ( .IN1(n1061), .IN2(n579), .IN3(n1318), .Q(n4853) );
  AO221X1 U5238 ( .IN1(n543), .IN2(n66), .IN3(n1308), .IN4(n924), .IN5(n1315), 
        .Q(add_frac_out[2]) );
  AO221X1 U5239 ( .IN1(n489), .IN2(n65), .IN3(n1306), .IN4(n881), .IN5(n4854), 
        .Q(add_frac_out[29]) );
  AO21X1 U5240 ( .IN1(n1062), .IN2(n579), .IN3(n1316), .Q(n4854) );
  AO221X1 U5241 ( .IN1(n969), .IN2(n579), .IN3(n517), .IN4(n1310), .IN5(n4855), 
        .Q(add_frac_out[28]) );
  AO21X1 U5242 ( .IN1(n938), .IN2(n1306), .IN3(n1317), .Q(n4855) );
  AO221X1 U5243 ( .IN1(n970), .IN2(n579), .IN3(n518), .IN4(n1309), .IN5(n4856), 
        .Q(add_frac_out[27]) );
  AO21X1 U5244 ( .IN1(n939), .IN2(n1307), .IN3(n1318), .Q(n4856) );
  AO221X1 U5245 ( .IN1(n971), .IN2(n579), .IN3(n519), .IN4(n1308), .IN5(n4857), 
        .Q(add_frac_out[26]) );
  AO21X1 U5246 ( .IN1(n940), .IN2(n66), .IN3(n1316), .Q(n4857) );
  AO221X1 U5247 ( .IN1(n972), .IN2(n579), .IN3(n520), .IN4(n65), .IN5(n4858), 
        .Q(add_frac_out[25]) );
  AO21X1 U5248 ( .IN1(n941), .IN2(n1305), .IN3(n1317), .Q(n4858) );
  AO221X1 U5249 ( .IN1(n973), .IN2(n579), .IN3(n521), .IN4(n1310), .IN5(n4859), 
        .Q(add_frac_out[24]) );
  AO21X1 U5250 ( .IN1(n942), .IN2(n1306), .IN3(n1318), .Q(n4859) );
  AO221X1 U5251 ( .IN1(n974), .IN2(n579), .IN3(n522), .IN4(n1309), .IN5(n4860), 
        .Q(add_frac_out[23]) );
  AO21X1 U5252 ( .IN1(n943), .IN2(n1307), .IN3(n1316), .Q(n4860) );
  AO221X1 U5253 ( .IN1(n975), .IN2(n579), .IN3(n523), .IN4(n1308), .IN5(n4861), 
        .Q(add_frac_out[22]) );
  AO21X1 U5254 ( .IN1(n944), .IN2(n66), .IN3(n1317), .Q(n4861) );
  AO221X1 U5255 ( .IN1(n976), .IN2(n579), .IN3(n524), .IN4(n65), .IN5(n4862), 
        .Q(add_frac_out[21]) );
  AO21X1 U5256 ( .IN1(n945), .IN2(n1305), .IN3(n1318), .Q(n4862) );
  AO221X1 U5257 ( .IN1(n977), .IN2(n579), .IN3(n525), .IN4(n1310), .IN5(n4863), 
        .Q(add_frac_out[20]) );
  AO21X1 U5258 ( .IN1(n946), .IN2(n1306), .IN3(n1316), .Q(n4863) );
  AO221X1 U5259 ( .IN1(n978), .IN2(n1306), .IN3(n65), .IN4(n551), .IN5(n1315), 
        .Q(add_frac_out[1]) );
  AO221X1 U5260 ( .IN1(n979), .IN2(n579), .IN3(n526), .IN4(n1309), .IN5(n4864), 
        .Q(add_frac_out[19]) );
  AO21X1 U5261 ( .IN1(n947), .IN2(n1307), .IN3(n1317), .Q(n4864) );
  AO221X1 U5262 ( .IN1(n980), .IN2(n579), .IN3(n527), .IN4(n1308), .IN5(n4865), 
        .Q(add_frac_out[18]) );
  AO21X1 U5263 ( .IN1(n948), .IN2(n66), .IN3(n1318), .Q(n4865) );
  AO221X1 U5264 ( .IN1(n981), .IN2(n579), .IN3(n528), .IN4(n65), .IN5(n4866), 
        .Q(add_frac_out[17]) );
  AO21X1 U5265 ( .IN1(n949), .IN2(n1305), .IN3(n1316), .Q(n4866) );
  AO221X1 U5266 ( .IN1(n982), .IN2(n579), .IN3(n529), .IN4(n1310), .IN5(n4867), 
        .Q(add_frac_out[16]) );
  AO21X1 U5267 ( .IN1(n950), .IN2(n1306), .IN3(n1317), .Q(n4867) );
  AO221X1 U5268 ( .IN1(n983), .IN2(n579), .IN3(n530), .IN4(n1309), .IN5(n4868), 
        .Q(add_frac_out[15]) );
  AO21X1 U5269 ( .IN1(n951), .IN2(n1307), .IN3(n1318), .Q(n4868) );
  AO221X1 U5270 ( .IN1(n984), .IN2(n579), .IN3(n531), .IN4(n1308), .IN5(n4869), 
        .Q(add_frac_out[14]) );
  AO21X1 U5271 ( .IN1(n952), .IN2(n66), .IN3(n1316), .Q(n4869) );
  AO221X1 U5272 ( .IN1(n985), .IN2(n579), .IN3(n532), .IN4(n65), .IN5(n4870), 
        .Q(add_frac_out[13]) );
  AO21X1 U5273 ( .IN1(n953), .IN2(n1305), .IN3(n1317), .Q(n4870) );
  AO221X1 U5274 ( .IN1(n986), .IN2(n579), .IN3(n533), .IN4(n1310), .IN5(n4871), 
        .Q(add_frac_out[12]) );
  AO21X1 U5275 ( .IN1(n954), .IN2(n1307), .IN3(n1315), .Q(n4871) );
  AO221X1 U5276 ( .IN1(n987), .IN2(n579), .IN3(n534), .IN4(n1309), .IN5(n4872), 
        .Q(add_frac_out[11]) );
  AO21X1 U5277 ( .IN1(n955), .IN2(n66), .IN3(n1315), .Q(n4872) );
  AO221X1 U5278 ( .IN1(n908), .IN2(n1305), .IN3(n535), .IN4(n1308), .IN5(n1315), .Q(add_frac_out[10]) );
  AO221X1 U5279 ( .IN1(n544), .IN2(n1305), .IN3(n1310), .IN4(n925), .IN5(n1315), .Q(add_frac_out[0]) );
  NAND3X0 U5280 ( .IN1(n441), .IN2(n758), .IN3(n4873), .QN(add_exp_out[9]) );
  NAND2X0 U5281 ( .IN1(\fpu_add_exp_dp/n2 ), .IN2(\fpu_add_exp_dp/n13 ), .QN(
        n4873) );
  NAND3X0 U5282 ( .IN1(n442), .IN2(n759), .IN3(n4874), .QN(add_exp_out[8]) );
  NAND2X0 U5283 ( .IN1(\fpu_add_exp_dp/n3 ), .IN2(\fpu_add_exp_dp/n14 ), .QN(
        n4874) );
  NAND3X0 U5284 ( .IN1(n732), .IN2(n434), .IN3(n4875), .QN(add_exp_out[7]) );
  NAND2X0 U5285 ( .IN1(\fpu_add_exp_dp/n4 ), .IN2(\fpu_add_exp_dp/n15 ), .QN(
        n4875) );
  NAND3X0 U5286 ( .IN1(n733), .IN2(n435), .IN3(n4876), .QN(add_exp_out[6]) );
  NAND2X0 U5287 ( .IN1(\fpu_add_exp_dp/n5 ), .IN2(\fpu_add_exp_dp/n16 ), .QN(
        n4876) );
  NAND3X0 U5288 ( .IN1(n734), .IN2(n436), .IN3(n4877), .QN(add_exp_out[5]) );
  NAND2X0 U5289 ( .IN1(\fpu_add_exp_dp/n6 ), .IN2(\fpu_add_exp_dp/n17 ), .QN(
        n4877) );
  NAND3X0 U5290 ( .IN1(n735), .IN2(n437), .IN3(n4878), .QN(add_exp_out[4]) );
  NAND2X0 U5291 ( .IN1(\fpu_add_exp_dp/n7 ), .IN2(\fpu_add_exp_dp/n18 ), .QN(
        n4878) );
  NAND3X0 U5292 ( .IN1(n736), .IN2(n438), .IN3(n4879), .QN(add_exp_out[3]) );
  NAND2X0 U5293 ( .IN1(\fpu_add_exp_dp/n8 ), .IN2(\fpu_add_exp_dp/n19 ), .QN(
        n4879) );
  NAND3X0 U5294 ( .IN1(n737), .IN2(n439), .IN3(n4880), .QN(add_exp_out[2]) );
  NAND2X0 U5295 ( .IN1(\fpu_add_exp_dp/n9 ), .IN2(\fpu_add_exp_dp/n20 ), .QN(
        n4880) );
  NAND3X0 U5296 ( .IN1(n738), .IN2(n440), .IN3(n4881), .QN(add_exp_out[1]) );
  NAND2X0 U5297 ( .IN1(\fpu_add_exp_dp/n21 ), .IN2(\fpu_add_exp_dp/n10 ), .QN(
        n4881) );
  NAND3X0 U5298 ( .IN1(n443), .IN2(n760), .IN3(n4882), .QN(add_exp_out[10]) );
  NAND2X0 U5299 ( .IN1(\fpu_add_exp_dp/n12 ), .IN2(\fpu_add_exp_dp/n1 ), .QN(
        n4882) );
  NAND3X0 U5300 ( .IN1(n764), .IN2(n454), .IN3(n4883), .QN(add_exp_out[0]) );
  NAND2X0 U5301 ( .IN1(\fpu_add_exp_dp/n22 ), .IN2(\fpu_add_exp_dp/n11 ), .QN(
        n4883) );
  INVX0 U5302 ( .INP(n4884), .ZN(add_exc_out[3]) );
  NAND2X0 U5303 ( .IN1(\fpu_add_ctl/n2 ), .IN2(n4884), .QN(add_exc_out[0]) );
  OA21X1 U5304 ( .IN1(\fpu_add_ctl/n5 ), .IN2(\fpu_add_frac_dp/n129 ), .IN3(
        \fpu_add_ctl/n4 ), .Q(n4884) );
  AOI21X1 U5305 ( .IN1(n1314), .IN2(n4809), .IN3(\fpu_add_ctl/n210 ), .QN(
        a6stg_fadd_in) );
  MUX21X1 U5306 ( .IN1(\fpu_add_ctl/n66 ), .IN2(n4885), .S(\fpu_add_ctl/n315 ), 
        .Q(n4809) );
  NAND2X0 U5307 ( .IN1(n642), .IN2(n339), .QN(n4885) );
  INVX0 U5308 ( .INP(n4417), .ZN(a1stg_step) );
  NAND2X0 U5309 ( .IN1(n4418), .IN2(n1313), .QN(n4417) );
  NOR2X0 U5310 ( .IN1(\fpu_add_ctl/n269 ), .IN2(add_dest_rdy), .QN(n3973) );
  NAND2X0 U5311 ( .IN1(n355), .IN2(n4886), .QN(n4418) );
  NAND4X0 U5312 ( .IN1(\fpu_add_ctl/n936 ), .IN2(\fpu_add_ctl/n314 ), .IN3(
        n4887), .IN4(n158), .QN(n4886) );
  NAND2X0 U5313 ( .IN1(\fpu_add_ctl/n318 ), .IN2(\fpu_add_ctl/n312 ), .QN(
        n4887) );
  NOR2X0 U5314 ( .IN1(n4394), .IN2(n4817), .QN(a1stg_fsdtoix) );
  NOR2X0 U5315 ( .IN1(n4802), .IN2(n4408), .QN(n4817) );
  AND2X1 U5316 ( .IN1(n4391), .IN2(n4389), .Q(n4394) );
  NAND3X0 U5317 ( .IN1(\fpu_add_ctl/n303 ), .IN2(n254), .IN3(n4888), .QN(n4389) );
  NAND3X0 U5318 ( .IN1(\fpu_add_ctl/n312 ), .IN2(n585), .IN3(n4888), .QN(n4391) );
  NOR4X0 U5319 ( .IN1(n595), .IN2(n84), .IN3(n172), .IN4(n18), .QN(n4888) );
  INVX0 U5320 ( .INP(n4070), .ZN(a1stg_fdtos) );
  NAND2X0 U5321 ( .IN1(n4816), .IN2(\fpu_add_ctl/n314 ), .QN(n4070) );
  INVX0 U5322 ( .INP(n4656), .ZN(n4816) );
  NAND4X0 U5323 ( .IN1(n4408), .IN2(\fpu_add_ctl/n303 ), .IN3(n4406), .IN4(n18), .QN(n4656) );
  INVX0 U5324 ( .INP(n4390), .ZN(n4408) );
  NAND2X0 U5325 ( .IN1(n158), .IN2(n829), .QN(n4390) );
  INVX0 U5326 ( .INP(n4046), .ZN(a1stg_faddsubs) );
  NAND2X0 U5327 ( .IN1(n4802), .IN2(n4409), .QN(n4046) );
  AND3X1 U5328 ( .IN1(n4406), .IN2(n172), .IN3(\fpu_add_ctl/n303 ), .Q(n4409)
         );
  NOR3X0 U5329 ( .IN1(n84), .IN2(n254), .IN3(n595), .QN(n4406) );
  INVX0 U5330 ( .INP(n4392), .ZN(n4802) );
  NAND2X0 U5331 ( .IN1(\fpu_add_ctl/n320 ), .IN2(\fpu_add_ctl/n936 ), .QN(
        n4392) );
endmodule

