
module fpu_div ( inq_op, inq_rnd_mode, inq_id, inq_in1, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0, 
        inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_div, 
        div_dest_rdy, fdiv_clken_l, fdiv_clken_l_div_exp_buf1, arst_l, grst_l, 
        rclk, div_pipe_active, d1stg_step, d8stg_fdiv_in, div_id_out_in, 
        div_exc_out, d8stg_fdivd, d8stg_fdivs, div_sign_out, div_exp_outa, 
        div_frac_outa, se, si, so );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  output [9:0] div_id_out_in;
  output [4:0] div_exc_out;
  output [10:0] div_exp_outa;
  output [51:0] div_frac_outa;
  input inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0,
         inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_53_0_neq_0,
         inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0,
         inq_in2_exp_neq_ffs, inq_div, div_dest_rdy, fdiv_clken_l,
         fdiv_clken_l_div_exp_buf1, arst_l, grst_l, rclk, se, si;
  output div_pipe_active, d1stg_step, d8stg_fdiv_in, d8stg_fdivd, d8stg_fdivs,
         div_sign_out, so;
  wire   d234stg_fdiv, d3stg_fdiv, d6stg_fdivs, d7stg_fdivd,
         div_expadd1_in1_dbl, div_expadd1_in1_sng, div_expadd1_in2_exp_in2_dbl,
         div_expadd1_in2_exp_in2_sng, div_expadd2_in1_exp_out,
         div_expadd2_no_decr_inv, \fpu_div_ctl/div_nx_out ,
         \fpu_div_ctl/div_id_out[9] , \fpu_div_ctl/div_id_out[8] ,
         \fpu_div_ctl/div_id_out[7] , \fpu_div_ctl/div_id_out[6] ,
         \fpu_div_ctl/div_id_out[5] , \fpu_div_ctl/div_id_out[4] ,
         \fpu_div_ctl/div_id_out[3] , \fpu_div_ctl/div_id_out[2] ,
         \fpu_div_ctl/div_id_out[1] , \fpu_div_ctl/div_id_out[0] ,
         \fpu_div_ctl/div_rnd_mode[1] , \fpu_div_ctl/div_cnt[0] ,
         \fpu_div_ctl/d3stg_opdec[1] , \fpu_div_ctl/d3stg_opdec[0] ,
         \fpu_div_ctl/d1stg_op[2] , \fpu_div_ctl/d1stg_op[3] ,
         \fpu_div_ctl/d1stg_op[4] , \fpu_div_ctl/d1stg_op[6] ,
         \fpu_div_ctl/d1stg_op[7] , \fpu_div_ctl/d1stg_div ,
         \fpu_div_ctl/d2stg_2zero_in , \fpu_div_ctl/d2stg_zero_in ,
         \fpu_div_ctl/d2stg_zero_in2 , \fpu_div_ctl/d2stg_infnan_in ,
         \fpu_div_ctl/d2stg_2inf_in , \fpu_div_ctl/d2stg_inf_in1 ,
         \fpu_div_ctl/d2stg_nan_in , \fpu_div_ctl/d2stg_nan_in2 ,
         \fpu_div_ctl/d2stg_snan_in1 , \fpu_div_ctl/d2stg_norm_dbl_in2 ,
         \fpu_div_ctl/d2stg_norm_sng_in2 , \fpu_div_ctl/d2stg_denorm_dbl_in2 ,
         \fpu_div_ctl/d2stg_denorm_sng_in2 , \fpu_div_ctl/d1stg_dblopa[4] ,
         \fpu_div_ctl/d1stg_sngopa[4] , \fpu_div_ctl/dffrl_div_ctl/N4 ,
         \fpu_div_ctl/i_d2stg_denorm_sng_in2/N3 ,
         \fpu_div_ctl/i_d2stg_denorm_dbl_in2/N3 ,
         \fpu_div_ctl/i_d2stg_norm_sng_in2/N3 ,
         \fpu_div_ctl/i_d2stg_norm_dbl_in2/N3 ,
         \fpu_div_ctl/i_d2stg_snan_in1/N3 , \fpu_div_ctl/i_d2stg_qnan_in1/N3 ,
         \fpu_div_ctl/i_d2stg_nan_in2/N3 , \fpu_div_ctl/i_d2stg_nan_in/N3 ,
         \fpu_div_ctl/i_d2stg_inf_in1/N3 , \fpu_div_ctl/i_d2stg_2inf_in/N3 ,
         \fpu_div_ctl/i_d2stg_zero_in2/N3 , \fpu_div_ctl/i_d2stg_2zero_in/N3 ,
         \fpu_div_ctl/i_d1stg_op/N21 , \fpu_div_ctl/i_d1stg_op/N20 ,
         \fpu_div_ctl/i_d1stg_op/N19 , \fpu_div_ctl/i_d1stg_op/N18 ,
         \fpu_div_ctl/i_d1stg_op/N17 , \fpu_div_ctl/i_d1stg_op/N16 ,
         \fpu_div_ctl/i_d1stg_op/N15 , \fpu_div_ctl/i_d1stg_op/N14 ,
         \fpu_div_ctl/i_d1stg_div/N7 , \fpu_div_ctl/i_d2stg_opdec/N11 ,
         \fpu_div_ctl/i_d234stg_fdiv/N7 , \fpu_div_ctl/i_d3stg_opdec/N11 ,
         \fpu_div_ctl/i_d3stg_opdec/N10 , \fpu_div_ctl/i_d3stg_opdec/N9 ,
         \fpu_div_ctl/i_d4stg_opdec/N11 , \fpu_div_ctl/i_d6stg_opdec/N11 ,
         \fpu_div_ctl/i_d6stg_opdec/N10 , \fpu_div_ctl/i_d6stg_opdec/N9 ,
         \fpu_div_ctl/i_d7stg_opdec/N11 , \fpu_div_ctl/i_d7stg_opdec/N9 ,
         \fpu_div_ctl/i_div_pipe_active/N7 ,
         \fpu_div_ctl/i_div_expadd1_in1_dbl/N3 ,
         \fpu_div_ctl/i_div_expadd1_in1_sng/N3 ,
         \fpu_div_ctl/i_div_expadd2_in1_exp_out/N7 ,
         \fpu_div_exp_dp/ckbuf_div_exp_dp/clken ,
         \fpu_div_exp_dp/ckbuf_div_exp_dp/N1 , n2, n14, n15, n16, n17, n18,
         n19, n21, n22, n25, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n40, n41, n47, n50, n52, n54, n58, n59, n86, n88, n89, n90, n93, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n117, n124, n125, n126, n127, n131, n138, n141, n142, n144, n145,
         n146, n148, n149, n150, n151, n152, n164, n168, n173, n177, n179,
         n181, n182, n184, n185, n191, n192, n193, n194, n196, n201, n205,
         n208, n209, n218, n246, n247, n248, n253, n272, n282, n285, n286,
         n289, n290, n291, n292, n351, n352, n354, n355, n370, n373, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n520, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n939, n979, n1047, n1349, n1351, n1353, n1354, n1355,
         n1356, \fpu_div_frac_dp/n2333 , \fpu_div_frac_dp/n2330 ,
         \fpu_div_frac_dp/n609 , \fpu_div_frac_dp/n602 ,
         \fpu_div_frac_dp/n997 , \fpu_div_frac_dp/n996 ,
         \fpu_div_frac_dp/n995 , \fpu_div_frac_dp/n994 ,
         \fpu_div_frac_dp/n993 , \fpu_div_frac_dp/n992 ,
         \fpu_div_frac_dp/n991 , \fpu_div_frac_dp/n990 ,
         \fpu_div_frac_dp/n989 , \fpu_div_frac_dp/n988 ,
         \fpu_div_frac_dp/n987 , \fpu_div_frac_dp/n985 ,
         \fpu_div_frac_dp/n984 , \fpu_div_frac_dp/n983 ,
         \fpu_div_frac_dp/n982 , \fpu_div_frac_dp/n981 ,
         \fpu_div_frac_dp/n980 , \fpu_div_frac_dp/n978 ,
         \fpu_div_frac_dp/n968 , \fpu_div_frac_dp/n967 ,
         \fpu_div_frac_dp/n960 , \fpu_div_frac_dp/n168 ,
         \fpu_div_frac_dp/n1439 , \fpu_div_frac_dp/n1438 ,
         \fpu_div_frac_dp/n1437 , \fpu_div_frac_dp/n1436 ,
         \fpu_div_frac_dp/n1435 , \fpu_div_frac_dp/n1434 ,
         \fpu_div_frac_dp/n1433 , \fpu_div_frac_dp/n1432 ,
         \fpu_div_frac_dp/n1431 , \fpu_div_frac_dp/n1430 ,
         \fpu_div_frac_dp/n1429 , \fpu_div_frac_dp/n1428 ,
         \fpu_div_frac_dp/n1427 , \fpu_div_frac_dp/n1426 ,
         \fpu_div_frac_dp/n1425 , \fpu_div_frac_dp/n1424 ,
         \fpu_div_frac_dp/n1423 , \fpu_div_frac_dp/n1422 ,
         \fpu_div_frac_dp/n1421 , \fpu_div_frac_dp/n1420 ,
         \fpu_div_frac_dp/n1419 , \fpu_div_frac_dp/n1418 ,
         \fpu_div_frac_dp/n1417 , \fpu_div_frac_dp/n1416 ,
         \fpu_div_frac_dp/n1415 , \fpu_div_frac_dp/n1414 ,
         \fpu_div_frac_dp/n1413 , \fpu_div_frac_dp/n1412 ,
         \fpu_div_frac_dp/n1411 , \fpu_div_frac_dp/n1410 ,
         \fpu_div_frac_dp/n1409 , \fpu_div_frac_dp/n1408 ,
         \fpu_div_frac_dp/n1407 , \fpu_div_frac_dp/n1406 ,
         \fpu_div_frac_dp/n1405 , \fpu_div_frac_dp/n1404 ,
         \fpu_div_frac_dp/n1403 , \fpu_div_frac_dp/n1402 ,
         \fpu_div_frac_dp/n1401 , \fpu_div_frac_dp/n1400 ,
         \fpu_div_frac_dp/n1399 , \fpu_div_frac_dp/n1398 ,
         \fpu_div_frac_dp/n1397 , \fpu_div_frac_dp/n1396 ,
         \fpu_div_frac_dp/n1395 , \fpu_div_frac_dp/n1394 ,
         \fpu_div_frac_dp/n1393 , \fpu_div_frac_dp/n1392 ,
         \fpu_div_frac_dp/n1391 , \fpu_div_frac_dp/n1390 ,
         \fpu_div_frac_dp/n1389 , \fpu_div_frac_dp/n1388 ,
         \fpu_div_frac_dp/n1387 , \fpu_div_frac_dp/n1386 ,
         \fpu_div_frac_dp/n1385 , \fpu_div_frac_dp/n1384 ,
         \fpu_div_frac_dp/n1383 , \fpu_div_frac_dp/n1382 ,
         \fpu_div_frac_dp/n1381 , \fpu_div_frac_dp/n1380 ,
         \fpu_div_frac_dp/n1379 , \fpu_div_frac_dp/n1378 ,
         \fpu_div_frac_dp/n1377 , \fpu_div_frac_dp/n1376 ,
         \fpu_div_frac_dp/n1375 , \fpu_div_frac_dp/n1374 ,
         \fpu_div_frac_dp/n1373 , \fpu_div_frac_dp/n1372 ,
         \fpu_div_frac_dp/n1371 , \fpu_div_frac_dp/n1370 ,
         \fpu_div_frac_dp/n1369 , \fpu_div_frac_dp/n1368 ,
         \fpu_div_frac_dp/n1367 , \fpu_div_frac_dp/n1366 ,
         \fpu_div_frac_dp/n1365 , \fpu_div_frac_dp/n1364 ,
         \fpu_div_frac_dp/n1363 , \fpu_div_frac_dp/n1362 ,
         \fpu_div_frac_dp/n1361 , \fpu_div_frac_dp/n1360 ,
         \fpu_div_frac_dp/n1359 , \fpu_div_frac_dp/n1358 ,
         \fpu_div_frac_dp/n1357 , \fpu_div_frac_dp/n1356 ,
         \fpu_div_frac_dp/n1355 , \fpu_div_frac_dp/n1354 ,
         \fpu_div_frac_dp/n1353 , \fpu_div_frac_dp/n1352 ,
         \fpu_div_frac_dp/n1351 , \fpu_div_frac_dp/n1350 ,
         \fpu_div_frac_dp/n1349 , \fpu_div_frac_dp/n1348 ,
         \fpu_div_frac_dp/n1347 , \fpu_div_frac_dp/n1346 ,
         \fpu_div_frac_dp/n1345 , \fpu_div_frac_dp/n1344 ,
         \fpu_div_frac_dp/n1343 , \fpu_div_frac_dp/n1342 ,
         \fpu_div_frac_dp/n1341 , \fpu_div_frac_dp/n1340 ,
         \fpu_div_frac_dp/n1339 , \fpu_div_frac_dp/n1338 ,
         \fpu_div_frac_dp/n1337 , \fpu_div_frac_dp/n1336 ,
         \fpu_div_frac_dp/n1335 , \fpu_div_frac_dp/n1334 ,
         \fpu_div_frac_dp/n1333 , \fpu_div_frac_dp/n1332 ,
         \fpu_div_frac_dp/n1331 , \fpu_div_frac_dp/n1330 ,
         \fpu_div_frac_dp/n1329 , \fpu_div_frac_dp/n1328 ,
         \fpu_div_frac_dp/n1327 , \fpu_div_frac_dp/n1326 ,
         \fpu_div_frac_dp/n1325 , \fpu_div_frac_dp/n1324 ,
         \fpu_div_frac_dp/n1323 , \fpu_div_frac_dp/n1322 ,
         \fpu_div_frac_dp/n1321 , \fpu_div_frac_dp/n1320 ,
         \fpu_div_frac_dp/n1319 , \fpu_div_frac_dp/n1318 ,
         \fpu_div_frac_dp/n1317 , \fpu_div_frac_dp/n1316 ,
         \fpu_div_frac_dp/n1315 , \fpu_div_frac_dp/n1314 ,
         \fpu_div_frac_dp/n1313 , \fpu_div_frac_dp/n1312 ,
         \fpu_div_frac_dp/n1311 , \fpu_div_frac_dp/n1310 ,
         \fpu_div_frac_dp/n1309 , \fpu_div_frac_dp/n1308 ,
         \fpu_div_frac_dp/n1307 , \fpu_div_frac_dp/n1306 ,
         \fpu_div_frac_dp/n1305 , \fpu_div_frac_dp/n1304 ,
         \fpu_div_frac_dp/n1303 , \fpu_div_frac_dp/n1302 ,
         \fpu_div_frac_dp/n1301 , \fpu_div_frac_dp/n1300 ,
         \fpu_div_frac_dp/n1299 , \fpu_div_frac_dp/n1298 ,
         \fpu_div_frac_dp/n1297 , \fpu_div_frac_dp/n1296 ,
         \fpu_div_frac_dp/n1295 , \fpu_div_frac_dp/n1294 ,
         \fpu_div_frac_dp/n1293 , \fpu_div_frac_dp/n1292 ,
         \fpu_div_frac_dp/n1291 , \fpu_div_frac_dp/n1290 ,
         \fpu_div_frac_dp/n1289 , \fpu_div_frac_dp/n1288 ,
         \fpu_div_frac_dp/n1287 , \fpu_div_frac_dp/n1286 ,
         \fpu_div_frac_dp/n1285 , \fpu_div_frac_dp/n1284 ,
         \fpu_div_frac_dp/n1283 , \fpu_div_frac_dp/n1282 ,
         \fpu_div_frac_dp/n1281 , \fpu_div_frac_dp/n1280 ,
         \fpu_div_frac_dp/n1279 , \fpu_div_frac_dp/n1278 ,
         \fpu_div_frac_dp/n1277 , \fpu_div_frac_dp/n1275 ,
         \fpu_div_frac_dp/n1274 , \fpu_div_frac_dp/n1273 ,
         \fpu_div_frac_dp/n1272 , \fpu_div_frac_dp/n1271 ,
         \fpu_div_frac_dp/n1270 , \fpu_div_frac_dp/n1269 ,
         \fpu_div_frac_dp/n1268 , \fpu_div_frac_dp/n1267 ,
         \fpu_div_frac_dp/n1266 , \fpu_div_frac_dp/n1265 ,
         \fpu_div_frac_dp/n1264 , \fpu_div_frac_dp/n1263 ,
         \fpu_div_frac_dp/n1262 , \fpu_div_frac_dp/n1261 ,
         \fpu_div_frac_dp/n1260 , \fpu_div_frac_dp/n1259 ,
         \fpu_div_frac_dp/n1258 , \fpu_div_frac_dp/n1257 ,
         \fpu_div_frac_dp/n1256 , \fpu_div_frac_dp/n1255 ,
         \fpu_div_frac_dp/n1254 , \fpu_div_frac_dp/n1253 ,
         \fpu_div_frac_dp/n1252 , \fpu_div_frac_dp/n1251 ,
         \fpu_div_frac_dp/n1250 , \fpu_div_frac_dp/n1249 ,
         \fpu_div_frac_dp/n1248 , \fpu_div_frac_dp/n1247 ,
         \fpu_div_frac_dp/n1246 , \fpu_div_frac_dp/n1245 ,
         \fpu_div_frac_dp/n1244 , \fpu_div_frac_dp/n1243 ,
         \fpu_div_frac_dp/n1242 , \fpu_div_frac_dp/n1241 ,
         \fpu_div_frac_dp/n1240 , \fpu_div_frac_dp/n1239 ,
         \fpu_div_frac_dp/n1238 , \fpu_div_frac_dp/n1237 ,
         \fpu_div_frac_dp/n1236 , \fpu_div_frac_dp/n1235 ,
         \fpu_div_frac_dp/n1234 , \fpu_div_frac_dp/n1233 ,
         \fpu_div_frac_dp/n1232 , \fpu_div_frac_dp/n1231 ,
         \fpu_div_frac_dp/n1230 , \fpu_div_frac_dp/n1229 ,
         \fpu_div_frac_dp/n1228 , \fpu_div_frac_dp/n1227 ,
         \fpu_div_frac_dp/n1226 , \fpu_div_frac_dp/n1225 ,
         \fpu_div_frac_dp/n1224 , \fpu_div_frac_dp/n1223 ,
         \fpu_div_frac_dp/n1222 , \fpu_div_frac_dp/n1221 ,
         \fpu_div_frac_dp/n1220 , \fpu_div_frac_dp/n1219 ,
         \fpu_div_frac_dp/n1218 , \fpu_div_frac_dp/n1217 ,
         \fpu_div_frac_dp/n1216 , \fpu_div_frac_dp/n1215 ,
         \fpu_div_frac_dp/n1214 , \fpu_div_frac_dp/n1213 ,
         \fpu_div_frac_dp/n1212 , \fpu_div_frac_dp/n1211 ,
         \fpu_div_frac_dp/n1210 , \fpu_div_frac_dp/n1209 ,
         \fpu_div_frac_dp/n1208 , \fpu_div_frac_dp/n1207 ,
         \fpu_div_frac_dp/n1206 , \fpu_div_frac_dp/n1205 ,
         \fpu_div_frac_dp/n1204 , \fpu_div_frac_dp/n1203 ,
         \fpu_div_frac_dp/n1202 , \fpu_div_frac_dp/n1201 ,
         \fpu_div_frac_dp/n1200 , \fpu_div_frac_dp/n1199 ,
         \fpu_div_frac_dp/n1198 , \fpu_div_frac_dp/n1197 ,
         \fpu_div_frac_dp/n1196 , \fpu_div_frac_dp/n1195 ,
         \fpu_div_frac_dp/n1194 , \fpu_div_frac_dp/n1193 ,
         \fpu_div_frac_dp/n1192 , \fpu_div_frac_dp/n1191 ,
         \fpu_div_frac_dp/n1190 , \fpu_div_frac_dp/n1189 ,
         \fpu_div_frac_dp/n1188 , \fpu_div_frac_dp/n1187 ,
         \fpu_div_frac_dp/n1186 , \fpu_div_frac_dp/n1185 ,
         \fpu_div_frac_dp/n1184 , \fpu_div_frac_dp/n1183 ,
         \fpu_div_frac_dp/n1182 , \fpu_div_frac_dp/n1181 ,
         \fpu_div_frac_dp/n1180 , \fpu_div_frac_dp/n1179 ,
         \fpu_div_frac_dp/n1178 , \fpu_div_frac_dp/n1177 ,
         \fpu_div_frac_dp/n1176 , \fpu_div_frac_dp/n1175 ,
         \fpu_div_frac_dp/n1174 , \fpu_div_frac_dp/n1173 ,
         \fpu_div_frac_dp/n1172 , \fpu_div_frac_dp/n1171 ,
         \fpu_div_frac_dp/n1170 , \fpu_div_frac_dp/n1169 ,
         \fpu_div_frac_dp/n1168 , \fpu_div_frac_dp/n1167 ,
         \fpu_div_frac_dp/n1166 , \fpu_div_frac_dp/n1165 ,
         \fpu_div_frac_dp/n1164 , \fpu_div_frac_dp/n1163 ,
         \fpu_div_frac_dp/n1162 , \fpu_div_frac_dp/n1161 ,
         \fpu_div_frac_dp/n1160 , \fpu_div_frac_dp/n1159 ,
         \fpu_div_frac_dp/n1158 , \fpu_div_frac_dp/n1157 ,
         \fpu_div_frac_dp/n1156 , \fpu_div_frac_dp/n1155 ,
         \fpu_div_frac_dp/n1154 , \fpu_div_frac_dp/n1153 ,
         \fpu_div_frac_dp/n1152 , \fpu_div_frac_dp/n1151 ,
         \fpu_div_frac_dp/n1150 , \fpu_div_frac_dp/n1149 ,
         \fpu_div_frac_dp/n1148 , \fpu_div_frac_dp/n1147 ,
         \fpu_div_frac_dp/n1146 , \fpu_div_frac_dp/n1145 ,
         \fpu_div_frac_dp/n1144 , \fpu_div_frac_dp/n1143 ,
         \fpu_div_frac_dp/n1142 , \fpu_div_frac_dp/n1141 ,
         \fpu_div_frac_dp/n1140 , \fpu_div_frac_dp/n1139 ,
         \fpu_div_frac_dp/n1138 , \fpu_div_frac_dp/n1137 ,
         \fpu_div_frac_dp/n1136 , \fpu_div_frac_dp/n1135 ,
         \fpu_div_frac_dp/n1134 , \fpu_div_frac_dp/n1133 ,
         \fpu_div_frac_dp/n1132 , \fpu_div_frac_dp/n1131 ,
         \fpu_div_frac_dp/n1130 , \fpu_div_frac_dp/n1129 ,
         \fpu_div_frac_dp/n1128 , \fpu_div_frac_dp/n1127 ,
         \fpu_div_frac_dp/n1126 , \fpu_div_frac_dp/n1125 ,
         \fpu_div_frac_dp/n1124 , \fpu_div_frac_dp/n1123 ,
         \fpu_div_frac_dp/n1122 , \fpu_div_frac_dp/n1121 ,
         \fpu_div_frac_dp/n1120 , \fpu_div_frac_dp/n1119 ,
         \fpu_div_frac_dp/n1118 , \fpu_div_frac_dp/n1117 ,
         \fpu_div_frac_dp/n1116 , \fpu_div_frac_dp/n1115 ,
         \fpu_div_frac_dp/n1114 , \fpu_div_frac_dp/n1113 ,
         \fpu_div_frac_dp/n1112 , \fpu_div_frac_dp/n1111 ,
         \fpu_div_frac_dp/n1110 , \fpu_div_frac_dp/n1109 ,
         \fpu_div_frac_dp/n1108 , \fpu_div_frac_dp/n1107 ,
         \fpu_div_frac_dp/n1106 , \fpu_div_frac_dp/n1105 ,
         \fpu_div_frac_dp/n1104 , \fpu_div_frac_dp/n1103 ,
         \fpu_div_frac_dp/n1102 , \fpu_div_frac_dp/n1101 ,
         \fpu_div_frac_dp/n1100 , \fpu_div_frac_dp/n1099 ,
         \fpu_div_frac_dp/n1098 , \fpu_div_frac_dp/n1097 ,
         \fpu_div_frac_dp/n1096 , \fpu_div_frac_dp/n1095 ,
         \fpu_div_frac_dp/n1094 , \fpu_div_frac_dp/n1093 ,
         \fpu_div_frac_dp/n1092 , \fpu_div_frac_dp/n1091 ,
         \fpu_div_frac_dp/n1090 , \fpu_div_frac_dp/n1089 ,
         \fpu_div_frac_dp/n1088 , \fpu_div_frac_dp/n1087 ,
         \fpu_div_frac_dp/n1086 , \fpu_div_frac_dp/n1085 ,
         \fpu_div_frac_dp/n1084 , \fpu_div_frac_dp/n1083 ,
         \fpu_div_frac_dp/n1082 , \fpu_div_frac_dp/n1081 ,
         \fpu_div_frac_dp/n1080 , \fpu_div_frac_dp/n1079 ,
         \fpu_div_frac_dp/n1078 , \fpu_div_frac_dp/n1077 ,
         \fpu_div_frac_dp/n1076 , \fpu_div_frac_dp/n1075 ,
         \fpu_div_frac_dp/n1074 , \fpu_div_frac_dp/n1073 ,
         \fpu_div_frac_dp/n1072 , \fpu_div_frac_dp/n1071 ,
         \fpu_div_frac_dp/n1070 , \fpu_div_frac_dp/n1069 ,
         \fpu_div_frac_dp/n1068 , \fpu_div_frac_dp/n1067 ,
         \fpu_div_frac_dp/n1066 , \fpu_div_frac_dp/n1065 ,
         \fpu_div_frac_dp/n1064 , \fpu_div_frac_dp/n1063 ,
         \fpu_div_frac_dp/n1062 , \fpu_div_frac_dp/n1061 ,
         \fpu_div_frac_dp/n1060 , \fpu_div_frac_dp/n1059 ,
         \fpu_div_frac_dp/n1058 , \fpu_div_frac_dp/n1057 ,
         \fpu_div_frac_dp/n1056 , \fpu_div_frac_dp/n487 ,
         \fpu_div_frac_dp/n486 , \fpu_div_frac_dp/n485 ,
         \fpu_div_frac_dp/n484 , \fpu_div_frac_dp/n483 ,
         \fpu_div_frac_dp/n482 , \fpu_div_frac_dp/n481 ,
         \fpu_div_frac_dp/n480 , \fpu_div_frac_dp/n479 ,
         \fpu_div_frac_dp/n478 , \fpu_div_frac_dp/n477 ,
         \fpu_div_frac_dp/n476 , \fpu_div_frac_dp/n475 ,
         \fpu_div_frac_dp/n474 , \fpu_div_frac_dp/n473 ,
         \fpu_div_frac_dp/n472 , \fpu_div_frac_dp/n471 ,
         \fpu_div_frac_dp/n470 , \fpu_div_frac_dp/n469 ,
         \fpu_div_frac_dp/n468 , \fpu_div_frac_dp/n467 ,
         \fpu_div_frac_dp/n466 , \fpu_div_frac_dp/n465 ,
         \fpu_div_frac_dp/n464 , \fpu_div_frac_dp/n463 ,
         \fpu_div_frac_dp/n462 , \fpu_div_frac_dp/n461 ,
         \fpu_div_frac_dp/n460 , \fpu_div_frac_dp/n459 ,
         \fpu_div_frac_dp/n458 , \fpu_div_frac_dp/n457 ,
         \fpu_div_frac_dp/n456 , \fpu_div_frac_dp/n455 ,
         \fpu_div_frac_dp/n454 , \fpu_div_frac_dp/n453 ,
         \fpu_div_frac_dp/n452 , \fpu_div_frac_dp/n451 ,
         \fpu_div_frac_dp/n450 , \fpu_div_frac_dp/n449 ,
         \fpu_div_frac_dp/n448 , \fpu_div_frac_dp/n447 ,
         \fpu_div_frac_dp/n446 , \fpu_div_frac_dp/n445 ,
         \fpu_div_frac_dp/n444 , \fpu_div_frac_dp/n443 ,
         \fpu_div_frac_dp/n442 , \fpu_div_frac_dp/n441 ,
         \fpu_div_frac_dp/n440 , \fpu_div_frac_dp/n439 ,
         \fpu_div_frac_dp/n438 , \fpu_div_frac_dp/n437 ,
         \fpu_div_frac_dp/n436 , \fpu_div_frac_dp/n435 ,
         \fpu_div_frac_dp/n434 , \fpu_div_frac_dp/n433 ,
         \fpu_div_frac_dp/n432 , \fpu_div_frac_dp/n431 ,
         \fpu_div_frac_dp/n430 , \fpu_div_frac_dp/n429 ,
         \fpu_div_frac_dp/n428 , \fpu_div_frac_dp/n427 ,
         \fpu_div_frac_dp/n426 , \fpu_div_frac_dp/n425 ,
         \fpu_div_frac_dp/n424 , \fpu_div_frac_dp/n422 ,
         \fpu_div_frac_dp/n421 , \fpu_div_frac_dp/n420 ,
         \fpu_div_frac_dp/n419 , \fpu_div_frac_dp/n418 ,
         \fpu_div_frac_dp/n417 , \fpu_div_frac_dp/n416 ,
         \fpu_div_frac_dp/n415 , \fpu_div_frac_dp/n414 ,
         \fpu_div_frac_dp/n413 , \fpu_div_frac_dp/n412 ,
         \fpu_div_frac_dp/n411 , \fpu_div_frac_dp/n410 ,
         \fpu_div_frac_dp/n409 , \fpu_div_frac_dp/n408 ,
         \fpu_div_frac_dp/n407 , \fpu_div_frac_dp/n406 ,
         \fpu_div_frac_dp/n405 , \fpu_div_frac_dp/n404 ,
         \fpu_div_frac_dp/n403 , \fpu_div_frac_dp/n402 ,
         \fpu_div_frac_dp/n401 , \fpu_div_frac_dp/n400 ,
         \fpu_div_frac_dp/n399 , \fpu_div_frac_dp/n398 ,
         \fpu_div_frac_dp/n397 , \fpu_div_frac_dp/n396 ,
         \fpu_div_frac_dp/n395 , \fpu_div_frac_dp/n394 ,
         \fpu_div_frac_dp/n393 , \fpu_div_frac_dp/n392 ,
         \fpu_div_frac_dp/n391 , \fpu_div_frac_dp/n390 ,
         \fpu_div_frac_dp/n389 , \fpu_div_frac_dp/n388 ,
         \fpu_div_frac_dp/n387 , \fpu_div_frac_dp/n386 ,
         \fpu_div_frac_dp/n385 , \fpu_div_frac_dp/n384 ,
         \fpu_div_frac_dp/n383 , \fpu_div_frac_dp/n382 ,
         \fpu_div_frac_dp/n381 , \fpu_div_frac_dp/n380 ,
         \fpu_div_frac_dp/n379 , \fpu_div_frac_dp/n378 ,
         \fpu_div_frac_dp/n377 , \fpu_div_frac_dp/n374 ,
         \fpu_div_frac_dp/n373 , \fpu_div_frac_dp/n372 ,
         \fpu_div_frac_dp/n371 , \fpu_div_frac_dp/n368 ,
         \fpu_div_frac_dp/n367 , \fpu_div_frac_dp/n366 ,
         \fpu_div_frac_dp/n364 , \fpu_div_frac_dp/n363 ,
         \fpu_div_frac_dp/n362 , \fpu_div_frac_dp/n361 ,
         \fpu_div_frac_dp/n360 , \fpu_div_frac_dp/n359 ,
         \fpu_div_frac_dp/n358 , \fpu_div_frac_dp/n354 ,
         \fpu_div_frac_dp/n350 , \fpu_div_frac_dp/n349 ,
         \fpu_div_frac_dp/n347 , \fpu_div_frac_dp/n345 ,
         \fpu_div_frac_dp/n344 , \fpu_div_frac_dp/n343 ,
         \fpu_div_frac_dp/n326 , \fpu_div_frac_dp/n325 ,
         \fpu_div_frac_dp/n324 , \fpu_div_frac_dp/n214 ,
         \fpu_div_frac_dp/n213 , \fpu_div_frac_dp/n212 ,
         \fpu_div_frac_dp/n211 , \fpu_div_frac_dp/n210 ,
         \fpu_div_frac_dp/n209 , \fpu_div_frac_dp/n208 ,
         \fpu_div_frac_dp/n207 , \fpu_div_frac_dp/n206 ,
         \fpu_div_frac_dp/n205 , \fpu_div_frac_dp/n204 ,
         \fpu_div_frac_dp/n203 , \fpu_div_frac_dp/n202 ,
         \fpu_div_frac_dp/n201 , \fpu_div_frac_dp/n200 ,
         \fpu_div_frac_dp/n199 , \fpu_div_frac_dp/n198 ,
         \fpu_div_frac_dp/n197 , \fpu_div_frac_dp/n196 ,
         \fpu_div_frac_dp/n195 , \fpu_div_frac_dp/n194 ,
         \fpu_div_frac_dp/n193 , \fpu_div_frac_dp/n192 ,
         \fpu_div_frac_dp/n191 , \fpu_div_frac_dp/n189 ,
         \fpu_div_frac_dp/n166 , \fpu_div_frac_dp/n165 ,
         \fpu_div_frac_dp/n164 , \fpu_div_frac_dp/n163 ,
         \fpu_div_frac_dp/n162 , \fpu_div_frac_dp/n160 ,
         \fpu_div_frac_dp/n158 , \fpu_div_frac_dp/n154 ,
         \fpu_div_frac_dp/n151 , \fpu_div_frac_dp/n148 ,
         \fpu_div_frac_dp/n147 , \fpu_div_frac_dp/n145 ,
         \fpu_div_frac_dp/n144 , \fpu_div_frac_dp/n142 ,
         \fpu_div_frac_dp/n141 , \fpu_div_frac_dp/n139 ,
         \fpu_div_frac_dp/n138 , \fpu_div_frac_dp/n136 ,
         \fpu_div_frac_dp/n135 , \fpu_div_frac_dp/n133 ,
         \fpu_div_frac_dp/n132 , \fpu_div_frac_dp/n130 ,
         \fpu_div_frac_dp/n129 , \fpu_div_frac_dp/n127 ,
         \fpu_div_frac_dp/n126 , \fpu_div_frac_dp/n124 ,
         \fpu_div_frac_dp/n123 , \fpu_div_frac_dp/n121 ,
         \fpu_div_frac_dp/n120 , \fpu_div_frac_dp/n118 ,
         \fpu_div_frac_dp/n117 , \fpu_div_frac_dp/n115 ,
         \fpu_div_frac_dp/n114 , \fpu_div_frac_dp/n112 ,
         \fpu_div_frac_dp/n111 , \fpu_div_frac_dp/n109 ,
         \fpu_div_frac_dp/n108 , \fpu_div_frac_dp/n106 ,
         \fpu_div_frac_dp/n105 , \fpu_div_frac_dp/n103 ,
         \fpu_div_frac_dp/n102 , \fpu_div_frac_dp/n100 , \fpu_div_frac_dp/n99 ,
         \fpu_div_frac_dp/n96 , \fpu_div_frac_dp/n94 , \fpu_div_frac_dp/n93 ,
         \fpu_div_frac_dp/n92 , \fpu_div_frac_dp/n83 , \fpu_div_frac_dp/n79 ,
         \fpu_div_frac_dp/n76 , \fpu_div_frac_dp/n64 , \fpu_div_frac_dp/n61 ,
         \fpu_div_frac_dp/n58 , \fpu_div_frac_dp/n43 , \fpu_div_frac_dp/n40 ,
         \fpu_div_frac_dp/n20 , \fpu_div_frac_dp/n19 , \fpu_div_frac_dp/n17 ,
         \fpu_div_frac_dp/n16 , \fpu_div_frac_dp/n14 , \fpu_div_frac_dp/n13 ,
         \fpu_div_frac_dp/n11 , \fpu_div_frac_dp/n10 , \fpu_div_frac_dp/n8 ,
         \fpu_div_frac_dp/n6 , \fpu_div_frac_dp/n4 , \fpu_div_frac_dp/n1 ,
         \fpu_div_frac_dp/i_div_shl_data/N3 ,
         \fpu_div_frac_dp/i_div_shl_data/N4 ,
         \fpu_div_frac_dp/i_div_shl_data/N5 ,
         \fpu_div_frac_dp/i_div_shl_data/N6 ,
         \fpu_div_frac_dp/i_div_shl_data/N7 ,
         \fpu_div_frac_dp/i_div_shl_data/N8 ,
         \fpu_div_frac_dp/i_div_shl_data/N9 ,
         \fpu_div_frac_dp/i_div_shl_data/N10 ,
         \fpu_div_frac_dp/i_div_shl_data/N11 ,
         \fpu_div_frac_dp/i_div_shl_data/N12 ,
         \fpu_div_frac_dp/i_div_shl_data/N13 ,
         \fpu_div_frac_dp/i_div_shl_data/N14 ,
         \fpu_div_frac_dp/i_div_shl_data/N15 ,
         \fpu_div_frac_dp/i_div_shl_data/N16 ,
         \fpu_div_frac_dp/i_div_shl_data/N17 ,
         \fpu_div_frac_dp/i_div_shl_data/N18 ,
         \fpu_div_frac_dp/i_div_shl_data/N19 ,
         \fpu_div_frac_dp/i_div_shl_data/N20 ,
         \fpu_div_frac_dp/i_div_shl_data/N21 ,
         \fpu_div_frac_dp/i_div_shl_data/N22 ,
         \fpu_div_frac_dp/i_div_shl_data/N23 ,
         \fpu_div_frac_dp/i_div_shl_data/N24 ,
         \fpu_div_frac_dp/i_div_shl_data/N25 ,
         \fpu_div_frac_dp/i_div_shl_data/N26 ,
         \fpu_div_frac_dp/i_div_shl_data/N27 ,
         \fpu_div_frac_dp/i_div_shl_data/N28 ,
         \fpu_div_frac_dp/i_div_shl_data/N29 ,
         \fpu_div_frac_dp/i_div_shl_data/N31 ,
         \fpu_div_frac_dp/i_div_shl_data/N32 ,
         \fpu_div_frac_dp/i_div_shl_data/N33 ,
         \fpu_div_frac_dp/i_div_shl_data/N34 ,
         \fpu_div_frac_dp/i_div_shl_data/N35 ,
         \fpu_div_frac_dp/i_div_shl_data/N36 ,
         \fpu_div_frac_dp/i_div_shl_data/N37 ,
         \fpu_div_frac_dp/i_div_shl_data/N38 ,
         \fpu_div_frac_dp/i_div_shl_data/N39 ,
         \fpu_div_frac_dp/i_div_shl_data/N40 ,
         \fpu_div_frac_dp/i_div_shl_data/N41 ,
         \fpu_div_frac_dp/i_div_shl_data/N42 ,
         \fpu_div_frac_dp/i_div_shl_data/N43 ,
         \fpu_div_frac_dp/i_div_shl_data/N44 ,
         \fpu_div_frac_dp/i_div_shl_data/N45 ,
         \fpu_div_frac_dp/i_div_shl_data/N46 ,
         \fpu_div_frac_dp/i_div_shl_data/N47 ,
         \fpu_div_frac_dp/i_div_shl_data/N48 ,
         \fpu_div_frac_dp/i_div_shl_data/N49 ,
         \fpu_div_frac_dp/i_div_shl_data/N50 ,
         \fpu_div_frac_dp/i_div_shl_data/N51 ,
         \fpu_div_frac_dp/i_div_shl_data/N52 ,
         \fpu_div_frac_dp/i_div_shl_data/N53 ,
         \fpu_div_frac_dp/i_div_shl_data/N54 ,
         \fpu_div_frac_dp/i_div_shl_data/N55 ,
         \fpu_div_frac_dp/i_dstg_xtra_regs/N4 ,
         \fpu_div_frac_dp/i_dstg_xtra_regs/N5 ,
         \fpu_div_frac_dp/i_dstg_xtra_regs/N6 ,
         \fpu_div_frac_dp/i_dstg_xtra_regs/N7 ,
         \fpu_div_frac_dp/i_dstg_xtra_regs/N9 ,
         \fpu_div_frac_dp/i_div_norm_inv/N3 ,
         \fpu_div_frac_dp/i_div_norm_inv/N4 ,
         \fpu_div_frac_dp/i_div_norm_inv/N5 ,
         \fpu_div_frac_dp/i_div_norm_inv/N6 ,
         \fpu_div_frac_dp/i_div_norm_inv/N7 ,
         \fpu_div_frac_dp/i_div_norm_inv/N8 ,
         \fpu_div_frac_dp/i_div_norm_inv/N9 ,
         \fpu_div_frac_dp/i_div_norm_inv/N10 ,
         \fpu_div_frac_dp/i_div_norm_inv/N11 ,
         \fpu_div_frac_dp/i_div_norm_inv/N12 ,
         \fpu_div_frac_dp/i_div_norm_inv/N13 ,
         \fpu_div_frac_dp/i_div_norm_inv/N14 ,
         \fpu_div_frac_dp/i_div_norm_inv/N15 ,
         \fpu_div_frac_dp/i_div_norm_inv/N16 ,
         \fpu_div_frac_dp/i_div_norm_inv/N17 ,
         \fpu_div_frac_dp/i_div_norm_inv/N18 ,
         \fpu_div_frac_dp/i_div_norm_inv/N19 ,
         \fpu_div_frac_dp/i_div_norm_inv/N20 ,
         \fpu_div_frac_dp/i_div_norm_inv/N21 ,
         \fpu_div_frac_dp/i_div_norm_inv/N22 ,
         \fpu_div_frac_dp/i_div_norm_inv/N23 ,
         \fpu_div_frac_dp/i_div_norm_inv/N24 ,
         \fpu_div_frac_dp/i_div_norm_inv/N25 ,
         \fpu_div_frac_dp/i_div_norm_inv/N26 ,
         \fpu_div_frac_dp/i_div_norm_inv/N27 ,
         \fpu_div_frac_dp/i_div_norm_inv/N28 ,
         \fpu_div_frac_dp/i_div_norm_inv/N29 ,
         \fpu_div_frac_dp/i_div_norm_inv/N30 ,
         \fpu_div_frac_dp/i_div_norm_inv/N31 ,
         \fpu_div_frac_dp/i_div_norm_inv/N32 ,
         \fpu_div_frac_dp/i_div_norm_inv/N33 ,
         \fpu_div_frac_dp/i_div_norm_inv/N34 ,
         \fpu_div_frac_dp/i_div_norm_inv/N35 ,
         \fpu_div_frac_dp/i_div_norm_inv/N36 ,
         \fpu_div_frac_dp/i_div_norm_inv/N37 ,
         \fpu_div_frac_dp/i_div_norm_inv/N38 ,
         \fpu_div_frac_dp/i_div_norm_inv/N39 ,
         \fpu_div_frac_dp/i_div_norm_inv/N40 ,
         \fpu_div_frac_dp/i_div_norm_inv/N41 ,
         \fpu_div_frac_dp/i_div_norm_inv/N42 ,
         \fpu_div_frac_dp/i_div_norm_inv/N43 ,
         \fpu_div_frac_dp/i_div_norm_inv/N44 ,
         \fpu_div_frac_dp/i_div_norm_inv/N45 ,
         \fpu_div_frac_dp/i_div_norm_inv/N46 ,
         \fpu_div_frac_dp/i_div_norm_inv/N47 ,
         \fpu_div_frac_dp/i_div_norm_inv/N48 ,
         \fpu_div_frac_dp/i_div_norm_inv/N49 ,
         \fpu_div_frac_dp/i_div_norm_inv/N50 ,
         \fpu_div_frac_dp/i_div_norm_inv/N51 ,
         \fpu_div_frac_dp/i_div_norm_inv/N52 ,
         \fpu_div_frac_dp/i_div_norm_inv/N53 ,
         \fpu_div_frac_dp/i_div_norm_inv/N54 ,
         \fpu_div_frac_dp/i_div_norm_inv/N55 ,
         \fpu_div_frac_dp/ckbuf_div_frac_dp/N1 ,
         \fpu_div_frac_dp/div_shl_data[52] ,
         \fpu_div_frac_dp/div_norm_inv[45] ,
         \fpu_div_frac_dp/div_norm_inv[43] ,
         \fpu_div_frac_dp/div_norm_inv[41] ,
         \fpu_div_frac_dp/div_norm_inv[37] ,
         \fpu_div_frac_dp/div_norm_inv[32] ,
         \fpu_div_frac_dp/div_norm_inv[26] ,
         \fpu_div_frac_dp/div_norm_inv[25] ,
         \fpu_div_frac_dp/div_norm_inv[23] ,
         \fpu_div_frac_dp/div_norm_inv[21] ,
         \fpu_div_frac_dp/div_norm_inv[14] ,
         \fpu_div_frac_dp/div_norm_inv[13] , \fpu_div_frac_dp/div_norm_inv[6] ,
         \fpu_div_frac_dp/div_norm_inv[5] , \fpu_div_frac_dp/div_norm_inv[0] ,
         \fpu_div_frac_dp/rclk , \fpu_div_frac_dp/d1stg_step , n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291;
  wire   [12:0] div_exp1;
  wire   [12:0] div_exp_out;
  assign div_exp_outa[10] = div_exp_out[10];
  assign div_exp_outa[9] = div_exp_out[9];
  assign div_exp_outa[8] = div_exp_out[8];
  assign div_exp_outa[7] = div_exp_out[7];
  assign div_exp_outa[6] = div_exp_out[6];
  assign div_exp_outa[5] = div_exp_out[5];
  assign div_exp_outa[4] = div_exp_out[4];
  assign div_exp_outa[3] = div_exp_out[3];
  assign div_exp_outa[2] = div_exp_out[2];
  assign div_exp_outa[1] = div_exp_out[1];
  assign div_exp_outa[0] = div_exp_out[0];
  assign so = 1'b0;
  assign d1stg_step = \fpu_div_frac_dp/d1stg_step ;

  DFFARX1 \fpu_div_ctl/dffrl_div_ctl/q_reg[0]  ( .D(
        \fpu_div_ctl/dffrl_div_ctl/N4 ), .CLK(rclk), .RSTB(arst_l), .Q(n1781), 
        .QN(n152) );
  LATCHX1 \fpu_div_exp_dp/ckbuf_div_exp_dp/clken_reg  ( .CLK(
        \fpu_div_frac_dp/rclk ), .D(\fpu_div_exp_dp/ckbuf_div_exp_dp/N1 ), .Q(
        \fpu_div_exp_dp/ckbuf_div_exp_dp/clken ), .QN(n151) );
  DFFX1 \fpu_div_exp_dp/i_div_exp1/q_reg[12]  ( .D(n514), .CLK(n577), .Q(n1782), .QN(n607) );
  DFFX1 \fpu_div_ctl/i_d5stg_opdec/q_reg[0]  ( .D(n485), .CLK(rclk), .Q(n1461), 
        .QN(n611) );
  DFFX1 \fpu_div_ctl/i_divd_cnt_lt_52a/q_reg[0]  ( .D(n513), .CLK(rclk), .Q(
        n1856), .QN(n150) );
  DFFX1 \fpu_div_ctl/i_d1stg_div/q_reg[0]  ( .D(\fpu_div_ctl/i_d1stg_div/N7 ), 
        .CLK(rclk), .Q(\fpu_div_ctl/d1stg_div ), .QN(n149) );
  DFFX1 \fpu_div_ctl/i_d1stg_op/q_reg[0]  ( .D(\fpu_div_ctl/i_d1stg_op/N14 ), 
        .CLK(rclk), .Q(n1785), .QN(n148) );
  DFFX1 \fpu_div_ctl/i_d1stg_op/q_reg[1]  ( .D(\fpu_div_ctl/i_d1stg_op/N15 ), 
        .CLK(rclk), .Q(n1784), .QN(n177) );
  DFFX1 \fpu_div_ctl/i_d1stg_op/q_reg[2]  ( .D(\fpu_div_ctl/i_d1stg_op/N16 ), 
        .CLK(rclk), .Q(\fpu_div_ctl/d1stg_op[2] ), .QN(n146) );
  DFFX1 \fpu_div_ctl/i_d1stg_op/q_reg[3]  ( .D(\fpu_div_ctl/i_d1stg_op/N17 ), 
        .CLK(rclk), .Q(\fpu_div_ctl/d1stg_op[3] ), .QN(n145) );
  DFFX1 \fpu_div_ctl/i_d1stg_op/q_reg[4]  ( .D(\fpu_div_ctl/i_d1stg_op/N18 ), 
        .CLK(rclk), .Q(\fpu_div_ctl/d1stg_op[4] ), .QN(n144) );
  DFFX1 \fpu_div_ctl/i_d1stg_op/q_reg[5]  ( .D(\fpu_div_ctl/i_d1stg_op/N19 ), 
        .CLK(rclk), .QN(n179) );
  DFFX1 \fpu_div_ctl/i_d1stg_op/q_reg[6]  ( .D(\fpu_div_ctl/i_d1stg_op/N20 ), 
        .CLK(rclk), .Q(\fpu_div_ctl/d1stg_op[6] ), .QN(n142) );
  DFFX1 \fpu_div_ctl/i_d1stg_op/q_reg[7]  ( .D(\fpu_div_ctl/i_d1stg_op/N21 ), 
        .CLK(rclk), .Q(\fpu_div_ctl/d1stg_op[7] ), .QN(n141) );
  DFFSSRX1 \fpu_div_ctl/i_d2stg_opdec/q_reg[1]  ( .D(n1354), .RSTB(n355), 
        .SETB(1'b1), .CLK(rclk), .Q(div_expadd1_in2_exp_in2_sng), .QN(n182) );
  DFFX1 \fpu_div_ctl/i_d3stg_opdec/q_reg[1]  ( .D(
        \fpu_div_ctl/i_d3stg_opdec/N10 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d3stg_opdec[1] ) );
  DFFSSRX1 \fpu_div_ctl/i_d4stg_opdec/q_reg[1]  ( .D(n1354), .RSTB(
        \fpu_div_ctl/d3stg_opdec[1] ), .SETB(1'b1), .CLK(rclk), .Q(n1851), 
        .QN(n138) );
  DFFX1 \fpu_div_ctl/i_d5stg_opdec/q_reg[1]  ( .D(n486), .CLK(rclk), .Q(n1396), 
        .QN(n581) );
  DFFX1 \fpu_div_ctl/i_d6stg_opdec/q_reg[1]  ( .D(
        \fpu_div_ctl/i_d6stg_opdec/N10 ), .CLK(rclk), .Q(d6stg_fdivs) );
  DFFSSRX1 \fpu_div_ctl/i_d7stg_opdec/q_reg[1]  ( .D(n1354), .RSTB(d6stg_fdivs), .SETB(1'b1), .CLK(rclk), .Q(n1391), .QN(n630) );
  DFFSSRX1 \fpu_div_ctl/i_d2stg_opdec/q_reg[0]  ( .D(n1354), .RSTB(n354), 
        .SETB(1'b1), .CLK(rclk), .Q(div_expadd1_in2_exp_in2_dbl), .QN(n181) );
  DFFX1 \fpu_div_ctl/i_d3stg_opdec/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d3stg_opdec/N9 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d3stg_opdec[0] ) );
  DFFSSRX1 \fpu_div_ctl/i_d4stg_opdec/q_reg[0]  ( .D(n1354), .RSTB(
        \fpu_div_ctl/d3stg_opdec[0] ), .SETB(1'b1), .CLK(rclk), .Q(n1852), 
        .QN(n131) );
  DFFX1 \fpu_div_ctl/i_d2stg_opdec/q_reg[2]  ( .D(
        \fpu_div_ctl/i_d2stg_opdec/N11 ), .CLK(rclk), .Q(n619), .QN(n1549) );
  DFFX1 \fpu_div_ctl/i_d3stg_opdec/q_reg[2]  ( .D(
        \fpu_div_ctl/i_d3stg_opdec/N11 ), .CLK(rclk), .Q(d3stg_fdiv), .QN(n184) );
  DFFX1 \fpu_div_ctl/i_d4stg_opdec/q_reg[2]  ( .D(
        \fpu_div_ctl/i_d4stg_opdec/N11 ), .CLK(rclk), .Q(n1433), .QN(n185) );
  DFFSSRX1 \fpu_div_ctl/i_d5stg_opdec/q_reg[2]  ( .D(n272), .RSTB(n185), 
        .SETB(n1354), .CLK(rclk), .Q(n191), .QN(n1373) );
  DFFX1 \fpu_div_ctl/i_d6stg_opdec/q_reg[2]  ( .D(
        \fpu_div_ctl/i_d6stg_opdec/N11 ), .CLK(rclk), .Q(n1552), .QN(n193) );
  DFFX1 \fpu_div_ctl/i_d7stg_opdec/q_reg[2]  ( .D(
        \fpu_div_ctl/i_d7stg_opdec/N11 ), .CLK(rclk), .Q(n1393), .QN(n194) );
  DFFSSRX1 \fpu_div_ctl/i_d8stg_opdec/q_reg[2]  ( .D(n939), .RSTB(n194), 
        .SETB(n1354), .CLK(rclk), .Q(n196) );
  DFFX1 \fpu_div_ctl/i_divd_cnt_lt_52/q_reg[0]  ( .D(n466), .CLK(rclk), .Q(
        n1857), .QN(n127) );
  DFFX1 \fpu_div_ctl/i_divs_cnt_lt_23a/q_reg[0]  ( .D(n467), .CLK(rclk), .Q(
        n1854), .QN(n126) );
  DFFX1 \fpu_div_ctl/i_divs_cnt_lt_23/q_reg[0]  ( .D(n468), .CLK(rclk), .Q(
        n1853), .QN(n125) );
  DFFX1 \fpu_div_ctl/i_d8stg_opdec/q_reg[1]  ( .D(n476), .CLK(rclk), .Q(
        d8stg_fdivs), .QN(n124) );
  DFFX1 \fpu_div_ctl/i_div_expadd2_in1_exp_out/q_reg[0]  ( .D(
        \fpu_div_ctl/i_div_expadd2_in1_exp_out/N7 ), .CLK(rclk), .Q(
        div_expadd2_in1_exp_out), .QN(n578) );
  DFFX1 \fpu_div_ctl/i_div_cnt/q_reg[5]  ( .D(n479), .CLK(rclk), .Q(n1545), 
        .QN(n620) );
  DFFX1 \fpu_div_ctl/i_div_cnt/q_reg[4]  ( .D(n480), .CLK(rclk), .Q(n1541), 
        .QN(n602) );
  DFFX1 \fpu_div_ctl/i_div_cnt/q_reg[3]  ( .D(n481), .CLK(rclk), .Q(n1395), 
        .QN(n586) );
  DFFX1 \fpu_div_ctl/i_div_cnt/q_reg[2]  ( .D(n482), .CLK(rclk), .Q(n1542), 
        .QN(n612) );
  DFFX1 \fpu_div_ctl/i_div_cnt/q_reg[1]  ( .D(n483), .CLK(rclk), .Q(n1372), 
        .QN(n594) );
  DFFX1 \fpu_div_ctl/i_div_cnt/q_reg[0]  ( .D(n484), .CLK(rclk), .Q(
        \fpu_div_ctl/div_cnt[0] ), .QN(n616) );
  DFFX1 \fpu_div_ctl/i_div_pipe_active/q_reg[0]  ( .D(
        \fpu_div_ctl/i_div_pipe_active/N7 ), .CLK(rclk), .Q(div_pipe_active)
         );
  DFFX1 \fpu_div_ctl/i_d234stg_fdiv/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d234stg_fdiv/N7 ), .CLK(rclk), .Q(d234stg_fdiv), .QN(
        n117) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[0]  ( .D(n413), .CLK(n577), .Q(
        n1725) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[1]  ( .D(n414), .CLK(n577), .Q(
        n1730) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[2]  ( .D(n415), .CLK(n577), .Q(
        n1724) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[3]  ( .D(n416), .CLK(n577), .Q(
        n623), .QN(n208) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[4]  ( .D(n417), .CLK(n577), .Q(
        n1532) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[5]  ( .D(n418), .CLK(n577), .Q(
        n622), .QN(n209) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[6]  ( .D(n419), .CLK(n577), .Q(
        n1534) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[7]  ( .D(n420), .CLK(n577), .Q(
        n1640) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[8]  ( .D(n421), .CLK(n577), .Q(
        n1642) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[9]  ( .D(n422), .CLK(n577), .Q(
        n1676) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in2/q_reg[10]  ( .D(n423), .CLK(n577), .Q(
        n1491) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[0]  ( .D(n424), .CLK(n577), .Q(
        n1872), .QN(n107) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[1]  ( .D(n425), .CLK(n577), .Q(
        n1876), .QN(n106) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[2]  ( .D(n426), .CLK(n577), .Q(
        n1871), .QN(n105) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[3]  ( .D(n427), .CLK(n577), .Q(
        n1855), .QN(n104) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[4]  ( .D(n428), .CLK(n577), .Q(
        n1860), .QN(n103) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[5]  ( .D(n429), .CLK(n577), .Q(
        n1863), .QN(n102) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[6]  ( .D(n430), .CLK(n577), .Q(
        n1862), .QN(n101) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[7]  ( .D(n431), .CLK(n577), .Q(
        n1861), .QN(n100) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[8]  ( .D(n432), .CLK(n577), .Q(
        n1858), .QN(n99) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[9]  ( .D(n433), .CLK(n577), .Q(
        n1865), .QN(n98) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_in1/q_reg[10]  ( .D(n434), .CLK(n577), .Q(
        n1859), .QN(n97) );
  DFFX1 \fpu_div_ctl/i_div_exp_in2_exp_neq_ffs/q_reg[0]  ( .D(n451), .CLK(rclk), .Q(n1647), .QN(n585) );
  DFFX1 \fpu_div_ctl/i_div_exp_in2_exp_eq_0/q_reg[0]  ( .D(n453), .CLK(rclk), 
        .Q(n606), .QN(n168) );
  DFFX1 \fpu_div_ctl/i_div_frac_in2_53_32_neq_0/q_reg[0]  ( .D(n454), .CLK(
        rclk), .Q(n1679), .QN(n1353) );
  DFFX1 \fpu_div_ctl/i_div_frac_in2_50_0_neq_0/q_reg[0]  ( .D(n455), .CLK(rclk), .Q(n1682), .QN(n96) );
  DFFX1 \fpu_div_ctl/i_div_frac_in2_53_0_neq_0/q_reg[0]  ( .D(n456), .CLK(rclk), .Q(n1869), .QN(n95) );
  DFFX1 \fpu_div_ctl/i_div_frac_in2_54/q_reg[0]  ( .D(n457), .CLK(rclk), .Q(
        n1645), .QN(n621) );
  DFFX1 \fpu_div_ctl/i_d2stg_zero_in2/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_zero_in2/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_zero_in2 ), .QN(n93) );
  DFFX1 \fpu_div_ctl/i_div_frac_in2_51/q_reg[0]  ( .D(n458), .CLK(rclk), .Q(
        n1651), .QN(n624) );
  DFFX1 \fpu_div_ctl/i_div_exp_in1_exp_neq_ffs/q_reg[0]  ( .D(n459), .CLK(rclk), .Q(n1543), .QN(n591) );
  DFFX1 \fpu_div_ctl/i_div_exp_in1_exp_eq_0/q_reg[0]  ( .D(n460), .CLK(rclk), 
        .Q(n604), .QN(n164) );
  DFFX1 \fpu_div_ctl/i_div_frac_in1_53_32_neq_0/q_reg[0]  ( .D(n461), .CLK(
        rclk), .Q(n1490), .QN(n90) );
  DFFX1 \fpu_div_ctl/i_div_frac_in1_50_0_neq_0/q_reg[0]  ( .D(n462), .CLK(rclk), .Q(n1489), .QN(n89) );
  DFFX1 \fpu_div_ctl/i_div_frac_in1_53_0_neq_0/q_reg[0]  ( .D(n463), .CLK(rclk), .Q(n1868), .QN(n88) );
  DFFX1 \fpu_div_ctl/i_div_frac_in1_54/q_reg[0]  ( .D(n464), .CLK(rclk), .Q(
        n1648), .QN(n627) );
  DFFSSRX1 \fpu_div_ctl/i_d2stg_zero_in/q_reg[0]  ( .D(n1356), .RSTB(n253), 
        .SETB(n1047), .CLK(rclk), .Q(n86), .QN(\fpu_div_ctl/d2stg_zero_in ) );
  DFFX1 \fpu_div_ctl/i_d2stg_2zero_in/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_2zero_in/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_2zero_in ) );
  DFFX1 \fpu_div_ctl/i_div_frac_in1_51/q_reg[0]  ( .D(n465), .CLK(rclk), .Q(
        n1672), .QN(n628) );
  DFFX1 \fpu_div_ctl/i_d1stg_id/q_reg[0]  ( .D(n495), .CLK(rclk), .Q(n1723) );
  DFFSSRX1 \fpu_div_ctl/i_div_id_out/q_reg[0]  ( .D(n1047), .RSTB(
        div_id_out_in[0]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_div_ctl/div_id_out[0] ) );
  DFFX1 \fpu_div_ctl/i_d1stg_id/q_reg[1]  ( .D(n496), .CLK(rclk), .Q(n1722) );
  DFFSSRX1 \fpu_div_ctl/i_div_id_out/q_reg[1]  ( .D(n1047), .RSTB(
        div_id_out_in[1]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_div_ctl/div_id_out[1] ) );
  DFFX1 \fpu_div_ctl/i_d1stg_id/q_reg[2]  ( .D(n497), .CLK(rclk), .Q(n1715), 
        .QN(n608) );
  DFFX1 \fpu_div_ctl/i_d1stg_id/q_reg[3]  ( .D(n498), .CLK(rclk), .Q(n1551), 
        .QN(n1351) );
  DFFX1 \fpu_div_ctl/i_d1stg_id/q_reg[4]  ( .D(n499), .CLK(rclk), .Q(n1786), 
        .QN(n597) );
  DFFSSRX1 \fpu_div_ctl/i_div_id_out/q_reg[5]  ( .D(n1047), .RSTB(
        div_id_out_in[5]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_div_ctl/div_id_out[5] ) );
  DFFSSRX1 \fpu_div_ctl/i_div_id_out/q_reg[4]  ( .D(n1047), .RSTB(
        div_id_out_in[4]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_div_ctl/div_id_out[4] ) );
  DFFSSRX1 \fpu_div_ctl/i_div_id_out/q_reg[3]  ( .D(n1047), .RSTB(
        div_id_out_in[3]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_div_ctl/div_id_out[3] ) );
  DFFSSRX1 \fpu_div_ctl/i_div_id_out/q_reg[2]  ( .D(n1047), .RSTB(
        div_id_out_in[2]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_div_ctl/div_id_out[2] ) );
  DFFSSRX1 \fpu_div_ctl/i_div_id_out/q_reg[9]  ( .D(n1047), .RSTB(
        div_id_out_in[9]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_div_ctl/div_id_out[9] ) );
  DFFSSRX1 \fpu_div_ctl/i_div_id_out/q_reg[8]  ( .D(n1047), .RSTB(
        div_id_out_in[8]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_div_ctl/div_id_out[8] ) );
  DFFSSRX1 \fpu_div_ctl/i_div_id_out/q_reg[7]  ( .D(n1047), .RSTB(
        div_id_out_in[7]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_div_ctl/div_id_out[7] ) );
  DFFSSRX1 \fpu_div_ctl/i_div_id_out/q_reg[6]  ( .D(n1047), .RSTB(
        div_id_out_in[6]), .SETB(1'b1), .CLK(rclk), .Q(
        \fpu_div_ctl/div_id_out[6] ) );
  DFFX1 \fpu_div_ctl/i_d1stg_rnd_mode/q_reg[0]  ( .D(n500), .CLK(rclk), .Q(
        n1732) );
  DFFX1 \fpu_div_ctl/i_div_rnd_mode/q_reg[0]  ( .D(n477), .CLK(rclk), .Q(n593), 
        .QN(n201) );
  DFFX1 \fpu_div_ctl/i_d1stg_rnd_mode/q_reg[1]  ( .D(n501), .CLK(rclk), .Q(
        n1875), .QN(n59) );
  DFFX1 \fpu_div_ctl/i_div_rnd_mode/q_reg[1]  ( .D(n478), .CLK(rclk), .Q(
        \fpu_div_ctl/div_rnd_mode[1] ), .QN(n58) );
  DFFX1 \fpu_div_ctl/i_d1stg_dblopa/q_reg[0]  ( .D(n502), .CLK(rclk), .Q(n1720), .QN(n520) );
  DFFX1 \fpu_div_ctl/i_d2stg_denorm_dbl_in2/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_denorm_dbl_in2/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_denorm_dbl_in2 ) );
  DFFX1 \fpu_div_ctl/i_d2stg_norm_dbl_in2/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_norm_dbl_in2/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_norm_dbl_in2 ) );
  DFFX1 \fpu_div_ctl/i_d1stg_dblopa/q_reg[1]  ( .D(n503), .CLK(rclk), .Q(n1375), .QN(n54) );
  DFFX1 \fpu_div_ctl/i_d1stg_dblopa/q_reg[2]  ( .D(n504), .CLK(rclk), .Q(n1547), .QN(n615) );
  DFFX1 \fpu_div_ctl/i_d1stg_dblopa/q_reg[3]  ( .D(n505), .CLK(rclk), .Q(n1731), .QN(n52) );
  DFFX1 \fpu_div_ctl/i_d1stg_dblopa/q_reg[4]  ( .D(n506), .CLK(rclk), .Q(
        \fpu_div_ctl/d1stg_dblopa[4] ) );
  DFFX1 \fpu_div_ctl/i_div_expadd1_in1_dbl/q_reg[0]  ( .D(
        \fpu_div_ctl/i_div_expadd1_in1_dbl/N3 ), .CLK(rclk), .Q(
        div_expadd1_in1_dbl), .QN(n587) );
  DFFX1 \fpu_div_ctl/i_d1stg_sngopa/q_reg[0]  ( .D(n508), .CLK(rclk), .Q(n1643), .QN(n50) );
  DFFX1 \fpu_div_ctl/i_d2stg_denorm_sng_in2/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_denorm_sng_in2/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_denorm_sng_in2 ) );
  DFFX1 \fpu_div_ctl/i_d2stg_norm_sng_in2/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_norm_sng_in2/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_norm_sng_in2 ) );
  DFFX1 \fpu_div_ctl/i_d1stg_sngopa/q_reg[1]  ( .D(n509), .CLK(rclk), .Q(n1376), .QN(n47) );
  DFFX1 \fpu_div_ctl/i_d2stg_snan_in1/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_snan_in1/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_snan_in1 ), .QN(n629) );
  DFFSSRX1 \fpu_div_ctl/i_d2stg_snan_in2/q_reg[0]  ( .D(n373), .RSTB(n370), 
        .SETB(n1047), .CLK(rclk), .Q(n1349), .QN(n1877) );
  DFFSSRX1 \fpu_div_ctl/i_d2stg_qnan_in2/q_reg[0]  ( .D(n351), .RSTB(n352), 
        .SETB(n1047), .CLK(rclk), .Q(n617), .QN(n1878) );
  DFFX1 \fpu_div_ctl/i_d2stg_qnan_in1/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_qnan_in1/N3 ), .CLK(rclk), .QN(n173) );
  DFFX1 \fpu_div_ctl/i_d1stg_sngopa/q_reg[2]  ( .D(n510), .CLK(rclk), .Q(n1401), .QN(n600) );
  DFFX1 \fpu_div_ctl/i_d2stg_nan_in2/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_nan_in2/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_nan_in2 ) );
  DFFX1 \fpu_div_ctl/i_d2stg_nan_in/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_nan_in/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_nan_in ), .QN(n41) );
  DFFX1 \fpu_div_ctl/i_d2stg_inf_in1/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_inf_in1/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_inf_in1 ), .QN(n40) );
  DFFX1 \fpu_div_ctl/i_d2stg_2inf_in/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d2stg_2inf_in/N3 ), .CLK(rclk), .Q(
        \fpu_div_ctl/d2stg_2inf_in ) );
  DFFX1 \fpu_div_ctl/i_div_nv_out/q_reg[0]  ( .D(n450), .CLK(rclk), .Q(
        div_exc_out[4]) );
  DFFX1 \fpu_div_ctl/i_d1stg_sngopa/q_reg[3]  ( .D(n511), .CLK(rclk), .Q(n1538), .QN(n37) );
  DFFSSRX1 \fpu_div_ctl/i_d2stg_infnan_in/q_reg[0]  ( .D(n35), .RSTB(n979), 
        .SETB(n1047), .CLK(rclk), .Q(n36), .QN(\fpu_div_ctl/d2stg_infnan_in )
         );
  DFFSSRX1 \fpu_div_exp_dp/i_div_exp1/q_reg[0]  ( .D(
        div_expadd1_in2_exp_in2_dbl), .RSTB(n291), .SETB(n282), .CLK(n577), 
        .Q(div_exp1[0]), .QN(n605) );
  DFFX1 \fpu_div_exp_dp/i_div_exp1/q_reg[1]  ( .D(n487), .CLK(n577), .Q(n1575), 
        .QN(n609) );
  DFFSSRX1 \fpu_div_exp_dp/i_div_exp1/q_reg[2]  ( .D(
        div_expadd1_in2_exp_in2_dbl), .RSTB(n291), .SETB(n285), .CLK(n577), 
        .Q(n1716), .QN(n596) );
  DFFSSRX1 \fpu_div_exp_dp/i_div_exp1/q_reg[3]  ( .D(n291), .RSTB(
        div_expadd1_in2_exp_in2_sng), .SETB(n286), .CLK(n577), .Q(div_exp1[3]), 
        .QN(n610) );
  DFFX1 \fpu_div_exp_dp/i_div_exp1/q_reg[4]  ( .D(n488), .CLK(n577), .Q(n1409), 
        .QN(n592) );
  DFFSSRX1 \fpu_div_exp_dp/i_div_exp1/q_reg[5]  ( .D(
        div_expadd1_in2_exp_in2_dbl), .RSTB(n291), .SETB(n289), .CLK(n577), 
        .Q(div_exp1[5]), .QN(n590) );
  DFFX1 \fpu_div_exp_dp/i_div_exp1/q_reg[6]  ( .D(n489), .CLK(n577), .Q(n1808), 
        .QN(n34) );
  DFFX1 \fpu_div_exp_dp/i_div_exp1/q_reg[7]  ( .D(n490), .CLK(n577), .Q(n1809), 
        .QN(n33) );
  DFFSSRX1 \fpu_div_exp_dp/i_div_exp1/q_reg[8]  ( .D(n291), .RSTB(
        div_expadd1_in2_exp_in2_sng), .SETB(n290), .CLK(n577), .Q(div_exp1[8]), 
        .QN(n32) );
  DFFX1 \fpu_div_exp_dp/i_div_exp1/q_reg[9]  ( .D(n491), .CLK(n577), .Q(n1817), 
        .QN(n31) );
  DFFX1 \fpu_div_exp_dp/i_div_exp1/q_reg[10]  ( .D(n492), .CLK(n577), .Q(n1815), .QN(n30) );
  DFFSSRX1 \fpu_div_exp_dp/i_div_exp1/q_reg[11]  ( .D(
        div_expadd1_in2_exp_in2_dbl), .RSTB(n291), .SETB(n292), .CLK(n577), 
        .Q(div_exp1[11]), .QN(n29) );
  DFFX1 \fpu_div_ctl/i_div_of_mask/q_reg[0]  ( .D(n448), .CLK(rclk), .Q(n1719), 
        .QN(n28) );
  DFFX1 \fpu_div_ctl/i_div_dz_out/q_reg[0]  ( .D(n452), .CLK(rclk), .Q(
        div_exc_out[1]) );
  DFFX1 \fpu_div_ctl/i_d1stg_sngopa/q_reg[4]  ( .D(n512), .CLK(rclk), .Q(
        \fpu_div_ctl/d1stg_sngopa[4] ) );
  DFFX1 \fpu_div_ctl/i_div_expadd1_in1_sng/q_reg[0]  ( .D(
        \fpu_div_ctl/i_div_expadd1_in1_sng/N3 ), .CLK(rclk), .Q(
        div_expadd1_in1_sng), .QN(n601) );
  DFFX1 \fpu_div_ctl/i_d1stg_dblop/q_reg[0]  ( .D(n507), .CLK(rclk), .Q(n1870), 
        .QN(n25) );
  DFFX1 \fpu_div_ctl/i_d1stg_sign1/q_reg[0]  ( .D(n494), .CLK(rclk), .Q(n1641), 
        .QN(n626) );
  DFFX1 \fpu_div_ctl/i_d1stg_sign2/q_reg[0]  ( .D(n493), .CLK(rclk), .Q(n1539)
         );
  DFFX1 \fpu_div_ctl/i_div_sign_out/q_reg[0]  ( .D(n449), .CLK(rclk), .Q(
        div_sign_out), .QN(n625) );
  DFFX1 \fpu_div_ctl/i_d6stg_opdec/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d6stg_opdec/N9 ), .CLK(rclk), .Q(n1397), .QN(n192) );
  DFFX1 \fpu_div_ctl/i_d7stg_opdec/q_reg[0]  ( .D(
        \fpu_div_ctl/i_d7stg_opdec/N9 ), .CLK(rclk), .Q(d7stg_fdivd), .QN(n22)
         );
  DFFX1 \fpu_div_ctl/i_d8stg_opdec/q_reg[0]  ( .D(n475), .CLK(rclk), .Q(
        d8stg_fdivd), .QN(n21) );
  DFFX1 \fpu_div_ctl/i_d5stg_fdiva/q_reg[0]  ( .D(n469), .CLK(rclk), .Q(n1579), 
        .QN(n576) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[12]  ( .D(n515), .CLK(n577), .Q(
        div_exp_out[12]), .QN(n613) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[0]  ( .D(n446), .CLK(n577), .Q(
        div_exp_out[0]), .QN(n218) );
  DFFX1 \fpu_div_ctl/i_div_of_out_tmp2/q_reg[0]  ( .D(n447), .CLK(rclk), .Q(
        n1873), .QN(n19) );
  DFFX1 \fpu_div_ctl/i_div_expadd2_no_decr_inv/q_reg[0]  ( .D(n437), .CLK(rclk), .Q(div_expadd2_no_decr_inv), .QN(n18) );
  DFFX1 \fpu_div_ctl/i_div_out_52_inv/q_reg[0]  ( .D(n474), .CLK(rclk), .Q(
        n1783), .QN(n205) );
  DFFX1 \fpu_div_ctl/i_d7stg_lsb/q_reg[0]  ( .D(n470), .CLK(rclk), .Q(n1874), 
        .QN(n17) );
  DFFX1 \fpu_div_ctl/i_d7stg_grd/q_reg[0]  ( .D(n472), .CLK(rclk), .Q(n1717), 
        .QN(n16) );
  DFFX1 \fpu_div_ctl/i_d7stg_stk/q_reg[0]  ( .D(n473), .CLK(rclk), .Q(n1536), 
        .QN(n15) );
  DFFX1 \fpu_div_ctl/i_div_nx_out/q_reg[0]  ( .D(n471), .CLK(rclk), .Q(
        \fpu_div_ctl/div_nx_out ), .QN(n14) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[11]  ( .D(n438), .CLK(n577), .Q(
        n1371), .QN(n618) );
  DFFSSRX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[10]  ( .D(d7stg_fdivd), .RSTB(
        n1355), .SETB(n246), .CLK(n577), .Q(div_exp_out[10]), .QN(n599) );
  DFFSSRX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[9]  ( .D(d7stg_fdivd), .RSTB(
        n1355), .SETB(n247), .CLK(n577), .Q(div_exp_out[9]), .QN(n580) );
  DFFSSRX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[8]  ( .D(d7stg_fdivd), .RSTB(
        n1355), .SETB(n248), .CLK(n577), .Q(div_exp_out[8]), .QN(n584) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[7]  ( .D(n439), .CLK(n577), .Q(
        div_exp_out[7]), .QN(n598) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[6]  ( .D(n440), .CLK(n577), .Q(
        div_exp_out[6]), .QN(n614) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[5]  ( .D(n441), .CLK(n577), .Q(
        div_exp_out[5]), .QN(n603) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[4]  ( .D(n442), .CLK(n577), .Q(
        div_exp_out[4]), .QN(n583) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[3]  ( .D(n443), .CLK(n577), .Q(
        div_exp_out[3]), .QN(n582) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[2]  ( .D(n444), .CLK(n577), .Q(
        div_exp_out[2]), .QN(n579) );
  DFFX1 \fpu_div_exp_dp/i_div_exp_out/q_reg[1]  ( .D(n445), .CLK(n577), .Q(
        div_exp_out[1]), .QN(n595) );
  DFFX1 \fpu_div_ctl/i_div_of_out_tmp1/q_reg[0]  ( .D(n436), .CLK(rclk), .Q(
        n1867), .QN(n2) );
  DFFX1 \fpu_div_ctl/i_div_uf_out/q_reg[0]  ( .D(n435), .CLK(rclk), .Q(
        div_exc_out[2]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[54]  ( .D(
        \fpu_div_frac_dp/n1056 ), .CLK(n1899), .Q(n1864), .QN(
        \fpu_div_frac_dp/n1 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[54]  ( .D(
        \fpu_div_frac_dp/n1058 ), .CLK(n1899), .Q(n1644) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[54]  ( .D(
        \fpu_div_frac_dp/n1057 ), .CLK(n1899), .Q(n1460) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[53]  ( .D(
        \fpu_div_frac_dp/n1113 ), .CLK(n1899), .Q(n1637), .QN(
        \fpu_div_frac_dp/n4 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[53]  ( .D(
        \fpu_div_frac_dp/n1059 ), .CLK(n1899), .Q(n1443) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[0]  ( .D(\fpu_div_frac_dp/n1219 ), .CLK(n1898), .Q(div_frac_outa[0]), .QN(\fpu_div_frac_dp/n6 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[0]  ( .D(
        \fpu_div_frac_dp/n1166 ), .CLK(n1901), .Q(n1362) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[0]  ( .D(
        \fpu_div_frac_dp/n1112 ), .CLK(n1901), .Q(n1527), .QN(
        \fpu_div_frac_dp/n8 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[1]  ( .D(\fpu_div_frac_dp/n1218 ), .CLK(n1898), .Q(div_frac_outa[1]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[1]  ( .D(
        \fpu_div_frac_dp/n1165 ), .CLK(n1898), .Q(n1512), .QN(
        \fpu_div_frac_dp/n10 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[1]  ( .D(
        \fpu_div_frac_dp/n1111 ), .CLK(n1901), .Q(n1623), .QN(
        \fpu_div_frac_dp/n11 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[2]  ( .D(\fpu_div_frac_dp/n1217 ), .CLK(n1901), .Q(div_frac_outa[2]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[2]  ( .D(
        \fpu_div_frac_dp/n1164 ), .CLK(n1901), .Q(n1493), .QN(
        \fpu_div_frac_dp/n13 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[2]  ( .D(
        \fpu_div_frac_dp/n1110 ), .CLK(n1901), .Q(n1622), .QN(
        \fpu_div_frac_dp/n14 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[3]  ( .D(\fpu_div_frac_dp/n1216 ), .CLK(n1902), .Q(div_frac_outa[3]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[3]  ( .D(
        \fpu_div_frac_dp/n1163 ), .CLK(n1902), .Q(n1513), .QN(
        \fpu_div_frac_dp/n16 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[3]  ( .D(
        \fpu_div_frac_dp/n1109 ), .CLK(n1902), .Q(n1621), .QN(
        \fpu_div_frac_dp/n17 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[4]  ( .D(\fpu_div_frac_dp/n1215 ), .CLK(n1902), .Q(div_frac_outa[4]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[4]  ( .D(
        \fpu_div_frac_dp/n1162 ), .CLK(n1898), .Q(n1516), .QN(
        \fpu_div_frac_dp/n19 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[4]  ( .D(
        \fpu_div_frac_dp/n1108 ), .CLK(n1901), .Q(n1620), .QN(
        \fpu_div_frac_dp/n20 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[5]  ( .D(\fpu_div_frac_dp/n1214 ), .CLK(n1902), .Q(div_frac_outa[5]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[5]  ( .D(
        \fpu_div_frac_dp/n1161 ), .CLK(n1902), .Q(n1404) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[5]  ( .D(
        \fpu_div_frac_dp/n1107 ), .CLK(n1902), .Q(n1596) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[6]  ( .D(\fpu_div_frac_dp/n1213 ), .CLK(n1902), .Q(div_frac_outa[6]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[6]  ( .D(
        \fpu_div_frac_dp/n1160 ), .CLK(n1902), .Q(n1379) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[6]  ( .D(
        \fpu_div_frac_dp/n1106 ), .CLK(n1902), .Q(n1595) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[7]  ( .D(\fpu_div_frac_dp/n1212 ), .CLK(n1902), .Q(div_frac_outa[7]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[7]  ( .D(
        \fpu_div_frac_dp/n1159 ), .CLK(n1898), .Q(n1365) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[7]  ( .D(
        \fpu_div_frac_dp/n1105 ), .CLK(n1901), .Q(n1594) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[8]  ( .D(\fpu_div_frac_dp/n1211 ), .CLK(n1902), .Q(div_frac_outa[8]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[8]  ( .D(
        \fpu_div_frac_dp/n1158 ), .CLK(n1903), .Q(n1359) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[8]  ( .D(
        \fpu_div_frac_dp/n1104 ), .CLK(n1903), .Q(n1593) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[9]  ( .D(\fpu_div_frac_dp/n1210 ), .CLK(n1903), .Q(div_frac_outa[9]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[9]  ( .D(
        \fpu_div_frac_dp/n1157 ), .CLK(n1903), .Q(n1366) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[9]  ( .D(
        \fpu_div_frac_dp/n1103 ), .CLK(n1903), .Q(n1592) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[10]  ( .D(
        \fpu_div_frac_dp/n1209 ), .CLK(n1903), .Q(div_frac_outa[10]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[10]  ( .D(
        \fpu_div_frac_dp/n1156 ), .CLK(n1898), .Q(n1380) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[10]  ( .D(
        \fpu_div_frac_dp/n1102 ), .CLK(n1901), .Q(n1591) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[11]  ( .D(
        \fpu_div_frac_dp/n1208 ), .CLK(n1903), .Q(div_frac_outa[11]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[11]  ( .D(
        \fpu_div_frac_dp/n1155 ), .CLK(n1903), .Q(n1517), .QN(
        \fpu_div_frac_dp/n40 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[11]  ( .D(
        \fpu_div_frac_dp/n1101 ), .CLK(n1903), .Q(n1590) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[12]  ( .D(
        \fpu_div_frac_dp/n1207 ), .CLK(n1903), .Q(div_frac_outa[12]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[12]  ( .D(
        \fpu_div_frac_dp/n1154 ), .CLK(n1903), .Q(n1500), .QN(
        \fpu_div_frac_dp/n43 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[12]  ( .D(
        \fpu_div_frac_dp/n1100 ), .CLK(n1904), .Q(n1586) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[13]  ( .D(
        \fpu_div_frac_dp/n1206 ), .CLK(n1903), .Q(div_frac_outa[13]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[13]  ( .D(
        \fpu_div_frac_dp/n1153 ), .CLK(n1898), .Q(n1358) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[13]  ( .D(
        \fpu_div_frac_dp/n1099 ), .CLK(n1901), .Q(n1589) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[14]  ( .D(
        \fpu_div_frac_dp/n1205 ), .CLK(n1904), .Q(div_frac_outa[14]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[14]  ( .D(
        \fpu_div_frac_dp/n1152 ), .CLK(n1904), .Q(n1363) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[14]  ( .D(
        \fpu_div_frac_dp/n1098 ), .CLK(n1904), .Q(n1585) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[15]  ( .D(
        \fpu_div_frac_dp/n1204 ), .CLK(n1904), .Q(div_frac_outa[15]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[15]  ( .D(
        \fpu_div_frac_dp/n1151 ), .CLK(n1904), .Q(n1405) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[15]  ( .D(
        \fpu_div_frac_dp/n1097 ), .CLK(n1904), .Q(n1584) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[16]  ( .D(
        \fpu_div_frac_dp/n1203 ), .CLK(n1904), .Q(div_frac_outa[16]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[16]  ( .D(
        \fpu_div_frac_dp/n1150 ), .CLK(n1898), .Q(n1381) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[16]  ( .D(
        \fpu_div_frac_dp/n1096 ), .CLK(n1901), .Q(n1588) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[17]  ( .D(
        \fpu_div_frac_dp/n1202 ), .CLK(n1904), .Q(div_frac_outa[17]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[17]  ( .D(
        \fpu_div_frac_dp/n1149 ), .CLK(n1904), .Q(n1501), .QN(
        \fpu_div_frac_dp/n58 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[17]  ( .D(
        \fpu_div_frac_dp/n1095 ), .CLK(n1904), .Q(n1583) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[18]  ( .D(
        \fpu_div_frac_dp/n1201 ), .CLK(n1905), .Q(div_frac_outa[18]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[18]  ( .D(
        \fpu_div_frac_dp/n1148 ), .CLK(n1905), .Q(n1518), .QN(
        \fpu_div_frac_dp/n61 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[18]  ( .D(
        \fpu_div_frac_dp/n1094 ), .CLK(n1905), .Q(n1582) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[19]  ( .D(
        \fpu_div_frac_dp/n1200 ), .CLK(n1904), .Q(div_frac_outa[19]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[19]  ( .D(
        \fpu_div_frac_dp/n1147 ), .CLK(n1898), .Q(n1502), .QN(
        \fpu_div_frac_dp/n64 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[19]  ( .D(
        \fpu_div_frac_dp/n1093 ), .CLK(n1901), .Q(n1587) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[20]  ( .D(
        \fpu_div_frac_dp/n1199 ), .CLK(n1905), .Q(div_frac_outa[20]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[20]  ( .D(
        \fpu_div_frac_dp/n1146 ), .CLK(n1905), .Q(n1357) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[20]  ( .D(
        \fpu_div_frac_dp/n1092 ), .CLK(n1905), .Q(n1581) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[21]  ( .D(
        \fpu_div_frac_dp/n1198 ), .CLK(n1905), .Q(div_frac_outa[21]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[21]  ( .D(
        \fpu_div_frac_dp/n1145 ), .CLK(n1905), .Q(n1406) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[21]  ( .D(
        \fpu_div_frac_dp/n1091 ), .CLK(n1905), .Q(n1470) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[22]  ( .D(
        \fpu_div_frac_dp/n1197 ), .CLK(n1905), .Q(div_frac_outa[22]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[22]  ( .D(
        \fpu_div_frac_dp/n1144 ), .CLK(n1898), .Q(n1382) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[22]  ( .D(
        \fpu_div_frac_dp/n1090 ), .CLK(n1900), .Q(n1469) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[23]  ( .D(
        \fpu_div_frac_dp/n1196 ), .CLK(n1905), .Q(div_frac_outa[23]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[23]  ( .D(
        \fpu_div_frac_dp/n1143 ), .CLK(n1905), .Q(n1503), .QN(
        \fpu_div_frac_dp/n76 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[23]  ( .D(
        \fpu_div_frac_dp/n1089 ), .CLK(n1906), .Q(n1468) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[24]  ( .D(
        \fpu_div_frac_dp/n1195 ), .CLK(n1906), .Q(div_frac_outa[24]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[24]  ( .D(
        \fpu_div_frac_dp/n1142 ), .CLK(n1906), .Q(n1519), .QN(
        \fpu_div_frac_dp/n79 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[24]  ( .D(
        \fpu_div_frac_dp/n1088 ), .CLK(n1906), .Q(n1467) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[26]  ( .D(
        \fpu_div_frac_dp/n1193 ), .CLK(n1906), .Q(div_frac_outa[26]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[25]  ( .D(
        \fpu_div_frac_dp/n1194 ), .CLK(n1906), .Q(div_frac_outa[25]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[25]  ( .D(
        \fpu_div_frac_dp/n1141 ), .CLK(n1898), .Q(n1504), .QN(
        \fpu_div_frac_dp/n83 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[25]  ( .D(
        \fpu_div_frac_dp/n1087 ), .CLK(n1900), .Q(n1466) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[27]  ( .D(
        \fpu_div_frac_dp/n1192 ), .CLK(n1906), .Q(div_frac_outa[27]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[27]  ( .D(
        \fpu_div_frac_dp/n1139 ), .CLK(n1906), .Q(n1402) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[27]  ( .D(
        \fpu_div_frac_dp/n1085 ), .CLK(n1906), .Q(n1464) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[26]  ( .D(
        \fpu_div_frac_dp/n1140 ), .CLK(n1906), .Q(n1377) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[26]  ( .D(
        \fpu_div_frac_dp/n1086 ), .CLK(n1906), .Q(n1465) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[28]  ( .D(
        \fpu_div_frac_dp/n1191 ), .CLK(n1906), .Q(div_frac_outa[28]), .QN(
        \fpu_div_frac_dp/n993 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[28]  ( .D(
        \fpu_div_frac_dp/n1138 ), .CLK(n1898), .Q(n1361) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[28]  ( .D(
        \fpu_div_frac_dp/n1084 ), .CLK(n1900), .Q(n1463) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[29]  ( .D(
        \fpu_div_frac_dp/n1190 ), .CLK(n1907), .Q(div_frac_outa[29]), .QN(
        \fpu_div_frac_dp/n92 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[29]  ( .D(
        \fpu_div_frac_dp/n1137 ), .CLK(n1907), .Q(n1537), .QN(
        \fpu_div_frac_dp/n93 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[29]  ( .D(
        \fpu_div_frac_dp/n1083 ), .CLK(n1907), .Q(n1612), .QN(
        \fpu_div_frac_dp/n94 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[30]  ( .D(
        \fpu_div_frac_dp/n1189 ), .CLK(n1907), .Q(div_frac_outa[30]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[30]  ( .D(
        \fpu_div_frac_dp/n1136 ), .CLK(n1907), .Q(n1520), .QN(
        \fpu_div_frac_dp/n96 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[30]  ( .D(
        \fpu_div_frac_dp/n1082 ), .CLK(n1907), .Q(n1462) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[31]  ( .D(
        \fpu_div_frac_dp/n1188 ), .CLK(n1907), .Q(div_frac_outa[31]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[31]  ( .D(
        \fpu_div_frac_dp/n1135 ), .CLK(n1899), .Q(n1505), .QN(
        \fpu_div_frac_dp/n99 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[31]  ( .D(
        \fpu_div_frac_dp/n1081 ), .CLK(n1900), .Q(n1619), .QN(
        \fpu_div_frac_dp/n100 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[32]  ( .D(
        \fpu_div_frac_dp/n1187 ), .CLK(n1907), .Q(div_frac_outa[32]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[32]  ( .D(
        \fpu_div_frac_dp/n1134 ), .CLK(n1907), .Q(n1506), .QN(
        \fpu_div_frac_dp/n102 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[32]  ( .D(
        \fpu_div_frac_dp/n1080 ), .CLK(n1907), .Q(n1611), .QN(
        \fpu_div_frac_dp/n103 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[33]  ( .D(
        \fpu_div_frac_dp/n1186 ), .CLK(n1907), .Q(div_frac_outa[33]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[33]  ( .D(
        \fpu_div_frac_dp/n1133 ), .CLK(n1908), .Q(n1507), .QN(
        \fpu_div_frac_dp/n105 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[33]  ( .D(
        \fpu_div_frac_dp/n1079 ), .CLK(n1908), .Q(n1610), .QN(
        \fpu_div_frac_dp/n106 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[34]  ( .D(
        \fpu_div_frac_dp/n1185 ), .CLK(n1907), .Q(div_frac_outa[34]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[34]  ( .D(
        \fpu_div_frac_dp/n1132 ), .CLK(n1899), .Q(n1521), .QN(
        \fpu_div_frac_dp/n108 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[34]  ( .D(
        \fpu_div_frac_dp/n1078 ), .CLK(n1900), .Q(n1618), .QN(
        \fpu_div_frac_dp/n109 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[35]  ( .D(
        \fpu_div_frac_dp/n1184 ), .CLK(n1908), .Q(div_frac_outa[35]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[35]  ( .D(
        \fpu_div_frac_dp/n1131 ), .CLK(n1908), .Q(n1494), .QN(
        \fpu_div_frac_dp/n111 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[35]  ( .D(
        \fpu_div_frac_dp/n1077 ), .CLK(n1908), .Q(n1609), .QN(
        \fpu_div_frac_dp/n112 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[36]  ( .D(
        \fpu_div_frac_dp/n1183 ), .CLK(n1908), .Q(div_frac_outa[36]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[36]  ( .D(
        \fpu_div_frac_dp/n1130 ), .CLK(n1908), .Q(n1497), .QN(
        \fpu_div_frac_dp/n114 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[36]  ( .D(
        \fpu_div_frac_dp/n1076 ), .CLK(n1908), .Q(n1608), .QN(
        \fpu_div_frac_dp/n115 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[37]  ( .D(
        \fpu_div_frac_dp/n1182 ), .CLK(n1908), .Q(div_frac_outa[37]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[37]  ( .D(
        \fpu_div_frac_dp/n1129 ), .CLK(n1899), .Q(n1495), .QN(
        \fpu_div_frac_dp/n117 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[37]  ( .D(
        \fpu_div_frac_dp/n1075 ), .CLK(n1900), .Q(n1617), .QN(
        \fpu_div_frac_dp/n118 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[38]  ( .D(
        \fpu_div_frac_dp/n1181 ), .CLK(n1908), .Q(div_frac_outa[38]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[38]  ( .D(
        \fpu_div_frac_dp/n1128 ), .CLK(n1908), .Q(n1514), .QN(
        \fpu_div_frac_dp/n120 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[38]  ( .D(
        \fpu_div_frac_dp/n1074 ), .CLK(n1908), .Q(n1607), .QN(
        \fpu_div_frac_dp/n121 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[39]  ( .D(
        \fpu_div_frac_dp/n1180 ), .CLK(n1909), .Q(div_frac_outa[39]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[39]  ( .D(
        \fpu_div_frac_dp/n1127 ), .CLK(n1909), .Q(n1508), .QN(
        \fpu_div_frac_dp/n123 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[39]  ( .D(
        \fpu_div_frac_dp/n1073 ), .CLK(n1909), .Q(n1606), .QN(
        \fpu_div_frac_dp/n124 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[40]  ( .D(
        \fpu_div_frac_dp/n1179 ), .CLK(n1909), .Q(div_frac_outa[40]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[40]  ( .D(
        \fpu_div_frac_dp/n1126 ), .CLK(n1899), .Q(n1509), .QN(
        \fpu_div_frac_dp/n126 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[40]  ( .D(
        \fpu_div_frac_dp/n1072 ), .CLK(n1900), .Q(n1616), .QN(
        \fpu_div_frac_dp/n127 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[41]  ( .D(
        \fpu_div_frac_dp/n1178 ), .CLK(n1909), .Q(div_frac_outa[41]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[41]  ( .D(
        \fpu_div_frac_dp/n1125 ), .CLK(n1909), .Q(n1522), .QN(
        \fpu_div_frac_dp/n129 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[41]  ( .D(
        \fpu_div_frac_dp/n1071 ), .CLK(n1909), .Q(n1605), .QN(
        \fpu_div_frac_dp/n130 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[42]  ( .D(
        \fpu_div_frac_dp/n1177 ), .CLK(n1909), .Q(div_frac_outa[42]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[42]  ( .D(
        \fpu_div_frac_dp/n1124 ), .CLK(n1909), .Q(n1498), .QN(
        \fpu_div_frac_dp/n132 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[42]  ( .D(
        \fpu_div_frac_dp/n1070 ), .CLK(n1909), .Q(n1604), .QN(
        \fpu_div_frac_dp/n133 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[43]  ( .D(
        \fpu_div_frac_dp/n1176 ), .CLK(n1909), .Q(div_frac_outa[43]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[43]  ( .D(
        \fpu_div_frac_dp/n1123 ), .CLK(n1899), .Q(n1496), .QN(
        \fpu_div_frac_dp/n135 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[43]  ( .D(
        \fpu_div_frac_dp/n1069 ), .CLK(n1900), .Q(n1615), .QN(
        \fpu_div_frac_dp/n136 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[44]  ( .D(
        \fpu_div_frac_dp/n1175 ), .CLK(n1909), .Q(div_frac_outa[44]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[44]  ( .D(
        \fpu_div_frac_dp/n1122 ), .CLK(n1910), .Q(n1515), .QN(
        \fpu_div_frac_dp/n138 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[44]  ( .D(
        \fpu_div_frac_dp/n1068 ), .CLK(n1910), .Q(n1603), .QN(
        \fpu_div_frac_dp/n139 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[45]  ( .D(
        \fpu_div_frac_dp/n1174 ), .CLK(n1910), .Q(div_frac_outa[45]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[45]  ( .D(
        \fpu_div_frac_dp/n1121 ), .CLK(n1910), .Q(n1510), .QN(
        \fpu_div_frac_dp/n141 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[45]  ( .D(
        \fpu_div_frac_dp/n1067 ), .CLK(n1910), .Q(n1602), .QN(
        \fpu_div_frac_dp/n142 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[46]  ( .D(
        \fpu_div_frac_dp/n1173 ), .CLK(n1910), .Q(div_frac_outa[46]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[46]  ( .D(
        \fpu_div_frac_dp/n1120 ), .CLK(n1899), .Q(n1511), .QN(
        \fpu_div_frac_dp/n144 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[46]  ( .D(
        \fpu_div_frac_dp/n1066 ), .CLK(n1900), .Q(n1614), .QN(
        \fpu_div_frac_dp/n145 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[47]  ( .D(
        \fpu_div_frac_dp/n1172 ), .CLK(n1910), .Q(div_frac_outa[47]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[47]  ( .D(
        \fpu_div_frac_dp/n1119 ), .CLK(n1910), .Q(n1523), .QN(
        \fpu_div_frac_dp/n147 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[47]  ( .D(
        \fpu_div_frac_dp/n1065 ), .CLK(n1910), .Q(n1601), .QN(
        \fpu_div_frac_dp/n148 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[48]  ( .D(
        \fpu_div_frac_dp/n1171 ), .CLK(n1910), .Q(div_frac_outa[48]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[48]  ( .D(
        \fpu_div_frac_dp/n1118 ), .CLK(n1910), .Q(n1378) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[48]  ( .D(
        \fpu_div_frac_dp/n1064 ), .CLK(n1911), .Q(n1600), .QN(
        \fpu_div_frac_dp/n151 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[49]  ( .D(
        \fpu_div_frac_dp/n1170 ), .CLK(n1910), .Q(div_frac_outa[49]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[49]  ( .D(
        \fpu_div_frac_dp/n1117 ), .CLK(n1899), .Q(n1407) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[49]  ( .D(
        \fpu_div_frac_dp/n1063 ), .CLK(n1900), .Q(n1613), .QN(
        \fpu_div_frac_dp/n154 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[51]  ( .D(
        \fpu_div_frac_dp/n1168 ), .CLK(n1911), .Q(div_frac_outa[51]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[50]  ( .D(
        \fpu_div_frac_dp/n1169 ), .CLK(n1911), .Q(div_frac_outa[50]) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[50]  ( .D(
        \fpu_div_frac_dp/n1116 ), .CLK(n1911), .Q(n1364) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[50]  ( .D(
        \fpu_div_frac_dp/n1062 ), .CLK(n1911), .Q(n1599), .QN(
        \fpu_div_frac_dp/n158 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[52]  ( .D(
        \fpu_div_frac_dp/n1167 ), .CLK(n1911), .Q(n1383) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[52]  ( .D(
        \fpu_div_frac_dp/n1114 ), .CLK(n1900), .Q(n1636), .QN(
        \fpu_div_frac_dp/n160 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[52]  ( .D(
        \fpu_div_frac_dp/n1060 ), .CLK(n1900), .Q(n1399) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1/q_reg[51]  ( .D(
        \fpu_div_frac_dp/n1115 ), .CLK(n1911), .Q(n1526), .QN(
        \fpu_div_frac_dp/n162 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in1a/q_reg[51]  ( .D(
        \fpu_div_frac_dp/n1061 ), .CLK(n1911), .Q(n1598), .QN(
        \fpu_div_frac_dp/n163 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_out/q_reg[53]  ( .D(
        \fpu_div_frac_dp/n1220 ), .CLK(n1911), .Q(n1529), .QN(
        \fpu_div_frac_dp/n164 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[54]  ( .D(
        \fpu_div_frac_dp/n1221 ), .CLK(\fpu_div_frac_dp/n985 ), .Q(n1866), 
        .QN(\fpu_div_frac_dp/n165 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[53]  ( .D(
        \fpu_div_frac_dp/n1222 ), .CLK(\fpu_div_frac_dp/n985 ), .Q(n1635), 
        .QN(\fpu_div_frac_dp/n166 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[52]  ( .D(
        \fpu_div_frac_dp/n1223 ), .CLK(n1919), .Q(n1578), .QN(
        \fpu_div_frac_dp/n995 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[51]  ( .D(
        \fpu_div_frac_dp/n1224 ), .CLK(n1917), .Q(n1439), .QN(
        \fpu_div_frac_dp/n992 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[50]  ( .D(
        \fpu_div_frac_dp/n1225 ), .CLK(n1913), .Q(n1440), .QN(
        \fpu_div_frac_dp/n991 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[49]  ( .D(
        \fpu_div_frac_dp/n1226 ), .CLK(n1915), .Q(n1441), .QN(
        \fpu_div_frac_dp/n990 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[48]  ( .D(
        \fpu_div_frac_dp/n1227 ), .CLK(n1919), .Q(n1471) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[47]  ( .D(
        \fpu_div_frac_dp/n1228 ), .CLK(n1916), .Q(n1472) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[46]  ( .D(
        \fpu_div_frac_dp/n1229 ), .CLK(n1913), .Q(n1473) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[45]  ( .D(
        \fpu_div_frac_dp/n1230 ), .CLK(n1914), .Q(n1474) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[44]  ( .D(
        \fpu_div_frac_dp/n1231 ), .CLK(n1918), .Q(n1475) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[43]  ( .D(
        \fpu_div_frac_dp/n1232 ), .CLK(n1916), .Q(n1476) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[42]  ( .D(
        \fpu_div_frac_dp/n1233 ), .CLK(n1913), .Q(n1477) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[41]  ( .D(
        \fpu_div_frac_dp/n1234 ), .CLK(n1914), .Q(n1478) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[40]  ( .D(
        \fpu_div_frac_dp/n1235 ), .CLK(n1918), .Q(n1479) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[39]  ( .D(
        \fpu_div_frac_dp/n1236 ), .CLK(n1916), .Q(n1480) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[38]  ( .D(
        \fpu_div_frac_dp/n1237 ), .CLK(n1912), .Q(n1481) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[37]  ( .D(
        \fpu_div_frac_dp/n1238 ), .CLK(n1914), .Q(n1482) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[36]  ( .D(
        \fpu_div_frac_dp/n1239 ), .CLK(n1919), .Q(n1483) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[35]  ( .D(
        \fpu_div_frac_dp/n1240 ), .CLK(n1917), .Q(n1484) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[34]  ( .D(
        \fpu_div_frac_dp/n1241 ), .CLK(n1912), .Q(n1485) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[33]  ( .D(
        \fpu_div_frac_dp/n1242 ), .CLK(n1914), .Q(n1486) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[32]  ( .D(
        \fpu_div_frac_dp/n1243 ), .CLK(n1918), .Q(n1487) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[31]  ( .D(
        \fpu_div_frac_dp/n1244 ), .CLK(n1916), .Q(n1488) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[30]  ( .D(
        \fpu_div_frac_dp/n1245 ), .CLK(n1913), .Q(n1624), .QN(
        \fpu_div_frac_dp/n189 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[29]  ( .D(
        \fpu_div_frac_dp/n1246 ), .CLK(n1914), .Q(n1442), .QN(
        \fpu_div_frac_dp/n987 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[28]  ( .D(
        \fpu_div_frac_dp/n1247 ), .CLK(n1918), .Q(n1625), .QN(
        \fpu_div_frac_dp/n191 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[27]  ( .D(
        \fpu_div_frac_dp/n1248 ), .CLK(n1916), .Q(n1626), .QN(
        \fpu_div_frac_dp/n192 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[26]  ( .D(
        \fpu_div_frac_dp/n1249 ), .CLK(n1912), .Q(n1627), .QN(
        \fpu_div_frac_dp/n193 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[25]  ( .D(
        \fpu_div_frac_dp/n1250 ), .CLK(n1914), .Q(n1628), .QN(
        \fpu_div_frac_dp/n194 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[24]  ( .D(
        \fpu_div_frac_dp/n1251 ), .CLK(n1919), .Q(n1629), .QN(
        \fpu_div_frac_dp/n195 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[23]  ( .D(
        \fpu_div_frac_dp/n1252 ), .CLK(n1917), .Q(n1630), .QN(
        \fpu_div_frac_dp/n196 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[22]  ( .D(
        \fpu_div_frac_dp/n1253 ), .CLK(n1912), .Q(n1631), .QN(
        \fpu_div_frac_dp/n197 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[21]  ( .D(
        \fpu_div_frac_dp/n1254 ), .CLK(n1915), .Q(n1632), .QN(
        \fpu_div_frac_dp/n198 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[20]  ( .D(
        \fpu_div_frac_dp/n1255 ), .CLK(n1920), .Q(n1444), .QN(
        \fpu_div_frac_dp/n199 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[19]  ( .D(
        \fpu_div_frac_dp/n1256 ), .CLK(n1918), .Q(n1445), .QN(
        \fpu_div_frac_dp/n200 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[18]  ( .D(
        \fpu_div_frac_dp/n1257 ), .CLK(n1913), .Q(n1446), .QN(
        \fpu_div_frac_dp/n201 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[17]  ( .D(
        \fpu_div_frac_dp/n1258 ), .CLK(n1916), .Q(n1447), .QN(
        \fpu_div_frac_dp/n202 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[16]  ( .D(
        \fpu_div_frac_dp/n1259 ), .CLK(n1920), .Q(n1448), .QN(
        \fpu_div_frac_dp/n203 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[15]  ( .D(
        \fpu_div_frac_dp/n1260 ), .CLK(n1918), .Q(n1449), .QN(
        \fpu_div_frac_dp/n204 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[14]  ( .D(
        \fpu_div_frac_dp/n1261 ), .CLK(n1913), .Q(n1450), .QN(
        \fpu_div_frac_dp/n205 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[13]  ( .D(
        \fpu_div_frac_dp/n1262 ), .CLK(n1915), .Q(n1451), .QN(
        \fpu_div_frac_dp/n206 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[12]  ( .D(
        \fpu_div_frac_dp/n1263 ), .CLK(n1920), .Q(n1452), .QN(
        \fpu_div_frac_dp/n207 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[11]  ( .D(
        \fpu_div_frac_dp/n1264 ), .CLK(n1917), .Q(n1453), .QN(
        \fpu_div_frac_dp/n208 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[10]  ( .D(
        \fpu_div_frac_dp/n1265 ), .CLK(n1912), .Q(n1454), .QN(
        \fpu_div_frac_dp/n209 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[9]  ( .D(
        \fpu_div_frac_dp/n1266 ), .CLK(n1915), .Q(n1455), .QN(
        \fpu_div_frac_dp/n210 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[8]  ( .D(
        \fpu_div_frac_dp/n1267 ), .CLK(n1919), .Q(n1456), .QN(
        \fpu_div_frac_dp/n211 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[7]  ( .D(
        \fpu_div_frac_dp/n1268 ), .CLK(n1917), .Q(n1457), .QN(
        \fpu_div_frac_dp/n212 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[6]  ( .D(
        \fpu_div_frac_dp/n1269 ), .CLK(n1912), .Q(n1458), .QN(
        \fpu_div_frac_dp/n213 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[5]  ( .D(
        \fpu_div_frac_dp/n1270 ), .CLK(n1915), .Q(n1459), .QN(
        \fpu_div_frac_dp/n214 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[4]  ( .D(
        \fpu_div_frac_dp/n1271 ), .CLK(n1920), .Q(n1434) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[3]  ( .D(
        \fpu_div_frac_dp/n1272 ), .CLK(n1917), .Q(n1435) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[2]  ( .D(
        \fpu_div_frac_dp/n1273 ), .CLK(n1911), .Q(n1436) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[1]  ( .D(
        \fpu_div_frac_dp/n1274 ), .CLK(n1915), .Q(n1437) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_add_in2/q_reg[0]  ( .D(
        \fpu_div_frac_dp/n1275 ), .CLK(n1919), .Q(n1683), .QN(
        \fpu_div_frac_dp/n997 ) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[52]  ( .D(
        \fpu_div_frac_dp/n1277 ), .CLK(n1919), .Q(n1718) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[51]  ( .D(
        \fpu_div_frac_dp/n1278 ), .CLK(n1917), .Q(n1728) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[50]  ( .D(
        \fpu_div_frac_dp/n1279 ), .CLK(n1913), .Q(n1727) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[49]  ( .D(
        \fpu_div_frac_dp/n1280 ), .CLK(n1914), .Q(n1726) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[48]  ( .D(
        \fpu_div_frac_dp/n1281 ), .CLK(n1918), .Q(n1780) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[47]  ( .D(
        \fpu_div_frac_dp/n1282 ), .CLK(n1916), .Q(n1779) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[46]  ( .D(
        \fpu_div_frac_dp/n1283 ), .CLK(n1913), .Q(n1778) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[45]  ( .D(
        \fpu_div_frac_dp/n1284 ), .CLK(n1914), .Q(n1777) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[44]  ( .D(
        \fpu_div_frac_dp/n1285 ), .CLK(n1918), .Q(n1776) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[43]  ( .D(
        \fpu_div_frac_dp/n1286 ), .CLK(n1916), .Q(n1775) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[42]  ( .D(
        \fpu_div_frac_dp/n1287 ), .CLK(n1912), .Q(n1774) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[41]  ( .D(
        \fpu_div_frac_dp/n1288 ), .CLK(n1914), .Q(n1773) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[40]  ( .D(
        \fpu_div_frac_dp/n1289 ), .CLK(n1918), .Q(n1772) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[39]  ( .D(
        \fpu_div_frac_dp/n1290 ), .CLK(n1916), .Q(n1771) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[38]  ( .D(
        \fpu_div_frac_dp/n1291 ), .CLK(n1912), .Q(n1770) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[37]  ( .D(
        \fpu_div_frac_dp/n1292 ), .CLK(n1913), .Q(n1769) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[36]  ( .D(
        \fpu_div_frac_dp/n1293 ), .CLK(n1919), .Q(n1768) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[35]  ( .D(
        \fpu_div_frac_dp/n1294 ), .CLK(n1916), .Q(n1767) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[34]  ( .D(
        \fpu_div_frac_dp/n1295 ), .CLK(n1911), .Q(n1766) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[33]  ( .D(
        \fpu_div_frac_dp/n1296 ), .CLK(n1914), .Q(n1765) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[32]  ( .D(
        \fpu_div_frac_dp/n1297 ), .CLK(n1918), .Q(n1764) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[31]  ( .D(
        \fpu_div_frac_dp/n1298 ), .CLK(n1916), .Q(n1763) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[30]  ( .D(
        \fpu_div_frac_dp/n1299 ), .CLK(n1913), .Q(n1762) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[29]  ( .D(
        \fpu_div_frac_dp/n1300 ), .CLK(n1914), .Q(n1761) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[28]  ( .D(
        \fpu_div_frac_dp/n1301 ), .CLK(n1918), .Q(n1760) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[27]  ( .D(
        \fpu_div_frac_dp/n1302 ), .CLK(n1916), .Q(n1759) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[26]  ( .D(
        \fpu_div_frac_dp/n1303 ), .CLK(n1912), .Q(n1758) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[25]  ( .D(
        \fpu_div_frac_dp/n1304 ), .CLK(n1914), .Q(n1757) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[24]  ( .D(
        \fpu_div_frac_dp/n1305 ), .CLK(n1919), .Q(n1756) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[23]  ( .D(
        \fpu_div_frac_dp/n1306 ), .CLK(n1917), .Q(n1755) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[22]  ( .D(
        \fpu_div_frac_dp/n1307 ), .CLK(n1912), .Q(n1754) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[21]  ( .D(
        \fpu_div_frac_dp/n1308 ), .CLK(n1915), .Q(n1753) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[20]  ( .D(
        \fpu_div_frac_dp/n1309 ), .CLK(n1920), .Q(n1752) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[19]  ( .D(
        \fpu_div_frac_dp/n1310 ), .CLK(n1918), .Q(n1751) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[18]  ( .D(
        \fpu_div_frac_dp/n1311 ), .CLK(n1913), .Q(n1750) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[17]  ( .D(
        \fpu_div_frac_dp/n1312 ), .CLK(n1915), .Q(n1749) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[16]  ( .D(
        \fpu_div_frac_dp/n1313 ), .CLK(n1920), .Q(n1748) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[15]  ( .D(
        \fpu_div_frac_dp/n1314 ), .CLK(n1917), .Q(n1747) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[14]  ( .D(
        \fpu_div_frac_dp/n1315 ), .CLK(n1913), .Q(n1746) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[13]  ( .D(
        \fpu_div_frac_dp/n1316 ), .CLK(n1915), .Q(n1745) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[12]  ( .D(
        \fpu_div_frac_dp/n1317 ), .CLK(n1919), .Q(n1744) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[11]  ( .D(
        \fpu_div_frac_dp/n1318 ), .CLK(n1917), .Q(n1743) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[10]  ( .D(
        \fpu_div_frac_dp/n1319 ), .CLK(n1912), .Q(n1742) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[9]  ( .D(\fpu_div_frac_dp/n1320 ), .CLK(n1915), .Q(n1741) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[8]  ( .D(\fpu_div_frac_dp/n1321 ), .CLK(n1919), .Q(n1740) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[7]  ( .D(\fpu_div_frac_dp/n1322 ), .CLK(n1917), .Q(n1739) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[6]  ( .D(\fpu_div_frac_dp/n1323 ), .CLK(n1912), .Q(n1738) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[5]  ( .D(\fpu_div_frac_dp/n1324 ), .CLK(n1915), .Q(n1737) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[4]  ( .D(\fpu_div_frac_dp/n1325 ), .CLK(n1920), .Q(n1736) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[3]  ( .D(\fpu_div_frac_dp/n1326 ), .CLK(n1917), .Q(n1735) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[2]  ( .D(\fpu_div_frac_dp/n1327 ), .CLK(n1911), .Q(n1734) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[1]  ( .D(\fpu_div_frac_dp/n1328 ), .CLK(n1915), .Q(n1733) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_save/q_reg[0]  ( .D(\fpu_div_frac_dp/n1329 ), .CLK(n1919), .Q(n1729) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[52]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N55 ), .CLK(n1921), .Q(
        \fpu_div_frac_dp/div_shl_data[52] ) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[51]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N54 ), .CLK(n1921), .Q(n1721) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[50]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N53 ), .CLK(n1921), .Q(n1530) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[49]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N52 ), .CLK(n1921), .Q(n1567) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[48]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N51 ), .CLK(n1921), .Q(n1424) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[47]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N50 ), .CLK(n1921), .Q(n1565) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[46]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N49 ), .CLK(n1922), .Q(n1423) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[45]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N48 ), .CLK(n1922), .Q(n1566) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[44]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N47 ), .CLK(n1922), .Q(n1422) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[43]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N46 ), .CLK(n1922), .Q(n1563) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[42]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N45 ), .CLK(n1922), .Q(n1421) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[41]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N44 ), .CLK(n1922), .Q(n1564) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[40]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N43 ), .CLK(n1923), .Q(n1420) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[39]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N42 ), .CLK(n1923), .Q(n1561) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[38]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N41 ), .CLK(n1923), .Q(n1419) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[37]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N40 ), .CLK(n1923), .Q(n1562) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[36]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N39 ), .CLK(n1923), .Q(n1416) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[35]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N38 ), .CLK(n1923), .Q(n1557) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[34]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N37 ), .CLK(n1924), .Q(n1415) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[33]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N36 ), .CLK(n1924), .Q(n1558) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[32]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N35 ), .CLK(n1924), .Q(n1418) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[31]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N34 ), .CLK(n1924), .Q(n1559) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[30]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N33 ), .CLK(n1924), .Q(n1417) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[29]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N32 ), .CLK(n1924), .Q(n1560) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[28]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N31 ), .CLK(n1926), .Q(n1412) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[27]  ( .D(\fpu_div_frac_dp/n609 ), .CLK(n1926), .Q(n1553) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[26]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N29 ), .CLK(n1926), .Q(n1411) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[25]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N28 ), .CLK(n1926), .Q(n1554) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[24]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N27 ), .CLK(n1926), .Q(n1414) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[23]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N26 ), .CLK(n1926), .Q(n1555) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[22]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N25 ), .CLK(n1927), .Q(n1413) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[21]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N24 ), .CLK(n1927), .Q(n1556) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[20]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N23 ), .CLK(n1927), .Q(n1430) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[19]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N22 ), .CLK(n1927), .Q(n1571) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[18]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N21 ), .CLK(n1927), .Q(n1429) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[17]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N20 ), .CLK(n1927), .Q(n1572) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[16]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N19 ), .CLK(n1898), .Q(n1432) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[15]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N18 ), .CLK(n1904), .Q(n1573) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[14]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N17 ), .CLK(n1906), .Q(n1431) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[13]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N16 ), .CLK(n1908), .Q(n1574) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[12]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N15 ), .CLK(n1910), .Q(n1385) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[11]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N14 ), .CLK(n1913), .Q(n1370) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[10]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N13 ), .CLK(n1914), .Q(n1384) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[9]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N12 ), .CLK(n1899), .Q(n1426) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[8]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N11 ), .CLK(n1919), .Q(n1570) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[7]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N10 ), .CLK(n1916), .Q(n1427) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[6]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N9 ), .CLK(n1925), .Q(n1569) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[5]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N8 ), .CLK(n1925), .Q(n1428) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[4]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N7 ), .CLK(n1925), .Q(n1568) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[3]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N6 ), .CLK(n1925), .Q(n1425) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[2]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N5 ), .CLK(n1925), .Q(n1638), .QN(
        \fpu_div_frac_dp/n324 ) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[1]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N4 ), .CLK(n1925), .Q(n1533), .QN(
        \fpu_div_frac_dp/n325 ) );
  DFFX1 \fpu_div_frac_dp/i_div_shl_data/q_reg[0]  ( .D(
        \fpu_div_frac_dp/i_div_shl_data/N3 ), .CLK(n1920), .Q(n1646), .QN(
        \fpu_div_frac_dp/n326 ) );
  DFFX1 \fpu_div_frac_dp/i_dstg_xtra_regs/q_reg[11]  ( .D(
        \fpu_div_frac_dp/n602 ), .CLK(n1921), .Q(n1540), .QN(
        \fpu_div_frac_dp/n978 ) );
  DFFX1 \fpu_div_frac_dp/i_dstg_xtra_regs/q_reg[10]  ( .D(
        \fpu_div_frac_dp/i_dstg_xtra_regs/N7 ), .CLK(n1920), .Q(n1392), .QN(
        \fpu_div_frac_dp/n967 ) );
  DFFX1 \fpu_div_frac_dp/i_dstg_xtra_regs/q_reg[9]  ( .D(
        \fpu_div_frac_dp/i_dstg_xtra_regs/N6 ), .CLK(n1920), .Q(n1546), .QN(
        \fpu_div_frac_dp/n980 ) );
  DFFX1 \fpu_div_frac_dp/i_dstg_xtra_regs/q_reg[8]  ( .D(
        \fpu_div_frac_dp/i_dstg_xtra_regs/N5 ), .CLK(n1920), .Q(n1394), .QN(
        \fpu_div_frac_dp/n968 ) );
  DFFX1 \fpu_div_frac_dp/i_dstg_xtra_regs/q_reg[7]  ( .D(
        \fpu_div_frac_dp/i_dstg_xtra_regs/N4 ), .CLK(n1920), .Q(n1544), .QN(
        \fpu_div_frac_dp/n994 ) );
  DFFX1 \fpu_div_frac_dp/i_dstg_xtra_regs/q_reg[6]  ( .D(
        \fpu_div_frac_dp/i_dstg_xtra_regs/N9 ), .CLK(n1920), .Q(n1398), .QN(
        \fpu_div_frac_dp/n960 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[52]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N55 ), .CLK(n1921), .Q(n1368) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[51]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N54 ), .CLK(n1921), .Q(n1524) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[50]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N53 ), .CLK(n1921), .Q(n1389) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[49]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N52 ), .CLK(n1921), .Q(n1677) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[48]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N51 ), .CLK(n1921), .Q(n1403) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[47]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N50 ), .CLK(n1922), .Q(n1634) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[46]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N49 ), .CLK(n1922), .Q(n1684), .QN(
        \fpu_div_frac_dp/n343 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[45]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N48 ), .CLK(n1922), .Q(
        \fpu_div_frac_dp/div_norm_inv[45] ), .QN(\fpu_div_frac_dp/n344 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[44]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N47 ), .CLK(n1922), .Q(n1410), .QN(
        \fpu_div_frac_dp/n345 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[43]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N46 ), .CLK(n1922), .Q(
        \fpu_div_frac_dp/div_norm_inv[43] ), .QN(\fpu_div_frac_dp/n984 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[42]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N45 ), .CLK(n1922), .Q(n1633) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[41]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N44 ), .CLK(n1923), .Q(
        \fpu_div_frac_dp/div_norm_inv[41] ), .QN(\fpu_div_frac_dp/n347 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[40]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N43 ), .CLK(n1923), .Q(n1400) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[39]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N42 ), .CLK(n1923), .Q(n1577) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[38]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N41 ), .CLK(n1923), .Q(n1685), .QN(
        \fpu_div_frac_dp/n349 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[37]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N40 ), .CLK(n1923), .Q(
        \fpu_div_frac_dp/div_norm_inv[37] ), .QN(\fpu_div_frac_dp/n350 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[36]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N39 ), .CLK(n1923), .Q(n1367) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[35]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N38 ), .CLK(n1924), .Q(n1525) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[34]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N37 ), .CLK(n1924), .Q(n1390) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[33]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N36 ), .CLK(n1924), .Q(n1678) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[32]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N35 ), .CLK(n1924), .Q(
        \fpu_div_frac_dp/div_norm_inv[32] ), .QN(\fpu_div_frac_dp/n354 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[31]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N34 ), .CLK(n1924), .Q(n1388) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[30]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N33 ), .CLK(n1924), .Q(n1492) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[29]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N32 ), .CLK(n1925), .Q(n1680) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[28]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N31 ), .CLK(n1926), .Q(n1438) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[27]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N30 ), .CLK(n1926), .Q(n1597), .QN(
        \fpu_div_frac_dp/n981 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[26]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N29 ), .CLK(n1926), .Q(
        \fpu_div_frac_dp/div_norm_inv[26] ), .QN(\fpu_div_frac_dp/n358 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[25]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N28 ), .CLK(n1926), .Q(
        \fpu_div_frac_dp/div_norm_inv[25] ), .QN(\fpu_div_frac_dp/n359 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[24]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N27 ), .CLK(n1926), .Q(n1649), .QN(
        \fpu_div_frac_dp/n360 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[23]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N26 ), .CLK(n1927), .Q(
        \fpu_div_frac_dp/div_norm_inv[23] ), .QN(\fpu_div_frac_dp/n2330 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[22]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N25 ), .CLK(n1927), .Q(n1681), .QN(
        \fpu_div_frac_dp/n361 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[21]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N24 ), .CLK(n1927), .Q(
        \fpu_div_frac_dp/div_norm_inv[21] ), .QN(\fpu_div_frac_dp/n362 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[20]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N23 ), .CLK(n1927), .Q(n1386), .QN(
        \fpu_div_frac_dp/n363 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[19]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N22 ), .CLK(n1927), .Q(n1360), .QN(
        \fpu_div_frac_dp/n989 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[18]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N21 ), .CLK(n1927), .Q(n1535), .QN(
        \fpu_div_frac_dp/n364 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[17]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N20 ), .CLK(n1928), .Q(n1675) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[16]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N19 ), .CLK(n1903), .Q(n1408), .QN(
        \fpu_div_frac_dp/n366 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[15]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N18 ), .CLK(n1905), .Q(n1580), .QN(
        \fpu_div_frac_dp/n982 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[14]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N17 ), .CLK(n1907), .Q(
        \fpu_div_frac_dp/div_norm_inv[14] ), .QN(\fpu_div_frac_dp/n367 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[13]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N16 ), .CLK(n1909), .Q(
        \fpu_div_frac_dp/div_norm_inv[13] ), .QN(\fpu_div_frac_dp/n368 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[12]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N15 ), .CLK(n1911), .Q(n1576) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[11]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N14 ), .CLK(n1915), .Q(n1531), .QN(
        \fpu_div_frac_dp/n988 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[10]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N13 ), .CLK(n1912), .Q(n1374) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[9]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N12 ), .CLK(n1902), .Q(n1650), .QN(
        \fpu_div_frac_dp/n371 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[8]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N11 ), .CLK(n1917), .Q(n1674), .QN(
        \fpu_div_frac_dp/n372 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[7]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N10 ), .CLK(n1918), .Q(n1528), .QN(
        \fpu_div_frac_dp/n983 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[6]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N9 ), .CLK(n1925), .Q(
        \fpu_div_frac_dp/div_norm_inv[6] ), .QN(\fpu_div_frac_dp/n373 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[5]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N8 ), .CLK(n1925), .Q(
        \fpu_div_frac_dp/div_norm_inv[5] ), .QN(\fpu_div_frac_dp/n374 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[4]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N7 ), .CLK(n1925), .Q(n1387), .QN(
        \fpu_div_frac_dp/n2333 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[3]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N6 ), .CLK(n1925), .Q(n1369) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[2]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N5 ), .CLK(n1925), .Q(n1673), .QN(
        \fpu_div_frac_dp/n996 ) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[1]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N4 ), .CLK(n1926), .Q(n1499) );
  DFFX1 \fpu_div_frac_dp/i_div_norm_inv/q_reg[0]  ( .D(
        \fpu_div_frac_dp/i_div_norm_inv/N3 ), .CLK(n1921), .Q(
        \fpu_div_frac_dp/div_norm_inv[0] ), .QN(\fpu_div_frac_dp/n377 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[54]  ( .D(
        \fpu_div_frac_dp/n1330 ), .CLK(\fpu_div_frac_dp/n985 ), .Q(n1807), 
        .QN(\fpu_div_frac_dp/n378 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[53]  ( .D(
        \fpu_div_frac_dp/n1331 ), .CLK(\fpu_div_frac_dp/n985 ), .Q(n1849), 
        .QN(\fpu_div_frac_dp/n379 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[52]  ( .D(
        \fpu_div_frac_dp/n1332 ), .CLK(\fpu_div_frac_dp/n985 ), .Q(n1845), 
        .QN(\fpu_div_frac_dp/n380 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[51]  ( .D(
        \fpu_div_frac_dp/n1333 ), .CLK(\fpu_div_frac_dp/n985 ), .Q(n1671), 
        .QN(\fpu_div_frac_dp/n381 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[50]  ( .D(
        \fpu_div_frac_dp/n1334 ), .CLK(\fpu_div_frac_dp/n985 ), .Q(n1806), 
        .QN(\fpu_div_frac_dp/n382 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[49]  ( .D(
        \fpu_div_frac_dp/n1335 ), .CLK(\fpu_div_frac_dp/n985 ), .Q(n1653), 
        .QN(\fpu_div_frac_dp/n383 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[48]  ( .D(
        \fpu_div_frac_dp/n1336 ), .CLK(n1900), .Q(n1654), .QN(
        \fpu_div_frac_dp/n384 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[47]  ( .D(
        \fpu_div_frac_dp/n1337 ), .CLK(n1901), .Q(n1655), .QN(
        \fpu_div_frac_dp/n385 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[46]  ( .D(
        \fpu_div_frac_dp/n1338 ), .CLK(n1925), .Q(n1656), .QN(
        \fpu_div_frac_dp/n386 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[45]  ( .D(
        \fpu_div_frac_dp/n1339 ), .CLK(n1927), .Q(n1657), .QN(
        \fpu_div_frac_dp/n387 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[44]  ( .D(
        \fpu_div_frac_dp/n1340 ), .CLK(n1926), .Q(n1658), .QN(
        \fpu_div_frac_dp/n388 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[43]  ( .D(
        \fpu_div_frac_dp/n1341 ), .CLK(n1924), .Q(n1659), .QN(
        \fpu_div_frac_dp/n389 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[42]  ( .D(
        \fpu_div_frac_dp/n1342 ), .CLK(n1923), .Q(n1660), .QN(
        \fpu_div_frac_dp/n390 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[41]  ( .D(
        \fpu_div_frac_dp/n1343 ), .CLK(n1935), .Q(n1661), .QN(
        \fpu_div_frac_dp/n391 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[40]  ( .D(
        \fpu_div_frac_dp/n1344 ), .CLK(n1935), .Q(n1662), .QN(
        \fpu_div_frac_dp/n392 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[39]  ( .D(
        \fpu_div_frac_dp/n1345 ), .CLK(n1935), .Q(n1663), .QN(
        \fpu_div_frac_dp/n393 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[38]  ( .D(
        \fpu_div_frac_dp/n1346 ), .CLK(n1935), .Q(n1664), .QN(
        \fpu_div_frac_dp/n394 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[37]  ( .D(
        \fpu_div_frac_dp/n1347 ), .CLK(n1935), .Q(n1665), .QN(
        \fpu_div_frac_dp/n395 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[36]  ( .D(
        \fpu_div_frac_dp/n1348 ), .CLK(n1935), .Q(n1666), .QN(
        \fpu_div_frac_dp/n396 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[35]  ( .D(
        \fpu_div_frac_dp/n1349 ), .CLK(n1935), .Q(n1667), .QN(
        \fpu_div_frac_dp/n397 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[34]  ( .D(
        \fpu_div_frac_dp/n1350 ), .CLK(n1935), .Q(n1668), .QN(
        \fpu_div_frac_dp/n398 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[33]  ( .D(
        \fpu_div_frac_dp/n1351 ), .CLK(n1935), .Q(n1669), .QN(
        \fpu_div_frac_dp/n399 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[32]  ( .D(
        \fpu_div_frac_dp/n1352 ), .CLK(n1935), .Q(n1652), .QN(
        \fpu_div_frac_dp/n400 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[31]  ( .D(
        \fpu_div_frac_dp/n1353 ), .CLK(n1935), .Q(n1711), .QN(
        \fpu_div_frac_dp/n401 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[30]  ( .D(
        \fpu_div_frac_dp/n1354 ), .CLK(n1935), .Q(n1712), .QN(
        \fpu_div_frac_dp/n402 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[29]  ( .D(
        \fpu_div_frac_dp/n1355 ), .CLK(n1934), .Q(n1714), .QN(
        \fpu_div_frac_dp/n403 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[28]  ( .D(
        \fpu_div_frac_dp/n1356 ), .CLK(n1934), .Q(n1713), .QN(
        \fpu_div_frac_dp/n404 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[27]  ( .D(
        \fpu_div_frac_dp/n1357 ), .CLK(n1934), .Q(n1692), .QN(
        \fpu_div_frac_dp/n405 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[26]  ( .D(
        \fpu_div_frac_dp/n1358 ), .CLK(n1934), .Q(n1693), .QN(
        \fpu_div_frac_dp/n406 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[25]  ( .D(
        \fpu_div_frac_dp/n1359 ), .CLK(n1934), .Q(n1694), .QN(
        \fpu_div_frac_dp/n407 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[24]  ( .D(
        \fpu_div_frac_dp/n1360 ), .CLK(n1934), .Q(n1695), .QN(
        \fpu_div_frac_dp/n408 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[23]  ( .D(
        \fpu_div_frac_dp/n1361 ), .CLK(n1934), .Q(n1696), .QN(
        \fpu_div_frac_dp/n409 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[22]  ( .D(
        \fpu_div_frac_dp/n1362 ), .CLK(n1934), .Q(n1697), .QN(
        \fpu_div_frac_dp/n410 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[21]  ( .D(
        \fpu_div_frac_dp/n1363 ), .CLK(n1934), .Q(n1698), .QN(
        \fpu_div_frac_dp/n411 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[20]  ( .D(
        \fpu_div_frac_dp/n1364 ), .CLK(n1934), .Q(n1699), .QN(
        \fpu_div_frac_dp/n412 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[19]  ( .D(
        \fpu_div_frac_dp/n1365 ), .CLK(n1934), .Q(n1700), .QN(
        \fpu_div_frac_dp/n413 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[18]  ( .D(
        \fpu_div_frac_dp/n1366 ), .CLK(n1934), .Q(n1701), .QN(
        \fpu_div_frac_dp/n414 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[17]  ( .D(
        \fpu_div_frac_dp/n1367 ), .CLK(n1933), .Q(n1702), .QN(
        \fpu_div_frac_dp/n415 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[16]  ( .D(
        \fpu_div_frac_dp/n1368 ), .CLK(n1933), .Q(n1703), .QN(
        \fpu_div_frac_dp/n416 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[15]  ( .D(
        \fpu_div_frac_dp/n1369 ), .CLK(n1933), .Q(n1704), .QN(
        \fpu_div_frac_dp/n417 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[14]  ( .D(
        \fpu_div_frac_dp/n1370 ), .CLK(n1933), .Q(n1705), .QN(
        \fpu_div_frac_dp/n418 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[13]  ( .D(
        \fpu_div_frac_dp/n1371 ), .CLK(n1933), .Q(n1706), .QN(
        \fpu_div_frac_dp/n419 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[12]  ( .D(
        \fpu_div_frac_dp/n1372 ), .CLK(n1933), .Q(n1707), .QN(
        \fpu_div_frac_dp/n420 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[11]  ( .D(
        \fpu_div_frac_dp/n1373 ), .CLK(n1933), .Q(n1708), .QN(
        \fpu_div_frac_dp/n421 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[10]  ( .D(
        \fpu_div_frac_dp/n1374 ), .CLK(n1933), .Q(n1818), .QN(
        \fpu_div_frac_dp/n422 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[9]  ( .D(\fpu_div_frac_dp/n1375 ), .CLK(n1933), .Q(n1639) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[8]  ( .D(\fpu_div_frac_dp/n1376 ), .CLK(n1933), .Q(n1709), .QN(\fpu_div_frac_dp/n424 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[7]  ( .D(\fpu_div_frac_dp/n1377 ), .CLK(n1933), .Q(n1710), .QN(\fpu_div_frac_dp/n425 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[6]  ( .D(\fpu_div_frac_dp/n1378 ), .CLK(n1933), .Q(n1686), .QN(\fpu_div_frac_dp/n426 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[5]  ( .D(\fpu_div_frac_dp/n1379 ), .CLK(n1932), .Q(n1687), .QN(\fpu_div_frac_dp/n427 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[4]  ( .D(\fpu_div_frac_dp/n1380 ), .CLK(n1932), .Q(n1688), .QN(\fpu_div_frac_dp/n428 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[3]  ( .D(\fpu_div_frac_dp/n1381 ), .CLK(n1932), .Q(n1689), .QN(\fpu_div_frac_dp/n429 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[2]  ( .D(\fpu_div_frac_dp/n1382 ), .CLK(n1932), .Q(n1690), .QN(\fpu_div_frac_dp/n430 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[1]  ( .D(\fpu_div_frac_dp/n1383 ), .CLK(n1932), .Q(n1691), .QN(\fpu_div_frac_dp/n431 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in2/q_reg[0]  ( .D(\fpu_div_frac_dp/n1384 ), .CLK(n1932), .Q(n1816), .QN(\fpu_div_frac_dp/n432 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[54]  ( .D(
        \fpu_div_frac_dp/n1385 ), .CLK(n1932), .Q(n1850), .QN(
        \fpu_div_frac_dp/n433 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[53]  ( .D(
        \fpu_div_frac_dp/n1386 ), .CLK(n1932), .Q(n1847), .QN(
        \fpu_div_frac_dp/n434 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[52]  ( .D(
        \fpu_div_frac_dp/n1387 ), .CLK(n1932), .Q(n1811), .QN(
        \fpu_div_frac_dp/n435 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[51]  ( .D(
        \fpu_div_frac_dp/n1388 ), .CLK(n1932), .Q(n1670), .QN(
        \fpu_div_frac_dp/n436 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[50]  ( .D(
        \fpu_div_frac_dp/n1389 ), .CLK(n1932), .Q(n1805), .QN(
        \fpu_div_frac_dp/n437 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[49]  ( .D(
        \fpu_div_frac_dp/n1390 ), .CLK(n1932), .Q(n1803), .QN(
        \fpu_div_frac_dp/n438 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[48]  ( .D(
        \fpu_div_frac_dp/n1391 ), .CLK(n1931), .Q(n1802), .QN(
        \fpu_div_frac_dp/n439 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[47]  ( .D(
        \fpu_div_frac_dp/n1392 ), .CLK(n1931), .Q(n1801), .QN(
        \fpu_div_frac_dp/n440 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[46]  ( .D(
        \fpu_div_frac_dp/n1393 ), .CLK(n1931), .Q(n1800), .QN(
        \fpu_div_frac_dp/n441 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[45]  ( .D(
        \fpu_div_frac_dp/n1394 ), .CLK(n1931), .Q(n1799), .QN(
        \fpu_div_frac_dp/n442 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[44]  ( .D(
        \fpu_div_frac_dp/n1395 ), .CLK(n1931), .Q(n1798), .QN(
        \fpu_div_frac_dp/n443 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[43]  ( .D(
        \fpu_div_frac_dp/n1396 ), .CLK(n1931), .Q(n1797), .QN(
        \fpu_div_frac_dp/n444 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[42]  ( .D(
        \fpu_div_frac_dp/n1397 ), .CLK(n1931), .Q(n1796), .QN(
        \fpu_div_frac_dp/n445 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[41]  ( .D(
        \fpu_div_frac_dp/n1398 ), .CLK(n1931), .Q(n1795), .QN(
        \fpu_div_frac_dp/n446 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[40]  ( .D(
        \fpu_div_frac_dp/n1399 ), .CLK(n1931), .Q(n1794), .QN(
        \fpu_div_frac_dp/n447 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[39]  ( .D(
        \fpu_div_frac_dp/n1400 ), .CLK(n1931), .Q(n1793), .QN(
        \fpu_div_frac_dp/n448 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[38]  ( .D(
        \fpu_div_frac_dp/n1401 ), .CLK(n1931), .Q(n1792), .QN(
        \fpu_div_frac_dp/n449 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[37]  ( .D(
        \fpu_div_frac_dp/n1402 ), .CLK(n1931), .Q(n1791), .QN(
        \fpu_div_frac_dp/n450 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[36]  ( .D(
        \fpu_div_frac_dp/n1403 ), .CLK(n1930), .Q(n1790), .QN(
        \fpu_div_frac_dp/n451 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[35]  ( .D(
        \fpu_div_frac_dp/n1404 ), .CLK(n1930), .Q(n1789), .QN(
        \fpu_div_frac_dp/n452 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[34]  ( .D(
        \fpu_div_frac_dp/n1405 ), .CLK(n1930), .Q(n1788), .QN(
        \fpu_div_frac_dp/n453 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[33]  ( .D(
        \fpu_div_frac_dp/n1406 ), .CLK(n1930), .Q(n1787), .QN(
        \fpu_div_frac_dp/n454 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[32]  ( .D(
        \fpu_div_frac_dp/n1407 ), .CLK(n1930), .Q(n1804), .QN(
        \fpu_div_frac_dp/n455 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[31]  ( .D(
        \fpu_div_frac_dp/n1408 ), .CLK(n1930), .Q(n1813), .QN(
        \fpu_div_frac_dp/n456 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[30]  ( .D(
        \fpu_div_frac_dp/n1409 ), .CLK(n1930), .Q(n1812), .QN(
        \fpu_div_frac_dp/n457 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[29]  ( .D(
        \fpu_div_frac_dp/n1410 ), .CLK(n1930), .Q(n1810), .QN(
        \fpu_div_frac_dp/n458 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[28]  ( .D(
        \fpu_div_frac_dp/n1411 ), .CLK(n1930), .Q(n1814), .QN(
        \fpu_div_frac_dp/n459 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[27]  ( .D(
        \fpu_div_frac_dp/n1412 ), .CLK(n1930), .Q(n1844), .QN(
        \fpu_div_frac_dp/n460 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[26]  ( .D(
        \fpu_div_frac_dp/n1413 ), .CLK(n1930), .Q(n1843), .QN(
        \fpu_div_frac_dp/n461 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[25]  ( .D(
        \fpu_div_frac_dp/n1414 ), .CLK(n1930), .Q(n1842), .QN(
        \fpu_div_frac_dp/n462 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[24]  ( .D(
        \fpu_div_frac_dp/n1415 ), .CLK(n1929), .Q(n1841), .QN(
        \fpu_div_frac_dp/n463 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[23]  ( .D(
        \fpu_div_frac_dp/n1416 ), .CLK(n1929), .Q(n1840), .QN(
        \fpu_div_frac_dp/n464 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[22]  ( .D(
        \fpu_div_frac_dp/n1417 ), .CLK(n1929), .Q(n1839), .QN(
        \fpu_div_frac_dp/n465 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[21]  ( .D(
        \fpu_div_frac_dp/n1418 ), .CLK(n1929), .Q(n1838), .QN(
        \fpu_div_frac_dp/n466 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[20]  ( .D(
        \fpu_div_frac_dp/n1419 ), .CLK(n1929), .Q(n1837), .QN(
        \fpu_div_frac_dp/n467 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[19]  ( .D(
        \fpu_div_frac_dp/n1420 ), .CLK(n1929), .Q(n1836), .QN(
        \fpu_div_frac_dp/n468 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[18]  ( .D(
        \fpu_div_frac_dp/n1421 ), .CLK(n1929), .Q(n1835), .QN(
        \fpu_div_frac_dp/n469 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[17]  ( .D(
        \fpu_div_frac_dp/n1422 ), .CLK(n1929), .Q(n1834), .QN(
        \fpu_div_frac_dp/n470 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[16]  ( .D(
        \fpu_div_frac_dp/n1423 ), .CLK(n1929), .Q(n1833), .QN(
        \fpu_div_frac_dp/n471 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[15]  ( .D(
        \fpu_div_frac_dp/n1424 ), .CLK(n1929), .Q(n1832), .QN(
        \fpu_div_frac_dp/n472 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[14]  ( .D(
        \fpu_div_frac_dp/n1425 ), .CLK(n1929), .Q(n1831), .QN(
        \fpu_div_frac_dp/n473 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[13]  ( .D(
        \fpu_div_frac_dp/n1426 ), .CLK(n1929), .Q(n1830), .QN(
        \fpu_div_frac_dp/n474 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[12]  ( .D(
        \fpu_div_frac_dp/n1427 ), .CLK(n1928), .Q(n1829), .QN(
        \fpu_div_frac_dp/n475 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[11]  ( .D(
        \fpu_div_frac_dp/n1428 ), .CLK(n1928), .Q(n1828), .QN(
        \fpu_div_frac_dp/n476 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[10]  ( .D(
        \fpu_div_frac_dp/n1429 ), .CLK(n1928), .Q(n1846), .QN(
        \fpu_div_frac_dp/n477 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[9]  ( .D(\fpu_div_frac_dp/n1430 ), .CLK(n1928), .Q(n1848), .QN(\fpu_div_frac_dp/n478 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[8]  ( .D(\fpu_div_frac_dp/n1431 ), .CLK(n1928), .Q(n1827), .QN(\fpu_div_frac_dp/n479 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[7]  ( .D(\fpu_div_frac_dp/n1432 ), .CLK(n1928), .Q(n1826), .QN(\fpu_div_frac_dp/n480 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[6]  ( .D(\fpu_div_frac_dp/n1433 ), .CLK(n1928), .Q(n1825), .QN(\fpu_div_frac_dp/n481 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[5]  ( .D(\fpu_div_frac_dp/n1434 ), .CLK(n1928), .Q(n1824), .QN(\fpu_div_frac_dp/n482 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[4]  ( .D(\fpu_div_frac_dp/n1435 ), .CLK(n1928), .Q(n1823), .QN(\fpu_div_frac_dp/n483 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[3]  ( .D(\fpu_div_frac_dp/n1436 ), .CLK(n1928), .Q(n1822), .QN(\fpu_div_frac_dp/n484 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[2]  ( .D(\fpu_div_frac_dp/n1437 ), .CLK(n1928), .Q(n1821), .QN(\fpu_div_frac_dp/n485 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[1]  ( .D(\fpu_div_frac_dp/n1438 ), .CLK(n1928), .Q(n1820), .QN(\fpu_div_frac_dp/n486 ) );
  DFFX1 \fpu_div_frac_dp/i_div_frac_in1/q_reg[0]  ( .D(\fpu_div_frac_dp/n1439 ), .CLK(n1922), .Q(n1819), .QN(\fpu_div_frac_dp/n487 ) );
  LATCHX1 \fpu_div_frac_dp/ckbuf_div_frac_dp/clken_reg  ( .CLK(
        \fpu_div_frac_dp/rclk ), .D(\fpu_div_frac_dp/ckbuf_div_frac_dp/N1 ), 
        .QN(\fpu_div_frac_dp/n168 ) );
  OR2X1 U1129 ( .IN1(n1888), .IN2(se), .Q(n1548) );
  OR2X1 U1130 ( .IN1(n185), .IN2(se), .Q(n1550) );
  INVX0 U1131 ( .INP(n1548), .ZN(n1879) );
  INVX0 U1132 ( .INP(n1548), .ZN(n1880) );
  INVX0 U1133 ( .INP(n1548), .ZN(n1881) );
  INVX0 U1134 ( .INP(n1548), .ZN(n1882) );
  INVX0 U1135 ( .INP(n1550), .ZN(n1883) );
  INVX0 U1136 ( .INP(n1550), .ZN(n1884) );
  INVX0 U1137 ( .INP(n1550), .ZN(n1885) );
  INVX0 U1138 ( .INP(n1550), .ZN(n1886) );
  INVX2 U1139 ( .INP(n2633), .ZN(n2560) );
  INVX2 U1140 ( .INP(n2628), .ZN(n2566) );
  INVX0 U1141 ( .INP(n1936), .ZN(n1928) );
  INVX0 U1142 ( .INP(n1936), .ZN(n1929) );
  INVX0 U1143 ( .INP(n1936), .ZN(n1930) );
  INVX0 U1144 ( .INP(n1936), .ZN(n1931) );
  INVX0 U1145 ( .INP(n1936), .ZN(n1932) );
  INVX0 U1146 ( .INP(n1936), .ZN(n1933) );
  INVX0 U1147 ( .INP(n1936), .ZN(n1934) );
  INVX0 U1148 ( .INP(n1936), .ZN(n1935) );
  INVX0 U1149 ( .INP(n1937), .ZN(n1925) );
  INVX0 U1150 ( .INP(n1937), .ZN(n1927) );
  INVX0 U1151 ( .INP(n1937), .ZN(n1926) );
  INVX0 U1152 ( .INP(n1937), .ZN(n1924) );
  INVX0 U1153 ( .INP(n1937), .ZN(n1923) );
  INVX0 U1154 ( .INP(n1937), .ZN(n1922) );
  INVX0 U1155 ( .INP(n1937), .ZN(n1921) );
  INVX0 U1156 ( .INP(n1937), .ZN(n1920) );
  INVX0 U1157 ( .INP(n1938), .ZN(n1912) );
  INVX0 U1158 ( .INP(n1937), .ZN(n1918) );
  INVX0 U1159 ( .INP(n1938), .ZN(n1914) );
  INVX0 U1160 ( .INP(n1937), .ZN(n1916) );
  INVX0 U1161 ( .INP(n1938), .ZN(n1915) );
  INVX0 U1162 ( .INP(n1938), .ZN(n1913) );
  INVX0 U1163 ( .INP(n1937), .ZN(n1917) );
  INVX0 U1164 ( .INP(n1937), .ZN(n1919) );
  INVX0 U1165 ( .INP(n1938), .ZN(n1911) );
  INVX0 U1166 ( .INP(n1938), .ZN(n1910) );
  INVX0 U1167 ( .INP(n1938), .ZN(n1909) );
  INVX0 U1168 ( .INP(n1938), .ZN(n1908) );
  INVX0 U1169 ( .INP(n1938), .ZN(n1907) );
  INVX0 U1170 ( .INP(n1938), .ZN(n1906) );
  INVX0 U1171 ( .INP(n1938), .ZN(n1905) );
  INVX0 U1172 ( .INP(n1938), .ZN(n1904) );
  INVX0 U1173 ( .INP(n1937), .ZN(n1900) );
  INVX0 U1174 ( .INP(n1936), .ZN(n1903) );
  INVX0 U1175 ( .INP(n1938), .ZN(n1902) );
  INVX0 U1176 ( .INP(n1937), .ZN(n1901) );
  INVX0 U1177 ( .INP(n1936), .ZN(n1898) );
  INVX0 U1178 ( .INP(n1938), .ZN(n1899) );
  INVX0 U1179 ( .INP(n1887), .ZN(n1896) );
  INVX0 U1180 ( .INP(n1887), .ZN(n1895) );
  INVX0 U1181 ( .INP(n1887), .ZN(n1888) );
  INVX0 U1182 ( .INP(n1887), .ZN(n1889) );
  INVX0 U1183 ( .INP(n1887), .ZN(n1890) );
  INVX0 U1184 ( .INP(n1887), .ZN(n1892) );
  INVX0 U1185 ( .INP(n1887), .ZN(n1891) );
  INVX0 U1186 ( .INP(n1887), .ZN(n1893) );
  INVX0 U1187 ( .INP(n1887), .ZN(n1894) );
  INVX0 U1188 ( .INP(n1887), .ZN(n1897) );
  INVX0 U1189 ( .INP(\fpu_div_frac_dp/n985 ), .ZN(n1937) );
  INVX0 U1190 ( .INP(\fpu_div_frac_dp/n985 ), .ZN(n1936) );
  INVX0 U1191 ( .INP(\fpu_div_frac_dp/n985 ), .ZN(n1938) );
  OR2X1 U1192 ( .IN1(\fpu_div_frac_dp/d1stg_step ), .IN2(se), .Q(n1887) );
  NOR2X0 U1193 ( .IN1(n151), .IN2(\fpu_div_frac_dp/rclk ), .QN(n577) );
  OAI22X1 U1194 ( .IN1(n1939), .IN2(n1940), .IN3(n1941), .IN4(n613), .QN(n515)
         );
  AO22X1 U1195 ( .IN1(n1942), .IN2(n1782), .IN3(n1943), .IN4(n1944), .Q(n514)
         );
  XNOR3X1 U1196 ( .IN1(n1945), .IN2(n1946), .IN3(n1947), .Q(n1943) );
  OR2X1 U1197 ( .IN1(n117), .IN2(n607), .Q(n1947) );
  OA22X1 U1198 ( .IN1(n1948), .IN2(n1949), .IN3(n1950), .IN4(n1946), .Q(n1945)
         );
  NOR2X0 U1199 ( .IN1(n1951), .IN2(n1952), .QN(n1949) );
  AO22X1 U1200 ( .IN1(n1953), .IN2(n1954), .IN3(n1955), .IN4(n1856), .Q(n513)
         );
  AO21X1 U1201 ( .IN1(n1956), .IN2(n1538), .IN3(n1957), .Q(n511) );
  AO21X1 U1202 ( .IN1(n1956), .IN2(n1401), .IN3(n1957), .Q(n510) );
  AO21X1 U1203 ( .IN1(n1956), .IN2(n1376), .IN3(n1957), .Q(n509) );
  AO21X1 U1204 ( .IN1(n1956), .IN2(n1643), .IN3(n1957), .Q(n508) );
  AO21X1 U1205 ( .IN1(n1956), .IN2(n1870), .IN3(n1958), .Q(n507) );
  AO21X1 U1206 ( .IN1(n1956), .IN2(n1731), .IN3(n1958), .Q(n505) );
  AO21X1 U1207 ( .IN1(n1956), .IN2(n1547), .IN3(n1958), .Q(n504) );
  AO21X1 U1208 ( .IN1(n1956), .IN2(n1375), .IN3(n1958), .Q(n503) );
  AO21X1 U1209 ( .IN1(n1956), .IN2(n1720), .IN3(n1958), .Q(n502) );
  AO22X1 U1210 ( .IN1(n1956), .IN2(n1875), .IN3(inq_rnd_mode[1]), .IN4(n1959), 
        .Q(n501) );
  AO22X1 U1211 ( .IN1(n1956), .IN2(n1732), .IN3(inq_rnd_mode[0]), .IN4(n1959), 
        .Q(n500) );
  AO22X1 U1212 ( .IN1(n1956), .IN2(n1786), .IN3(inq_id[4]), .IN4(n1959), .Q(
        n499) );
  AO22X1 U1213 ( .IN1(n1956), .IN2(n1551), .IN3(inq_id[3]), .IN4(n1959), .Q(
        n498) );
  AO22X1 U1214 ( .IN1(n1956), .IN2(n1715), .IN3(inq_id[2]), .IN4(n1959), .Q(
        n497) );
  AO22X1 U1215 ( .IN1(n1956), .IN2(n1722), .IN3(inq_id[1]), .IN4(n1959), .Q(
        n496) );
  AO22X1 U1216 ( .IN1(n1956), .IN2(n1723), .IN3(inq_id[0]), .IN4(n1959), .Q(
        n495) );
  AO22X1 U1217 ( .IN1(n1956), .IN2(n1641), .IN3(inq_in1[63]), .IN4(n1959), .Q(
        n494) );
  AO22X1 U1218 ( .IN1(n1956), .IN2(n1539), .IN3(inq_in2[63]), .IN4(n1959), .Q(
        n493) );
  AO22X1 U1219 ( .IN1(n1942), .IN2(n1815), .IN3(n1960), .IN4(n1944), .Q(n492)
         );
  XNOR3X1 U1220 ( .IN1(n1961), .IN2(n1962), .IN3(n1963), .Q(n1960) );
  AO22X1 U1221 ( .IN1(n1942), .IN2(n1817), .IN3(n1944), .IN4(n1964), .Q(n491)
         );
  XOR3X1 U1222 ( .IN1(n1965), .IN2(n1966), .IN3(n1967), .Q(n1964) );
  AO22X1 U1223 ( .IN1(n1942), .IN2(n1809), .IN3(n1968), .IN4(n1944), .Q(n490)
         );
  XOR3X1 U1224 ( .IN1(n1969), .IN2(n1970), .IN3(n1971), .Q(n1968) );
  AO22X1 U1225 ( .IN1(n1942), .IN2(n1808), .IN3(n1972), .IN4(n1944), .Q(n489)
         );
  XOR3X1 U1226 ( .IN1(n1973), .IN2(n1974), .IN3(n1975), .Q(n1972) );
  AO222X1 U1227 ( .IN1(n1976), .IN2(n1944), .IN3(n291), .IN4(n1977), .IN5(
        n1942), .IN6(n1409), .Q(n488) );
  NAND2X0 U1228 ( .IN1(n181), .IN2(n182), .QN(n1977) );
  XNOR3X1 U1229 ( .IN1(n1978), .IN2(n1979), .IN3(n1980), .Q(n1976) );
  AO22X1 U1230 ( .IN1(n1942), .IN2(n1575), .IN3(n1944), .IN4(n1981), .Q(n487)
         );
  XOR3X1 U1231 ( .IN1(n1982), .IN2(n1983), .IN3(n1984), .Q(n1981) );
  INVX0 U1232 ( .INP(n1985), .ZN(n1944) );
  AO22X1 U1233 ( .IN1(n1986), .IN2(n1396), .IN3(n1987), .IN4(n1851), .Q(n486)
         );
  AO22X1 U1234 ( .IN1(n1986), .IN2(n1461), .IN3(n1987), .IN4(n1852), .Q(n485)
         );
  MUX21X1 U1235 ( .IN1(n1988), .IN2(n1989), .S(n616), .Q(n484) );
  MUX21X1 U1236 ( .IN1(n1990), .IN2(n1991), .S(n1372), .Q(n483) );
  AO21X1 U1237 ( .IN1(n1989), .IN2(n616), .IN3(n1988), .Q(n1991) );
  NOR2X0 U1238 ( .IN1(n616), .IN2(n1992), .QN(n1990) );
  INVX0 U1239 ( .INP(n1989), .ZN(n1992) );
  AO22X1 U1240 ( .IN1(n1988), .IN2(n1542), .IN3(n1993), .IN4(n1989), .Q(n482)
         );
  AND2X1 U1241 ( .IN1(n1994), .IN2(n1995), .Q(n1993) );
  AO22X1 U1242 ( .IN1(n1988), .IN2(n1395), .IN3(n1996), .IN4(n1989), .Q(n481)
         );
  AO22X1 U1243 ( .IN1(n1988), .IN2(n1541), .IN3(n1989), .IN4(n1997), .Q(n480)
         );
  AO22X1 U1244 ( .IN1(n1988), .IN2(n1545), .IN3(n1989), .IN4(n1998), .Q(n479)
         );
  NOR2X0 U1245 ( .IN1(n1999), .IN2(n2000), .QN(n1989) );
  AND3X1 U1246 ( .IN1(n185), .IN2(n2000), .IN3(n1354), .Q(n1988) );
  OAI22X1 U1247 ( .IN1(n2001), .IN2(n58), .IN3(n2002), .IN4(n59), .QN(n478) );
  AO22X1 U1248 ( .IN1(n593), .IN2(n2003), .IN3(n2004), .IN4(n1732), .Q(n477)
         );
  NOR2X0 U1249 ( .IN1(n1999), .IN2(n2005), .QN(n476) );
  MUX21X1 U1250 ( .IN1(n124), .IN2(n630), .S(n939), .Q(n2005) );
  NOR2X0 U1251 ( .IN1(n1999), .IN2(n2006), .QN(n475) );
  MUX21X1 U1252 ( .IN1(n21), .IN2(n22), .S(n939), .Q(n2006) );
  AO22X1 U1253 ( .IN1(n2007), .IN2(n1783), .IN3(n2008), .IN4(n2009), .Q(n474)
         );
  NOR2X0 U1254 ( .IN1(se), .IN2(n194), .QN(n2008) );
  AO22X1 U1255 ( .IN1(n2010), .IN2(n2011), .IN3(n2012), .IN4(n1536), .Q(n473)
         );
  NAND2X0 U1256 ( .IN1(n2013), .IN2(n2014), .QN(n2011) );
  MUX21X1 U1257 ( .IN1(n2015), .IN2(n2016), .S(n2017), .Q(n2013) );
  NAND2X0 U1258 ( .IN1(n192), .IN2(div_frac_outa[28]), .QN(n2015) );
  AO22X1 U1259 ( .IN1(n2012), .IN2(n1717), .IN3(n2018), .IN4(n2010), .Q(n472)
         );
  MUX21X1 U1260 ( .IN1(n2019), .IN2(n2020), .S(n2017), .Q(n2018) );
  INVX0 U1261 ( .INP(n2016), .ZN(n2019) );
  MUX21X1 U1262 ( .IN1(\fpu_div_frac_dp/n92 ), .IN2(\fpu_div_frac_dp/n6 ), .S(
        n1397), .Q(n2016) );
  NOR2X0 U1263 ( .IN1(se), .IN2(n2021), .QN(n471) );
  MUX21X1 U1264 ( .IN1(n14), .IN2(n2022), .S(n1393), .Q(n2021) );
  AO22X1 U1265 ( .IN1(n2012), .IN2(n1874), .IN3(n2023), .IN4(n2010), .Q(n470)
         );
  MUX21X1 U1266 ( .IN1(n2020), .IN2(n2024), .S(n2017), .Q(n2023) );
  MUX21X1 U1267 ( .IN1(div_frac_outa[31]), .IN2(div_frac_outa[2]), .S(n1397), 
        .Q(n2024) );
  MUX21X1 U1268 ( .IN1(div_frac_outa[1]), .IN2(div_frac_outa[30]), .S(n192), 
        .Q(n2020) );
  NOR2X0 U1269 ( .IN1(n1552), .IN2(se), .QN(n2012) );
  AO22X1 U1270 ( .IN1(n1986), .IN2(n1579), .IN3(n1987), .IN4(n1433), .Q(n469)
         );
  AO22X1 U1271 ( .IN1(n2025), .IN2(n1954), .IN3(n1955), .IN4(n1853), .Q(n468)
         );
  AO22X1 U1272 ( .IN1(n2025), .IN2(n1954), .IN3(n1955), .IN4(n1854), .Q(n467)
         );
  NAND2X0 U1273 ( .IN1(n138), .IN2(n2026), .QN(n2025) );
  NAND4X0 U1274 ( .IN1(n2027), .IN2(n2028), .IN3(n2029), .IN4(n1396), .QN(
        n2026) );
  AO21X1 U1275 ( .IN1(n2030), .IN2(n2031), .IN3(n2032), .Q(n2029) );
  NAND3X0 U1276 ( .IN1(n1994), .IN2(n1372), .IN3(n616), .QN(n2031) );
  AO22X1 U1277 ( .IN1(n1953), .IN2(n1954), .IN3(n1955), .IN4(n1857), .Q(n466)
         );
  AND2X1 U1278 ( .IN1(n1986), .IN2(n2033), .Q(n1955) );
  NOR2X0 U1279 ( .IN1(n1999), .IN2(n272), .QN(n1986) );
  AO21X1 U1280 ( .IN1(n1354), .IN2(n939), .IN3(n1987), .Q(n1954) );
  AND2X1 U1281 ( .IN1(n1354), .IN2(n272), .Q(n1987) );
  NAND2X0 U1282 ( .IN1(n131), .IN2(n2034), .QN(n1953) );
  NAND3X0 U1283 ( .IN1(n2035), .IN2(n1461), .IN3(n2027), .QN(n2034) );
  NAND3X0 U1284 ( .IN1(n1997), .IN2(n2036), .IN3(n1998), .QN(n2035) );
  INVX0 U1285 ( .INP(n2028), .ZN(n1998) );
  XOR2X1 U1286 ( .IN1(n2037), .IN2(n1545), .Q(n2028) );
  NAND2X0 U1287 ( .IN1(n2038), .IN2(n1541), .QN(n2037) );
  AO21X1 U1288 ( .IN1(n1995), .IN2(n1994), .IN3(n1996), .Q(n2036) );
  INVX0 U1289 ( .INP(n2030), .ZN(n1996) );
  AO21X1 U1290 ( .IN1(n586), .IN2(n1995), .IN3(n2038), .Q(n2030) );
  OR2X1 U1291 ( .IN1(n1542), .IN2(n2039), .Q(n1994) );
  INVX0 U1292 ( .INP(n2032), .ZN(n1997) );
  XOR2X1 U1293 ( .IN1(n602), .IN2(n2038), .Q(n2032) );
  NOR2X0 U1294 ( .IN1(n1995), .IN2(n586), .QN(n2038) );
  NAND2X0 U1295 ( .IN1(n2039), .IN2(n1542), .QN(n1995) );
  NOR2X0 U1296 ( .IN1(n616), .IN2(n594), .QN(n2039) );
  AO22X1 U1297 ( .IN1(n1895), .IN2(n1672), .IN3(inq_in1[51]), .IN4(n2040), .Q(
        n465) );
  AO22X1 U1298 ( .IN1(n1897), .IN2(n1648), .IN3(inq_in1[54]), .IN4(n2040), .Q(
        n464) );
  AO22X1 U1299 ( .IN1(n1897), .IN2(n1868), .IN3(inq_in1_53_0_neq_0), .IN4(
        n2040), .Q(n463) );
  AO22X1 U1300 ( .IN1(n1896), .IN2(n1489), .IN3(inq_in1_50_0_neq_0), .IN4(
        n2040), .Q(n462) );
  AO22X1 U1301 ( .IN1(n1897), .IN2(n1490), .IN3(inq_in1_53_32_neq_0), .IN4(
        n2040), .Q(n461) );
  AO22X1 U1302 ( .IN1(n604), .IN2(n1897), .IN3(inq_in1_exp_eq_0), .IN4(n2040), 
        .Q(n460) );
  AO22X1 U1303 ( .IN1(n1896), .IN2(n1543), .IN3(inq_in1_exp_neq_ffs), .IN4(
        n2040), .Q(n459) );
  AO22X1 U1304 ( .IN1(n1897), .IN2(n1651), .IN3(inq_in2[51]), .IN4(n2040), .Q(
        n458) );
  AO22X1 U1305 ( .IN1(n1896), .IN2(n1645), .IN3(inq_in2[54]), .IN4(n2040), .Q(
        n457) );
  AO22X1 U1306 ( .IN1(n1896), .IN2(n1869), .IN3(inq_in2_53_0_neq_0), .IN4(
        n2040), .Q(n456) );
  AO22X1 U1307 ( .IN1(n1896), .IN2(n1682), .IN3(inq_in2_50_0_neq_0), .IN4(
        n2040), .Q(n455) );
  AO22X1 U1308 ( .IN1(n1896), .IN2(n1679), .IN3(inq_in2_53_32_neq_0), .IN4(
        n2040), .Q(n454) );
  AO22X1 U1309 ( .IN1(n606), .IN2(n1897), .IN3(inq_in2_exp_eq_0), .IN4(n2040), 
        .Q(n453) );
  AO22X1 U1310 ( .IN1(n2003), .IN2(div_exc_out[1]), .IN3(n2041), .IN4(
        \fpu_div_ctl/i_d2stg_zero_in2/N3 ), .Q(n452) );
  NOR2X0 U1311 ( .IN1(n2042), .IN2(n2043), .QN(n2041) );
  AO22X1 U1312 ( .IN1(n1896), .IN2(n1647), .IN3(inq_in2_exp_neq_ffs), .IN4(
        n2040), .Q(n451) );
  MUX21X1 U1313 ( .IN1(div_exc_out[4]), .IN2(n2044), .S(n2001), .Q(n450) );
  OR4X1 U1314 ( .IN1(n2045), .IN2(\fpu_div_ctl/i_d2stg_2inf_in/N3 ), .IN3(
        \fpu_div_ctl/i_d2stg_2zero_in/N3 ), .IN4(
        \fpu_div_ctl/i_d2stg_snan_in1/N3 ), .Q(n2044) );
  AOI21X1 U1315 ( .IN1(n373), .IN2(n370), .IN3(se), .QN(n2045) );
  AO21X1 U1316 ( .IN1(n2003), .IN2(div_sign_out), .IN3(n2046), .Q(n449) );
  NOR4X0 U1317 ( .IN1(n2002), .IN2(\fpu_div_ctl/d2stg_2inf_in ), .IN3(
        \fpu_div_ctl/d2stg_2zero_in ), .IN4(n2047), .QN(n2046) );
  MUX21X1 U1318 ( .IN1(n2048), .IN2(n2049), .S(n2050), .Q(n2047) );
  OA221X1 U1319 ( .IN1(\fpu_div_ctl/d2stg_nan_in2 ), .IN2(n173), .IN3(n629), 
        .IN4(n1877), .IN5(n1539), .Q(n2050) );
  AND3X1 U1320 ( .IN1(n617), .IN2(n1641), .IN3(n1349), .Q(n2049) );
  NAND3X0 U1321 ( .IN1(n2051), .IN2(n1641), .IN3(n1349), .QN(n2048) );
  NAND2X0 U1322 ( .IN1(n629), .IN2(n1878), .QN(n2051) );
  INVX0 U1323 ( .INP(n2004), .ZN(n2002) );
  OAI21X1 U1324 ( .IN1(n28), .IN2(n2001), .IN3(n2052), .QN(n448) );
  NAND4X0 U1325 ( .IN1(n2053), .IN2(n2004), .IN3(n253), .IN4(n979), .QN(n2052)
         );
  INVX0 U1326 ( .INP(n2054), .ZN(n979) );
  NOR2X0 U1327 ( .IN1(n2042), .IN2(se), .QN(n2004) );
  INVX0 U1328 ( .INP(n2043), .ZN(n2053) );
  AO21X1 U1329 ( .IN1(n2007), .IN2(n1873), .IN3(n1355), .Q(n447) );
  AO222X1 U1330 ( .IN1(n2055), .IN2(div_exp_out[0]), .IN3(n2056), .IN4(n2057), 
        .IN5(n1355), .IN6(n2058), .Q(n446) );
  XNOR3X1 U1331 ( .IN1(n2059), .IN2(n2060), .IN3(n2061), .Q(n2057) );
  AO221X1 U1332 ( .IN1(n2056), .IN2(n2062), .IN3(n2055), .IN4(div_exp_out[1]), 
        .IN5(n1355), .Q(n445) );
  XNOR3X1 U1333 ( .IN1(n2063), .IN2(n2064), .IN3(n2065), .Q(n2062) );
  AO221X1 U1334 ( .IN1(n2066), .IN2(n2056), .IN3(n2055), .IN4(div_exp_out[2]), 
        .IN5(n1355), .Q(n444) );
  XNOR3X1 U1335 ( .IN1(n2067), .IN2(n2061), .IN3(n2068), .Q(n2066) );
  AO221X1 U1336 ( .IN1(n2069), .IN2(n2056), .IN3(n2055), .IN4(div_exp_out[3]), 
        .IN5(n1355), .Q(n443) );
  XNOR3X1 U1337 ( .IN1(n2070), .IN2(n2071), .IN3(n2072), .Q(n2069) );
  AO221X1 U1338 ( .IN1(n2073), .IN2(n2056), .IN3(n2055), .IN4(div_exp_out[4]), 
        .IN5(n1355), .Q(n442) );
  XNOR3X1 U1339 ( .IN1(n2074), .IN2(n2075), .IN3(n2076), .Q(n2073) );
  AO221X1 U1340 ( .IN1(n2077), .IN2(n2056), .IN3(n2055), .IN4(div_exp_out[5]), 
        .IN5(n1355), .Q(n441) );
  XNOR3X1 U1341 ( .IN1(n2078), .IN2(n2061), .IN3(n2079), .Q(n2077) );
  AO221X1 U1342 ( .IN1(n2056), .IN2(n2080), .IN3(n2055), .IN4(div_exp_out[6]), 
        .IN5(n1355), .Q(n440) );
  XNOR3X1 U1343 ( .IN1(n2081), .IN2(n2063), .IN3(n2082), .Q(n2080) );
  AO221X1 U1344 ( .IN1(n2056), .IN2(n2083), .IN3(n2055), .IN4(div_exp_out[7]), 
        .IN5(n1355), .Q(n439) );
  XNOR3X1 U1345 ( .IN1(n2063), .IN2(n2084), .IN3(n2085), .Q(n2083) );
  AO22X1 U1346 ( .IN1(n2055), .IN2(n1371), .IN3(n2056), .IN4(n2086), .Q(n438)
         );
  XNOR3X1 U1347 ( .IN1(n2063), .IN2(n2087), .IN3(n2088), .Q(n2086) );
  NOR2X0 U1348 ( .IN1(se), .IN2(n2089), .QN(n437) );
  MUX21X1 U1349 ( .IN1(n2090), .IN2(n18), .S(n2000), .Q(n2089) );
  NAND3X0 U1350 ( .IN1(n1940), .IN2(n2091), .IN3(\fpu_div_frac_dp/n164 ), .QN(
        n2090) );
  NAND4X0 U1351 ( .IN1(n2092), .IN2(n1409), .IN3(n609), .IN4(n2093), .QN(n2091) );
  NOR2X0 U1352 ( .IN1(n2094), .IN2(n2095), .QN(n2093) );
  MUX21X1 U1353 ( .IN1(n2096), .IN2(n2097), .S(n605), .Q(n2095) );
  NAND3X0 U1354 ( .IN1(n590), .IN2(n1396), .IN3(n596), .QN(n2097) );
  NAND3X0 U1355 ( .IN1(n581), .IN2(n1716), .IN3(n610), .QN(n2096) );
  XOR3X1 U1356 ( .IN1(n2098), .IN2(n2099), .IN3(n2063), .Q(n1940) );
  OA22X1 U1357 ( .IN1(n576), .IN2(n607), .IN3(n578), .IN4(n613), .Q(n2099) );
  OA22X1 U1358 ( .IN1(n2063), .IN2(n2100), .IN3(n2087), .IN4(n2088), .Q(n2098)
         );
  AND2X1 U1359 ( .IN1(n2088), .IN2(n2087), .Q(n2100) );
  OA22X1 U1360 ( .IN1(n618), .IN2(n578), .IN3(n576), .IN4(n29), .Q(n2087) );
  AO22X1 U1361 ( .IN1(n2101), .IN2(n2102), .IN3(n2063), .IN4(n2103), .Q(n2088)
         );
  OR2X1 U1362 ( .IN1(n2102), .IN2(n2101), .Q(n2103) );
  AO21X1 U1363 ( .IN1(n1867), .IN2(n2007), .IN3(n2104), .Q(n436) );
  AND4X1 U1364 ( .IN1(n2105), .IN2(n2106), .IN3(n613), .IN4(n2107), .Q(n2104)
         );
  AO22X1 U1365 ( .IN1(n2007), .IN2(div_exc_out[2]), .IN3(n2105), .IN4(n2108), 
        .Q(n435) );
  NAND2X0 U1366 ( .IN1(n613), .IN2(n2109), .QN(n2108) );
  NAND3X0 U1367 ( .IN1(n2110), .IN2(n2111), .IN3(n218), .QN(n2109) );
  NAND2X0 U1368 ( .IN1(n2022), .IN2(n2014), .QN(n2111) );
  AND4X1 U1369 ( .IN1(n2112), .IN2(n2113), .IN3(n2114), .IN4(n2115), .Q(n2014)
         );
  NOR4X0 U1370 ( .IN1(n2116), .IN2(n2117), .IN3(n2118), .IN4(n2119), .QN(n2115) );
  NAND4X0 U1371 ( .IN1(\fpu_div_frac_dp/n96 ), .IN2(\fpu_div_frac_dp/n93 ), 
        .IN3(\fpu_div_frac_dp/n99 ), .IN4(n2120), .QN(n2119) );
  NOR3X0 U1372 ( .IN1(n1377), .IN2(n1402), .IN3(n1361), .QN(n2120) );
  NAND4X0 U1373 ( .IN1(\fpu_div_frac_dp/n79 ), .IN2(\fpu_div_frac_dp/n76 ), 
        .IN3(\fpu_div_frac_dp/n83 ), .IN4(n2121), .QN(n2118) );
  NOR4X0 U1374 ( .IN1(n1357), .IN2(n1362), .IN3(n1406), .IN4(n1382), .QN(n2121) );
  NAND4X0 U1375 ( .IN1(\fpu_div_frac_dp/n61 ), .IN2(\fpu_div_frac_dp/n58 ), 
        .IN3(\fpu_div_frac_dp/n64 ), .IN4(n2122), .QN(n2117) );
  NOR4X0 U1376 ( .IN1(n1358), .IN2(n1363), .IN3(n1405), .IN4(n1381), .QN(n2122) );
  NAND4X0 U1377 ( .IN1(\fpu_div_frac_dp/n40 ), .IN2(\fpu_div_frac_dp/n4 ), 
        .IN3(\fpu_div_frac_dp/n43 ), .IN4(n2123), .QN(n2116) );
  NOR4X0 U1378 ( .IN1(n1460), .IN2(n1359), .IN3(n1366), .IN4(n1380), .QN(n2123) );
  NOR4X0 U1379 ( .IN1(n2124), .IN2(n2125), .IN3(n2126), .IN4(n2127), .QN(n2114) );
  NAND3X0 U1380 ( .IN1(\fpu_div_frac_dp/n132 ), .IN2(\fpu_div_frac_dp/n13 ), 
        .IN3(\fpu_div_frac_dp/n135 ), .QN(n2127) );
  NAND4X0 U1381 ( .IN1(\fpu_div_frac_dp/n129 ), .IN2(\fpu_div_frac_dp/n126 ), 
        .IN3(\fpu_div_frac_dp/n123 ), .IN4(\fpu_div_frac_dp/n120 ), .QN(n2126)
         );
  NAND3X0 U1382 ( .IN1(\fpu_div_frac_dp/n114 ), .IN2(\fpu_div_frac_dp/n111 ), 
        .IN3(\fpu_div_frac_dp/n117 ), .QN(n2125) );
  NAND4X0 U1383 ( .IN1(\fpu_div_frac_dp/n108 ), .IN2(\fpu_div_frac_dp/n105 ), 
        .IN3(\fpu_div_frac_dp/n102 ), .IN4(\fpu_div_frac_dp/n10 ), .QN(n2124)
         );
  NOR4X0 U1384 ( .IN1(n2128), .IN2(n1364), .IN3(n1378), .IN4(n1407), .QN(n2113) );
  NAND4X0 U1385 ( .IN1(\fpu_div_frac_dp/n147 ), .IN2(\fpu_div_frac_dp/n144 ), 
        .IN3(\fpu_div_frac_dp/n141 ), .IN4(\fpu_div_frac_dp/n138 ), .QN(n2128)
         );
  NOR4X0 U1386 ( .IN1(n2129), .IN2(n1365), .IN3(n1404), .IN4(n1379), .QN(n2112) );
  NAND4X0 U1387 ( .IN1(\fpu_div_frac_dp/n19 ), .IN2(\fpu_div_frac_dp/n162 ), 
        .IN3(\fpu_div_frac_dp/n160 ), .IN4(\fpu_div_frac_dp/n16 ), .QN(n2129)
         );
  INVX0 U1388 ( .INP(n2130), .ZN(n2110) );
  NOR2X0 U1389 ( .IN1(n1393), .IN2(se), .QN(n2007) );
  AO22X1 U1390 ( .IN1(n1896), .IN2(n1859), .IN3(inq_in1[62]), .IN4(n2040), .Q(
        n434) );
  AO22X1 U1391 ( .IN1(n1896), .IN2(n1865), .IN3(inq_in1[61]), .IN4(n2040), .Q(
        n433) );
  AO22X1 U1392 ( .IN1(n1896), .IN2(n1858), .IN3(inq_in1[60]), .IN4(n2040), .Q(
        n432) );
  AO22X1 U1393 ( .IN1(n1896), .IN2(n1861), .IN3(inq_in1[59]), .IN4(n2040), .Q(
        n431) );
  AO22X1 U1394 ( .IN1(n1897), .IN2(n1862), .IN3(inq_in1[58]), .IN4(n2040), .Q(
        n430) );
  AO22X1 U1395 ( .IN1(n1896), .IN2(n1863), .IN3(inq_in1[57]), .IN4(n2040), .Q(
        n429) );
  AO22X1 U1396 ( .IN1(n1896), .IN2(n1860), .IN3(inq_in1[56]), .IN4(n2040), .Q(
        n428) );
  AO22X1 U1397 ( .IN1(n1896), .IN2(n1855), .IN3(inq_in1[55]), .IN4(n2040), .Q(
        n427) );
  AO22X1 U1398 ( .IN1(n1896), .IN2(n1871), .IN3(inq_in1[54]), .IN4(n2040), .Q(
        n426) );
  AO22X1 U1399 ( .IN1(n1896), .IN2(n1876), .IN3(inq_in1[53]), .IN4(n2040), .Q(
        n425) );
  AO22X1 U1400 ( .IN1(n1895), .IN2(n1872), .IN3(inq_in1[52]), .IN4(n2040), .Q(
        n424) );
  AO22X1 U1401 ( .IN1(n1896), .IN2(n1491), .IN3(inq_in2[62]), .IN4(n2040), .Q(
        n423) );
  AO22X1 U1402 ( .IN1(n1895), .IN2(n1676), .IN3(inq_in2[61]), .IN4(n2040), .Q(
        n422) );
  AO22X1 U1403 ( .IN1(n1895), .IN2(n1642), .IN3(inq_in2[60]), .IN4(n2040), .Q(
        n421) );
  AO22X1 U1404 ( .IN1(n1895), .IN2(n1640), .IN3(inq_in2[59]), .IN4(n2040), .Q(
        n420) );
  AO22X1 U1405 ( .IN1(n1895), .IN2(n1534), .IN3(inq_in2[58]), .IN4(n2040), .Q(
        n419) );
  AO22X1 U1406 ( .IN1(n622), .IN2(n1897), .IN3(inq_in2[57]), .IN4(n2040), .Q(
        n418) );
  AO22X1 U1407 ( .IN1(n1895), .IN2(n1532), .IN3(inq_in2[56]), .IN4(n2040), .Q(
        n417) );
  AO22X1 U1408 ( .IN1(n623), .IN2(n1897), .IN3(inq_in2[55]), .IN4(n2040), .Q(
        n416) );
  AO22X1 U1409 ( .IN1(n1895), .IN2(n1724), .IN3(inq_in2[54]), .IN4(n2040), .Q(
        n415) );
  AO22X1 U1410 ( .IN1(n1895), .IN2(n1730), .IN3(inq_in2[53]), .IN4(n2040), .Q(
        n414) );
  AO22X1 U1411 ( .IN1(n1895), .IN2(n1725), .IN3(inq_in2[52]), .IN4(n2040), .Q(
        n413) );
  NOR2X0 U1412 ( .IN1(n2131), .IN2(se), .QN(n2040) );
  OA22X1 U1413 ( .IN1(n1985), .IN2(n2132), .IN3(n29), .IN4(n2133), .Q(n292) );
  XNOR3X1 U1414 ( .IN1(n1946), .IN2(n1948), .IN3(n1950), .Q(n2132) );
  INVX0 U1415 ( .INP(n1952), .ZN(n1950) );
  AO22X1 U1416 ( .IN1(n1962), .IN2(n1963), .IN3(n1961), .IN4(n2134), .Q(n1952)
         );
  OR2X1 U1417 ( .IN1(n1962), .IN2(n1963), .Q(n2134) );
  AND3X1 U1418 ( .IN1(n2135), .IN2(n2136), .IN3(n587), .Q(n1961) );
  OR2X1 U1419 ( .IN1(n1491), .IN2(n181), .Q(n2136) );
  AOI22X1 U1420 ( .IN1(n1967), .IN2(n1966), .IN3(n1965), .IN4(n2137), .QN(
        n1963) );
  OR2X1 U1421 ( .IN1(n1966), .IN2(n1967), .Q(n2137) );
  AOI21X1 U1422 ( .IN1(n2135), .IN2(n1676), .IN3(n1951), .QN(n1965) );
  OAI22X1 U1423 ( .IN1(n98), .IN2(n587), .IN3(n31), .IN4(n117), .QN(n1966) );
  AO22X1 U1424 ( .IN1(n2138), .IN2(n2139), .IN3(n2140), .IN4(n2141), .Q(n1967)
         );
  NAND2X0 U1425 ( .IN1(n2142), .IN2(n2143), .QN(n2140) );
  INVX0 U1426 ( .INP(n2142), .ZN(n2139) );
  INVX0 U1427 ( .INP(n2143), .ZN(n2138) );
  OA22X1 U1428 ( .IN1(n587), .IN2(n97), .IN3(n117), .IN4(n30), .Q(n1962) );
  NOR2X0 U1429 ( .IN1(n29), .IN2(n117), .QN(n1948) );
  AND2X1 U1430 ( .IN1(n2144), .IN2(n2145), .Q(n291) );
  NAND3X0 U1431 ( .IN1(n41), .IN2(n40), .IN3(n93), .QN(n2145) );
  OA22X1 U1432 ( .IN1(n2146), .IN2(n1985), .IN3(n32), .IN4(n2133), .Q(n290) );
  XNOR3X1 U1433 ( .IN1(n2143), .IN2(n2142), .IN3(n2141), .Q(n2146) );
  AO22X1 U1434 ( .IN1(n1971), .IN2(n1970), .IN3(n2147), .IN4(n1969), .Q(n2141)
         );
  NAND3X0 U1435 ( .IN1(n601), .IN2(n184), .IN3(n2148), .QN(n1969) );
  OA22X1 U1436 ( .IN1(n182), .IN2(n1491), .IN3(n181), .IN4(n1640), .Q(n2148)
         );
  OR2X1 U1437 ( .IN1(n1970), .IN2(n1971), .Q(n2147) );
  OAI222X1 U1438 ( .IN1(n117), .IN2(n33), .IN3(n100), .IN4(n587), .IN5(n601), 
        .IN6(n97), .QN(n1970) );
  AO22X1 U1439 ( .IN1(n1975), .IN2(n1974), .IN3(n2149), .IN4(n1973), .Q(n1971)
         );
  OAI221X1 U1440 ( .IN1(n1676), .IN2(n182), .IN3(n1534), .IN4(n181), .IN5(n184), .QN(n1973) );
  OR2X1 U1441 ( .IN1(n1974), .IN2(n1975), .Q(n2149) );
  OAI222X1 U1442 ( .IN1(n117), .IN2(n34), .IN3(n101), .IN4(n587), .IN5(n601), 
        .IN6(n98), .QN(n1974) );
  AO22X1 U1443 ( .IN1(n2150), .IN2(n2151), .IN3(n2152), .IN4(n2153), .Q(n1975)
         );
  OR2X1 U1444 ( .IN1(n2151), .IN2(n2150), .Q(n2152) );
  OA22X1 U1445 ( .IN1(n99), .IN2(n587), .IN3(n32), .IN4(n117), .Q(n2142) );
  AO21X1 U1446 ( .IN1(n2135), .IN2(n1642), .IN3(n1951), .Q(n2143) );
  INVX0 U1447 ( .INP(n1946), .ZN(n1951) );
  NAND2X0 U1448 ( .IN1(n181), .IN2(n2135), .QN(n1946) );
  AND2X1 U1449 ( .IN1(n182), .IN2(n184), .Q(n2135) );
  OA22X1 U1450 ( .IN1(n1985), .IN2(n2154), .IN3(n590), .IN4(n2133), .Q(n289)
         );
  XNOR3X1 U1451 ( .IN1(n2153), .IN2(n2151), .IN3(n2150), .Q(n2154) );
  NAND3X0 U1452 ( .IN1(n2155), .IN2(n587), .IN3(n2156), .QN(n2150) );
  OA22X1 U1453 ( .IN1(n182), .IN2(n1642), .IN3(n622), .IN4(n181), .Q(n2156) );
  MUX21X1 U1454 ( .IN1(n184), .IN2(n185), .S(n1540), .Q(n2155) );
  OAI222X1 U1455 ( .IN1(n117), .IN2(n590), .IN3(n102), .IN4(n587), .IN5(n601), 
        .IN6(n99), .QN(n2151) );
  AO22X1 U1456 ( .IN1(n1980), .IN2(n2157), .IN3(n2158), .IN4(n1978), .Q(n2153)
         );
  NAND4X0 U1457 ( .IN1(n2159), .IN2(n601), .IN3(n2160), .IN4(n587), .QN(n1978)
         );
  OA22X1 U1458 ( .IN1(n182), .IN2(n1640), .IN3(n181), .IN4(n1532), .Q(n2160)
         );
  MUX21X1 U1459 ( .IN1(n184), .IN2(n185), .S(n1392), .Q(n2159) );
  NAND2X0 U1460 ( .IN1(n1979), .IN2(n2161), .QN(n2158) );
  INVX0 U1461 ( .INP(n1979), .ZN(n2157) );
  OA222X1 U1462 ( .IN1(n103), .IN2(n587), .IN3(n100), .IN4(n601), .IN5(n117), 
        .IN6(n592), .Q(n1979) );
  INVX0 U1463 ( .INP(n2161), .ZN(n1980) );
  OA22X1 U1464 ( .IN1(n2162), .IN2(n2163), .IN3(n2164), .IN4(n2165), .Q(n2161)
         );
  AND2X1 U1465 ( .IN1(n2163), .IN2(n2162), .Q(n2164) );
  OA22X1 U1466 ( .IN1(n1985), .IN2(n2166), .IN3(n610), .IN4(n2133), .Q(n286)
         );
  XOR3X1 U1467 ( .IN1(n2165), .IN2(n2163), .IN3(n2162), .Q(n2166) );
  AND3X1 U1468 ( .IN1(n2167), .IN2(n601), .IN3(n2168), .Q(n2162) );
  OA22X1 U1469 ( .IN1(n182), .IN2(n1534), .IN3(n623), .IN4(n181), .Q(n2168) );
  MUX21X1 U1470 ( .IN1(n184), .IN2(n185), .S(n1546), .Q(n2167) );
  OA222X1 U1471 ( .IN1(n104), .IN2(n587), .IN3(n101), .IN4(n601), .IN5(n117), 
        .IN6(n610), .Q(n2163) );
  AOI22X1 U1472 ( .IN1(n2169), .IN2(n2170), .IN3(n2171), .IN4(n2172), .QN(
        n2165) );
  NAND2X0 U1473 ( .IN1(n2173), .IN2(n2174), .QN(n2171) );
  INVX0 U1474 ( .INP(n2173), .ZN(n2170) );
  OA22X1 U1475 ( .IN1(n1985), .IN2(n2175), .IN3(n596), .IN4(n2133), .Q(n285)
         );
  XNOR3X1 U1476 ( .IN1(n2173), .IN2(n2174), .IN3(n2172), .Q(n2175) );
  AO22X1 U1477 ( .IN1(n1984), .IN2(n1983), .IN3(n1982), .IN4(n2176), .Q(n2172)
         );
  OR2X1 U1478 ( .IN1(n1983), .IN2(n1984), .Q(n2176) );
  OAI222X1 U1479 ( .IN1(n106), .IN2(n587), .IN3(n103), .IN4(n601), .IN5(n117), 
        .IN6(n609), .QN(n1983) );
  NAND3X0 U1480 ( .IN1(n2177), .IN2(n587), .IN3(n2178), .QN(n1984) );
  OA22X1 U1481 ( .IN1(n182), .IN2(n1532), .IN3(n181), .IN4(n1730), .Q(n2178)
         );
  MUX21X1 U1482 ( .IN1(n184), .IN2(n185), .S(n1544), .Q(n2177) );
  INVX0 U1483 ( .INP(n2169), .ZN(n2174) );
  NAND3X0 U1484 ( .IN1(n2179), .IN2(n587), .IN3(n2180), .QN(n2169) );
  OA22X1 U1485 ( .IN1(n181), .IN2(n1724), .IN3(n622), .IN4(n182), .Q(n2180) );
  MUX21X1 U1486 ( .IN1(n184), .IN2(n185), .S(n1394), .Q(n2179) );
  OA222X1 U1487 ( .IN1(n596), .IN2(n117), .IN3(n601), .IN4(n102), .IN5(n587), 
        .IN6(n105), .Q(n2173) );
  OA22X1 U1488 ( .IN1(n1985), .IN2(n2181), .IN3(n605), .IN4(n2133), .Q(n282)
         );
  AO21X1 U1489 ( .IN1(n2182), .IN2(n2183), .IN3(n1982), .Q(n2181) );
  NOR2X0 U1490 ( .IN1(n2183), .IN2(n2182), .QN(n1982) );
  AND3X1 U1491 ( .IN1(n2184), .IN2(n601), .IN3(n2185), .Q(n2183) );
  OA22X1 U1492 ( .IN1(n181), .IN2(n1725), .IN3(n623), .IN4(n182), .Q(n2185) );
  MUX21X1 U1493 ( .IN1(n184), .IN2(n185), .S(n1398), .Q(n2184) );
  OA222X1 U1494 ( .IN1(n601), .IN2(n104), .IN3(n605), .IN4(n117), .IN5(n587), 
        .IN6(n107), .Q(n2182) );
  NAND2X0 U1495 ( .IN1(n2144), .IN2(n2186), .QN(n1985) );
  NAND4X0 U1496 ( .IN1(n185), .IN2(n2187), .IN3(n184), .IN4(n2188), .QN(n2186)
         );
  NOR2X0 U1497 ( .IN1(n1942), .IN2(se), .QN(n2144) );
  INVX0 U1498 ( .INP(n2133), .ZN(n1942) );
  NAND4X0 U1499 ( .IN1(n185), .IN2(n2187), .IN3(n2189), .IN4(n1549), .QN(n2133) );
  NAND2X0 U1500 ( .IN1(n2027), .IN2(n1373), .QN(n272) );
  INVX0 U1501 ( .INP(n2190), .ZN(n2027) );
  OA22X1 U1502 ( .IN1(n2191), .IN2(n1939), .IN3(n2192), .IN4(n584), .Q(n248)
         );
  XOR3X1 U1503 ( .IN1(n2063), .IN2(n2193), .IN3(n2194), .Q(n2191) );
  OA22X1 U1504 ( .IN1(n2195), .IN2(n1939), .IN3(n2192), .IN4(n580), .Q(n247)
         );
  XOR3X1 U1505 ( .IN1(n2063), .IN2(n2196), .IN3(n2197), .Q(n2195) );
  OA22X1 U1506 ( .IN1(n2198), .IN2(n1939), .IN3(n2192), .IN4(n599), .Q(n246)
         );
  INVX0 U1507 ( .INP(n2055), .ZN(n2192) );
  NAND2X0 U1508 ( .IN1(n1941), .IN2(n2199), .QN(n2055) );
  NAND4X0 U1509 ( .IN1(n2200), .IN2(n613), .IN3(n2201), .IN4(n1047), .QN(n2199) );
  NAND3X0 U1510 ( .IN1(n193), .IN2(n2003), .IN3(n194), .QN(n1941) );
  INVX0 U1511 ( .INP(n2001), .ZN(n2003) );
  NAND2X0 U1512 ( .IN1(n2042), .IN2(n1047), .QN(n2001) );
  INVX0 U1513 ( .INP(n2056), .ZN(n1939) );
  OA221X1 U1514 ( .IN1(n2202), .IN2(n1552), .IN3(n194), .IN4(n613), .IN5(n1047), .Q(n2056) );
  OAI21X1 U1515 ( .IN1(n2201), .IN2(n2203), .IN3(n2042), .QN(n2202) );
  NAND2X0 U1516 ( .IN1(n2106), .IN2(n2204), .QN(n2201) );
  XOR3X1 U1517 ( .IN1(n2063), .IN2(n2101), .IN3(n2102), .Q(n2198) );
  AO22X1 U1518 ( .IN1(n2196), .IN2(n2197), .IN3(n2063), .IN4(n2205), .Q(n2102)
         );
  OR2X1 U1519 ( .IN1(n2197), .IN2(n2196), .Q(n2205) );
  AO22X1 U1520 ( .IN1(n2193), .IN2(n2194), .IN3(n2063), .IN4(n2206), .Q(n2197)
         );
  OR2X1 U1521 ( .IN1(n2194), .IN2(n2193), .Q(n2206) );
  AO22X1 U1522 ( .IN1(n2084), .IN2(n2085), .IN3(n2063), .IN4(n2207), .Q(n2194)
         );
  OR2X1 U1523 ( .IN1(n2085), .IN2(n2084), .Q(n2207) );
  AO22X1 U1524 ( .IN1(n2081), .IN2(n2082), .IN3(n2063), .IN4(n2208), .Q(n2085)
         );
  OR2X1 U1525 ( .IN1(n2082), .IN2(n2081), .Q(n2208) );
  AO22X1 U1526 ( .IN1(n2079), .IN2(n2061), .IN3(n2078), .IN4(n2209), .Q(n2082)
         );
  OR2X1 U1527 ( .IN1(n2079), .IN2(n2061), .Q(n2209) );
  OA22X1 U1528 ( .IN1(n603), .IN2(n578), .IN3(n590), .IN4(n576), .Q(n2078) );
  AO22X1 U1529 ( .IN1(n2075), .IN2(n2076), .IN3(n2210), .IN4(n2074), .Q(n2079)
         );
  OR2X1 U1530 ( .IN1(n2076), .IN2(n2075), .Q(n2210) );
  AO22X1 U1531 ( .IN1(n2070), .IN2(n2072), .IN3(n2071), .IN4(n2211), .Q(n2076)
         );
  OR2X1 U1532 ( .IN1(n2072), .IN2(n2070), .Q(n2211) );
  OA22X1 U1533 ( .IN1(n610), .IN2(n576), .IN3(n582), .IN4(n578), .Q(n2071) );
  AO22X1 U1534 ( .IN1(n2068), .IN2(n2061), .IN3(n2067), .IN4(n2212), .Q(n2072)
         );
  OR2X1 U1535 ( .IN1(n2068), .IN2(n2061), .Q(n2212) );
  OA22X1 U1536 ( .IN1(n596), .IN2(n576), .IN3(n579), .IN4(n578), .Q(n2067) );
  AO22X1 U1537 ( .IN1(n2064), .IN2(n2065), .IN3(n2063), .IN4(n2213), .Q(n2068)
         );
  OR2X1 U1538 ( .IN1(n2065), .IN2(n2064), .Q(n2213) );
  AO22X1 U1539 ( .IN1(n2059), .IN2(n2061), .IN3(n2060), .IN4(n2214), .Q(n2065)
         );
  OR2X1 U1540 ( .IN1(n2061), .IN2(n2059), .Q(n2214) );
  AO21X1 U1541 ( .IN1(n581), .IN2(n2074), .IN3(n2063), .Q(n2061) );
  OA22X1 U1542 ( .IN1(n605), .IN2(n576), .IN3(n578), .IN4(n218), .Q(n2059) );
  OA22X1 U1543 ( .IN1(n609), .IN2(n576), .IN3(n595), .IN4(n578), .Q(n2064) );
  AO21X1 U1544 ( .IN1(n611), .IN2(n2074), .IN3(n2063), .Q(n2070) );
  INVX0 U1545 ( .INP(n2215), .ZN(n2074) );
  OA22X1 U1546 ( .IN1(n592), .IN2(n576), .IN3(n583), .IN4(n578), .Q(n2075) );
  OA22X1 U1547 ( .IN1(n614), .IN2(n578), .IN3(n576), .IN4(n34), .Q(n2081) );
  OA22X1 U1548 ( .IN1(n598), .IN2(n578), .IN3(n576), .IN4(n33), .Q(n2084) );
  OA22X1 U1549 ( .IN1(n584), .IN2(n578), .IN3(n576), .IN4(n32), .Q(n2193) );
  OA22X1 U1550 ( .IN1(n580), .IN2(n578), .IN3(n576), .IN4(n31), .Q(n2196) );
  OA22X1 U1551 ( .IN1(n599), .IN2(n578), .IN3(n576), .IN4(n30), .Q(n2101) );
  NOR2X0 U1552 ( .IN1(n1579), .IN2(n2215), .QN(n2063) );
  NOR2X0 U1553 ( .IN1(n18), .IN2(n193), .QN(n2215) );
  AND3X1 U1554 ( .IN1(n613), .IN2(n2216), .IN3(n2105), .Q(n1355) );
  NOR2X0 U1555 ( .IN1(\fpu_div_frac_dp/rclk ), .IN2(\fpu_div_frac_dp/n168 ), 
        .QN(\fpu_div_frac_dp/n985 ) );
  INVX0 U1556 ( .INP(rclk), .ZN(\fpu_div_frac_dp/rclk ) );
  NOR2X0 U1557 ( .IN1(se), .IN2(n1597), .QN(\fpu_div_frac_dp/n609 ) );
  AO22X1 U1558 ( .IN1(inq_in1[0]), .IN2(n1881), .IN3(n1888), .IN4(n1819), .Q(
        \fpu_div_frac_dp/n1439 ) );
  AO22X1 U1559 ( .IN1(inq_in1[1]), .IN2(n1880), .IN3(n1888), .IN4(n1820), .Q(
        \fpu_div_frac_dp/n1438 ) );
  AO22X1 U1560 ( .IN1(inq_in1[2]), .IN2(n1879), .IN3(n1888), .IN4(n1821), .Q(
        \fpu_div_frac_dp/n1437 ) );
  AO22X1 U1561 ( .IN1(inq_in1[3]), .IN2(n1882), .IN3(n1888), .IN4(n1822), .Q(
        \fpu_div_frac_dp/n1436 ) );
  AO22X1 U1562 ( .IN1(inq_in1[4]), .IN2(n1881), .IN3(n1888), .IN4(n1823), .Q(
        \fpu_div_frac_dp/n1435 ) );
  AO22X1 U1563 ( .IN1(inq_in1[5]), .IN2(n1880), .IN3(n1888), .IN4(n1824), .Q(
        \fpu_div_frac_dp/n1434 ) );
  AO22X1 U1564 ( .IN1(inq_in1[6]), .IN2(n1879), .IN3(n1888), .IN4(n1825), .Q(
        \fpu_div_frac_dp/n1433 ) );
  AO22X1 U1565 ( .IN1(inq_in1[7]), .IN2(n1882), .IN3(n1888), .IN4(n1826), .Q(
        \fpu_div_frac_dp/n1432 ) );
  AO22X1 U1566 ( .IN1(inq_in1[8]), .IN2(n1881), .IN3(n1888), .IN4(n1827), .Q(
        \fpu_div_frac_dp/n1431 ) );
  AO22X1 U1567 ( .IN1(inq_in1[9]), .IN2(n1880), .IN3(n1888), .IN4(n1848), .Q(
        \fpu_div_frac_dp/n1430 ) );
  AO22X1 U1568 ( .IN1(inq_in1[10]), .IN2(n1879), .IN3(n1888), .IN4(n1846), .Q(
        \fpu_div_frac_dp/n1429 ) );
  AO22X1 U1569 ( .IN1(inq_in1[11]), .IN2(n1882), .IN3(n1888), .IN4(n1828), .Q(
        \fpu_div_frac_dp/n1428 ) );
  AO22X1 U1570 ( .IN1(inq_in1[12]), .IN2(n1881), .IN3(n1888), .IN4(n1829), .Q(
        \fpu_div_frac_dp/n1427 ) );
  AO22X1 U1571 ( .IN1(inq_in1[13]), .IN2(n1880), .IN3(n1889), .IN4(n1830), .Q(
        \fpu_div_frac_dp/n1426 ) );
  AO22X1 U1572 ( .IN1(inq_in1[14]), .IN2(n1879), .IN3(n1889), .IN4(n1831), .Q(
        \fpu_div_frac_dp/n1425 ) );
  AO22X1 U1573 ( .IN1(inq_in1[15]), .IN2(n1882), .IN3(n1889), .IN4(n1832), .Q(
        \fpu_div_frac_dp/n1424 ) );
  AO22X1 U1574 ( .IN1(inq_in1[16]), .IN2(n1881), .IN3(n1889), .IN4(n1833), .Q(
        \fpu_div_frac_dp/n1423 ) );
  AO22X1 U1575 ( .IN1(inq_in1[17]), .IN2(n1880), .IN3(n1889), .IN4(n1834), .Q(
        \fpu_div_frac_dp/n1422 ) );
  AO22X1 U1576 ( .IN1(inq_in1[18]), .IN2(n1879), .IN3(n1889), .IN4(n1835), .Q(
        \fpu_div_frac_dp/n1421 ) );
  AO22X1 U1577 ( .IN1(inq_in1[19]), .IN2(n1882), .IN3(n1889), .IN4(n1836), .Q(
        \fpu_div_frac_dp/n1420 ) );
  AO22X1 U1578 ( .IN1(inq_in1[20]), .IN2(n1881), .IN3(n1889), .IN4(n1837), .Q(
        \fpu_div_frac_dp/n1419 ) );
  AO22X1 U1579 ( .IN1(inq_in1[21]), .IN2(n1880), .IN3(n1889), .IN4(n1838), .Q(
        \fpu_div_frac_dp/n1418 ) );
  AO22X1 U1580 ( .IN1(inq_in1[22]), .IN2(n1879), .IN3(n1889), .IN4(n1839), .Q(
        \fpu_div_frac_dp/n1417 ) );
  AO22X1 U1581 ( .IN1(inq_in1[23]), .IN2(n1882), .IN3(n1889), .IN4(n1840), .Q(
        \fpu_div_frac_dp/n1416 ) );
  AO22X1 U1582 ( .IN1(inq_in1[24]), .IN2(n1881), .IN3(n1889), .IN4(n1841), .Q(
        \fpu_div_frac_dp/n1415 ) );
  AO22X1 U1583 ( .IN1(inq_in1[25]), .IN2(n1880), .IN3(n1889), .IN4(n1842), .Q(
        \fpu_div_frac_dp/n1414 ) );
  AO22X1 U1584 ( .IN1(inq_in1[26]), .IN2(n1879), .IN3(n1889), .IN4(n1843), .Q(
        \fpu_div_frac_dp/n1413 ) );
  AO22X1 U1585 ( .IN1(inq_in1[27]), .IN2(n1882), .IN3(n1889), .IN4(n1844), .Q(
        \fpu_div_frac_dp/n1412 ) );
  AO22X1 U1586 ( .IN1(inq_in1[28]), .IN2(n1881), .IN3(n1890), .IN4(n1814), .Q(
        \fpu_div_frac_dp/n1411 ) );
  AO22X1 U1587 ( .IN1(inq_in1[29]), .IN2(n1880), .IN3(n1890), .IN4(n1810), .Q(
        \fpu_div_frac_dp/n1410 ) );
  AO22X1 U1588 ( .IN1(inq_in1[30]), .IN2(n1879), .IN3(n1890), .IN4(n1812), .Q(
        \fpu_div_frac_dp/n1409 ) );
  AO22X1 U1589 ( .IN1(inq_in1[31]), .IN2(n1882), .IN3(n1890), .IN4(n1813), .Q(
        \fpu_div_frac_dp/n1408 ) );
  AO22X1 U1590 ( .IN1(inq_in1[32]), .IN2(n1881), .IN3(n1890), .IN4(n1804), .Q(
        \fpu_div_frac_dp/n1407 ) );
  AO22X1 U1591 ( .IN1(inq_in1[33]), .IN2(n1880), .IN3(n1890), .IN4(n1787), .Q(
        \fpu_div_frac_dp/n1406 ) );
  AO22X1 U1592 ( .IN1(inq_in1[34]), .IN2(n1879), .IN3(n1890), .IN4(n1788), .Q(
        \fpu_div_frac_dp/n1405 ) );
  AO22X1 U1593 ( .IN1(inq_in1[35]), .IN2(n1882), .IN3(n1890), .IN4(n1789), .Q(
        \fpu_div_frac_dp/n1404 ) );
  AO22X1 U1594 ( .IN1(inq_in1[36]), .IN2(n1881), .IN3(n1890), .IN4(n1790), .Q(
        \fpu_div_frac_dp/n1403 ) );
  AO22X1 U1595 ( .IN1(inq_in1[37]), .IN2(n1880), .IN3(n1890), .IN4(n1791), .Q(
        \fpu_div_frac_dp/n1402 ) );
  AO22X1 U1596 ( .IN1(inq_in1[38]), .IN2(n1879), .IN3(n1890), .IN4(n1792), .Q(
        \fpu_div_frac_dp/n1401 ) );
  AO22X1 U1597 ( .IN1(inq_in1[39]), .IN2(n1882), .IN3(n1890), .IN4(n1793), .Q(
        \fpu_div_frac_dp/n1400 ) );
  AO22X1 U1598 ( .IN1(inq_in1[40]), .IN2(n1881), .IN3(n1890), .IN4(n1794), .Q(
        \fpu_div_frac_dp/n1399 ) );
  AO22X1 U1599 ( .IN1(inq_in1[41]), .IN2(n1880), .IN3(n1890), .IN4(n1795), .Q(
        \fpu_div_frac_dp/n1398 ) );
  AO22X1 U1600 ( .IN1(inq_in1[42]), .IN2(n1879), .IN3(n1890), .IN4(n1796), .Q(
        \fpu_div_frac_dp/n1397 ) );
  AO22X1 U1601 ( .IN1(inq_in1[43]), .IN2(n1882), .IN3(n1891), .IN4(n1797), .Q(
        \fpu_div_frac_dp/n1396 ) );
  AO22X1 U1602 ( .IN1(inq_in1[44]), .IN2(n1881), .IN3(n1891), .IN4(n1798), .Q(
        \fpu_div_frac_dp/n1395 ) );
  AO22X1 U1603 ( .IN1(inq_in1[45]), .IN2(n1880), .IN3(n1891), .IN4(n1799), .Q(
        \fpu_div_frac_dp/n1394 ) );
  AO22X1 U1604 ( .IN1(inq_in1[46]), .IN2(n1879), .IN3(n1891), .IN4(n1800), .Q(
        \fpu_div_frac_dp/n1393 ) );
  AO22X1 U1605 ( .IN1(inq_in1[47]), .IN2(n1882), .IN3(n1891), .IN4(n1801), .Q(
        \fpu_div_frac_dp/n1392 ) );
  AO22X1 U1606 ( .IN1(inq_in1[48]), .IN2(n1881), .IN3(n1891), .IN4(n1802), .Q(
        \fpu_div_frac_dp/n1391 ) );
  AO22X1 U1607 ( .IN1(inq_in1[49]), .IN2(n1880), .IN3(n1891), .IN4(n1803), .Q(
        \fpu_div_frac_dp/n1390 ) );
  AO22X1 U1608 ( .IN1(inq_in1[50]), .IN2(n1879), .IN3(n1891), .IN4(n1805), .Q(
        \fpu_div_frac_dp/n1389 ) );
  AO22X1 U1609 ( .IN1(n1879), .IN2(inq_in1[51]), .IN3(n1891), .IN4(n1670), .Q(
        \fpu_div_frac_dp/n1388 ) );
  AO22X1 U1610 ( .IN1(n1882), .IN2(inq_in1[52]), .IN3(n1891), .IN4(n1811), .Q(
        \fpu_div_frac_dp/n1387 ) );
  AO22X1 U1611 ( .IN1(n1881), .IN2(inq_in1[53]), .IN3(n1891), .IN4(n1847), .Q(
        \fpu_div_frac_dp/n1386 ) );
  AO22X1 U1612 ( .IN1(n1880), .IN2(inq_in1[54]), .IN3(n1891), .IN4(n1850), .Q(
        \fpu_div_frac_dp/n1385 ) );
  AO22X1 U1613 ( .IN1(inq_in2[0]), .IN2(n1882), .IN3(n1891), .IN4(n1816), .Q(
        \fpu_div_frac_dp/n1384 ) );
  AO22X1 U1614 ( .IN1(inq_in2[1]), .IN2(n1881), .IN3(n1891), .IN4(n1691), .Q(
        \fpu_div_frac_dp/n1383 ) );
  AO22X1 U1615 ( .IN1(inq_in2[2]), .IN2(n1880), .IN3(n1892), .IN4(n1690), .Q(
        \fpu_div_frac_dp/n1382 ) );
  AO22X1 U1616 ( .IN1(inq_in2[3]), .IN2(n1879), .IN3(n1892), .IN4(n1689), .Q(
        \fpu_div_frac_dp/n1381 ) );
  AO22X1 U1617 ( .IN1(inq_in2[4]), .IN2(n1882), .IN3(n1892), .IN4(n1688), .Q(
        \fpu_div_frac_dp/n1380 ) );
  AO22X1 U1618 ( .IN1(inq_in2[5]), .IN2(n1881), .IN3(n1892), .IN4(n1687), .Q(
        \fpu_div_frac_dp/n1379 ) );
  AO22X1 U1619 ( .IN1(inq_in2[6]), .IN2(n1880), .IN3(n1892), .IN4(n1686), .Q(
        \fpu_div_frac_dp/n1378 ) );
  AO22X1 U1620 ( .IN1(inq_in2[7]), .IN2(n1879), .IN3(n1892), .IN4(n1710), .Q(
        \fpu_div_frac_dp/n1377 ) );
  AO22X1 U1621 ( .IN1(inq_in2[8]), .IN2(n1882), .IN3(n1892), .IN4(n1709), .Q(
        \fpu_div_frac_dp/n1376 ) );
  AO22X1 U1622 ( .IN1(inq_in2[9]), .IN2(n1881), .IN3(n1892), .IN4(n1639), .Q(
        \fpu_div_frac_dp/n1375 ) );
  AO22X1 U1623 ( .IN1(inq_in2[10]), .IN2(n1880), .IN3(n1892), .IN4(n1818), .Q(
        \fpu_div_frac_dp/n1374 ) );
  AO22X1 U1624 ( .IN1(inq_in2[11]), .IN2(n1879), .IN3(n1892), .IN4(n1708), .Q(
        \fpu_div_frac_dp/n1373 ) );
  AO22X1 U1625 ( .IN1(inq_in2[12]), .IN2(n1882), .IN3(n1892), .IN4(n1707), .Q(
        \fpu_div_frac_dp/n1372 ) );
  AO22X1 U1626 ( .IN1(inq_in2[13]), .IN2(n1881), .IN3(n1892), .IN4(n1706), .Q(
        \fpu_div_frac_dp/n1371 ) );
  AO22X1 U1627 ( .IN1(inq_in2[14]), .IN2(n1880), .IN3(n1892), .IN4(n1705), .Q(
        \fpu_div_frac_dp/n1370 ) );
  AO22X1 U1628 ( .IN1(inq_in2[15]), .IN2(n1879), .IN3(n1892), .IN4(n1704), .Q(
        \fpu_div_frac_dp/n1369 ) );
  AO22X1 U1629 ( .IN1(inq_in2[16]), .IN2(n1882), .IN3(n1892), .IN4(n1703), .Q(
        \fpu_div_frac_dp/n1368 ) );
  AO22X1 U1630 ( .IN1(inq_in2[17]), .IN2(n1881), .IN3(n1893), .IN4(n1702), .Q(
        \fpu_div_frac_dp/n1367 ) );
  AO22X1 U1631 ( .IN1(inq_in2[18]), .IN2(n1880), .IN3(n1893), .IN4(n1701), .Q(
        \fpu_div_frac_dp/n1366 ) );
  AO22X1 U1632 ( .IN1(inq_in2[19]), .IN2(n1879), .IN3(n1891), .IN4(n1700), .Q(
        \fpu_div_frac_dp/n1365 ) );
  AO22X1 U1633 ( .IN1(inq_in2[20]), .IN2(n1882), .IN3(n1893), .IN4(n1699), .Q(
        \fpu_div_frac_dp/n1364 ) );
  AO22X1 U1634 ( .IN1(inq_in2[21]), .IN2(n1881), .IN3(n1893), .IN4(n1698), .Q(
        \fpu_div_frac_dp/n1363 ) );
  AO22X1 U1635 ( .IN1(inq_in2[22]), .IN2(n1880), .IN3(n1893), .IN4(n1697), .Q(
        \fpu_div_frac_dp/n1362 ) );
  AO22X1 U1636 ( .IN1(inq_in2[23]), .IN2(n1879), .IN3(n1893), .IN4(n1696), .Q(
        \fpu_div_frac_dp/n1361 ) );
  AO22X1 U1637 ( .IN1(inq_in2[24]), .IN2(n1882), .IN3(n1893), .IN4(n1695), .Q(
        \fpu_div_frac_dp/n1360 ) );
  AO22X1 U1638 ( .IN1(inq_in2[25]), .IN2(n1881), .IN3(n1893), .IN4(n1694), .Q(
        \fpu_div_frac_dp/n1359 ) );
  AO22X1 U1639 ( .IN1(inq_in2[26]), .IN2(n1880), .IN3(n1893), .IN4(n1693), .Q(
        \fpu_div_frac_dp/n1358 ) );
  AO22X1 U1640 ( .IN1(inq_in2[27]), .IN2(n1879), .IN3(n1893), .IN4(n1692), .Q(
        \fpu_div_frac_dp/n1357 ) );
  AO22X1 U1641 ( .IN1(inq_in2[28]), .IN2(n1882), .IN3(n1893), .IN4(n1713), .Q(
        \fpu_div_frac_dp/n1356 ) );
  AO22X1 U1642 ( .IN1(inq_in2[29]), .IN2(n1881), .IN3(n1893), .IN4(n1714), .Q(
        \fpu_div_frac_dp/n1355 ) );
  AO22X1 U1643 ( .IN1(inq_in2[30]), .IN2(n1880), .IN3(n1893), .IN4(n1712), .Q(
        \fpu_div_frac_dp/n1354 ) );
  AO22X1 U1644 ( .IN1(inq_in2[31]), .IN2(n1879), .IN3(n1893), .IN4(n1711), .Q(
        \fpu_div_frac_dp/n1353 ) );
  AO22X1 U1645 ( .IN1(inq_in2[32]), .IN2(n1882), .IN3(n1894), .IN4(n1652), .Q(
        \fpu_div_frac_dp/n1352 ) );
  AO22X1 U1646 ( .IN1(inq_in2[33]), .IN2(n1881), .IN3(n1894), .IN4(n1669), .Q(
        \fpu_div_frac_dp/n1351 ) );
  AO22X1 U1647 ( .IN1(inq_in2[34]), .IN2(n1880), .IN3(n1893), .IN4(n1668), .Q(
        \fpu_div_frac_dp/n1350 ) );
  AO22X1 U1648 ( .IN1(inq_in2[35]), .IN2(n1879), .IN3(n1894), .IN4(n1667), .Q(
        \fpu_div_frac_dp/n1349 ) );
  AO22X1 U1649 ( .IN1(inq_in2[36]), .IN2(n1882), .IN3(n1894), .IN4(n1666), .Q(
        \fpu_div_frac_dp/n1348 ) );
  AO22X1 U1650 ( .IN1(inq_in2[37]), .IN2(n1881), .IN3(n1894), .IN4(n1665), .Q(
        \fpu_div_frac_dp/n1347 ) );
  AO22X1 U1651 ( .IN1(inq_in2[38]), .IN2(n1880), .IN3(n1894), .IN4(n1664), .Q(
        \fpu_div_frac_dp/n1346 ) );
  AO22X1 U1652 ( .IN1(inq_in2[39]), .IN2(n1879), .IN3(n1894), .IN4(n1663), .Q(
        \fpu_div_frac_dp/n1345 ) );
  AO22X1 U1653 ( .IN1(inq_in2[40]), .IN2(n1882), .IN3(n1894), .IN4(n1662), .Q(
        \fpu_div_frac_dp/n1344 ) );
  AO22X1 U1654 ( .IN1(inq_in2[41]), .IN2(n1881), .IN3(n1894), .IN4(n1661), .Q(
        \fpu_div_frac_dp/n1343 ) );
  AO22X1 U1655 ( .IN1(inq_in2[42]), .IN2(n1880), .IN3(n1894), .IN4(n1660), .Q(
        \fpu_div_frac_dp/n1342 ) );
  AO22X1 U1656 ( .IN1(inq_in2[43]), .IN2(n1879), .IN3(n1894), .IN4(n1659), .Q(
        \fpu_div_frac_dp/n1341 ) );
  AO22X1 U1657 ( .IN1(inq_in2[44]), .IN2(n1882), .IN3(n1894), .IN4(n1658), .Q(
        \fpu_div_frac_dp/n1340 ) );
  AO22X1 U1658 ( .IN1(inq_in2[45]), .IN2(n1881), .IN3(n1894), .IN4(n1657), .Q(
        \fpu_div_frac_dp/n1339 ) );
  AO22X1 U1659 ( .IN1(inq_in2[46]), .IN2(n1880), .IN3(n1894), .IN4(n1656), .Q(
        \fpu_div_frac_dp/n1338 ) );
  AO22X1 U1660 ( .IN1(inq_in2[47]), .IN2(n1879), .IN3(n1895), .IN4(n1655), .Q(
        \fpu_div_frac_dp/n1337 ) );
  AO22X1 U1661 ( .IN1(inq_in2[48]), .IN2(n1882), .IN3(n1895), .IN4(n1654), .Q(
        \fpu_div_frac_dp/n1336 ) );
  AO22X1 U1662 ( .IN1(inq_in2[49]), .IN2(n1881), .IN3(n1894), .IN4(n1653), .Q(
        \fpu_div_frac_dp/n1335 ) );
  AO22X1 U1663 ( .IN1(inq_in2[50]), .IN2(n1880), .IN3(n1895), .IN4(n1806), .Q(
        \fpu_div_frac_dp/n1334 ) );
  AO22X1 U1664 ( .IN1(n1879), .IN2(inq_in2[51]), .IN3(n1895), .IN4(n1671), .Q(
        \fpu_div_frac_dp/n1333 ) );
  AO22X1 U1665 ( .IN1(n1882), .IN2(inq_in2[52]), .IN3(n1895), .IN4(n1845), .Q(
        \fpu_div_frac_dp/n1332 ) );
  AO22X1 U1666 ( .IN1(n1881), .IN2(inq_in2[53]), .IN3(n1895), .IN4(n1849), .Q(
        \fpu_div_frac_dp/n1331 ) );
  AO22X1 U1667 ( .IN1(n1880), .IN2(inq_in2[54]), .IN3(n1888), .IN4(n1807), .Q(
        \fpu_div_frac_dp/n1330 ) );
  AO22X1 U1668 ( .IN1(n2189), .IN2(n1729), .IN3(n2217), .IN4(n2218), .Q(
        \fpu_div_frac_dp/n1329 ) );
  AO22X1 U1669 ( .IN1(n2189), .IN2(n1733), .IN3(n2217), .IN4(n2219), .Q(
        \fpu_div_frac_dp/n1328 ) );
  AO22X1 U1670 ( .IN1(n2189), .IN2(n1734), .IN3(n2220), .IN4(n2217), .Q(
        \fpu_div_frac_dp/n1327 ) );
  AO22X1 U1671 ( .IN1(n2189), .IN2(n1735), .IN3(n2217), .IN4(n2221), .Q(
        \fpu_div_frac_dp/n1326 ) );
  NOR2X0 U1672 ( .IN1(n2222), .IN2(n2223), .QN(n2217) );
  AO22X1 U1673 ( .IN1(n2189), .IN2(n1736), .IN3(n2224), .IN4(n2225), .Q(
        \fpu_div_frac_dp/n1325 ) );
  AO22X1 U1674 ( .IN1(n2189), .IN2(n1737), .IN3(n2224), .IN4(n2226), .Q(
        \fpu_div_frac_dp/n1324 ) );
  AO22X1 U1675 ( .IN1(n2189), .IN2(n1738), .IN3(n2224), .IN4(n2227), .Q(
        \fpu_div_frac_dp/n1323 ) );
  AO22X1 U1676 ( .IN1(n2189), .IN2(n1739), .IN3(n2224), .IN4(n2228), .Q(
        \fpu_div_frac_dp/n1322 ) );
  AO22X1 U1677 ( .IN1(n2189), .IN2(n1740), .IN3(n2224), .IN4(n2229), .Q(
        \fpu_div_frac_dp/n1321 ) );
  AO22X1 U1678 ( .IN1(n2189), .IN2(n1741), .IN3(n2224), .IN4(n2230), .Q(
        \fpu_div_frac_dp/n1320 ) );
  AO22X1 U1679 ( .IN1(n2189), .IN2(n1742), .IN3(n2224), .IN4(n2231), .Q(
        \fpu_div_frac_dp/n1319 ) );
  AO22X1 U1680 ( .IN1(n2189), .IN2(n1743), .IN3(n2224), .IN4(n2232), .Q(
        \fpu_div_frac_dp/n1318 ) );
  AO22X1 U1681 ( .IN1(n2189), .IN2(n1744), .IN3(n2224), .IN4(n2233), .Q(
        \fpu_div_frac_dp/n1317 ) );
  AO22X1 U1682 ( .IN1(n2189), .IN2(n1745), .IN3(n2224), .IN4(n2234), .Q(
        \fpu_div_frac_dp/n1316 ) );
  AO22X1 U1683 ( .IN1(n2189), .IN2(n1746), .IN3(n2224), .IN4(n2235), .Q(
        \fpu_div_frac_dp/n1315 ) );
  AO22X1 U1684 ( .IN1(n2189), .IN2(n1747), .IN3(n2224), .IN4(n2236), .Q(
        \fpu_div_frac_dp/n1314 ) );
  NOR2X0 U1685 ( .IN1(n2222), .IN2(n2237), .QN(n2224) );
  AO22X1 U1686 ( .IN1(n2189), .IN2(n1748), .IN3(n2238), .IN4(n2239), .Q(
        \fpu_div_frac_dp/n1313 ) );
  AO22X1 U1687 ( .IN1(n2189), .IN2(n1749), .IN3(n2238), .IN4(n2240), .Q(
        \fpu_div_frac_dp/n1312 ) );
  AO22X1 U1688 ( .IN1(n2189), .IN2(n1750), .IN3(n2238), .IN4(n2241), .Q(
        \fpu_div_frac_dp/n1311 ) );
  AO22X1 U1689 ( .IN1(n2189), .IN2(n1751), .IN3(n2238), .IN4(n2242), .Q(
        \fpu_div_frac_dp/n1310 ) );
  AO22X1 U1690 ( .IN1(n2189), .IN2(n1752), .IN3(n2238), .IN4(n2243), .Q(
        \fpu_div_frac_dp/n1309 ) );
  AO22X1 U1691 ( .IN1(n2189), .IN2(n1753), .IN3(n2244), .IN4(n2245), .Q(
        \fpu_div_frac_dp/n1308 ) );
  INVX0 U1692 ( .INP(n2246), .ZN(n2245) );
  AO22X1 U1693 ( .IN1(n2189), .IN2(n1754), .IN3(n2244), .IN4(n2247), .Q(
        \fpu_div_frac_dp/n1307 ) );
  INVX0 U1694 ( .INP(n2248), .ZN(n2247) );
  AO22X1 U1695 ( .IN1(n2189), .IN2(n1755), .IN3(n2244), .IN4(n2249), .Q(
        \fpu_div_frac_dp/n1306 ) );
  INVX0 U1696 ( .INP(n2250), .ZN(n2249) );
  AO22X1 U1697 ( .IN1(n2189), .IN2(n1756), .IN3(n2244), .IN4(n2251), .Q(
        \fpu_div_frac_dp/n1305 ) );
  INVX0 U1698 ( .INP(n2252), .ZN(n2251) );
  AO22X1 U1699 ( .IN1(n2189), .IN2(n1757), .IN3(n2244), .IN4(n2253), .Q(
        \fpu_div_frac_dp/n1304 ) );
  INVX0 U1700 ( .INP(n2254), .ZN(n2253) );
  AO22X1 U1701 ( .IN1(n2189), .IN2(n1758), .IN3(n2244), .IN4(n2255), .Q(
        \fpu_div_frac_dp/n1303 ) );
  INVX0 U1702 ( .INP(n2256), .ZN(n2255) );
  AO22X1 U1703 ( .IN1(n2189), .IN2(n1759), .IN3(n2244), .IN4(n2257), .Q(
        \fpu_div_frac_dp/n1302 ) );
  INVX0 U1704 ( .INP(n2258), .ZN(n2257) );
  AO22X1 U1705 ( .IN1(n2189), .IN2(n1760), .IN3(n2244), .IN4(n2259), .Q(
        \fpu_div_frac_dp/n1301 ) );
  INVX0 U1706 ( .INP(n2260), .ZN(n2259) );
  AO22X1 U1707 ( .IN1(n2189), .IN2(n1761), .IN3(n2244), .IN4(n2261), .Q(
        \fpu_div_frac_dp/n1300 ) );
  INVX0 U1708 ( .INP(n2262), .ZN(n2261) );
  AO22X1 U1709 ( .IN1(n2189), .IN2(n1762), .IN3(n2244), .IN4(n2263), .Q(
        \fpu_div_frac_dp/n1299 ) );
  INVX0 U1710 ( .INP(n2264), .ZN(n2263) );
  AO22X1 U1711 ( .IN1(n2189), .IN2(n1763), .IN3(n2244), .IN4(n2265), .Q(
        \fpu_div_frac_dp/n1298 ) );
  INVX0 U1712 ( .INP(n2266), .ZN(n2265) );
  AO22X1 U1713 ( .IN1(n2189), .IN2(n1764), .IN3(n2244), .IN4(n2267), .Q(
        \fpu_div_frac_dp/n1297 ) );
  AO22X1 U1714 ( .IN1(n2189), .IN2(n1765), .IN3(n2244), .IN4(n2268), .Q(
        \fpu_div_frac_dp/n1296 ) );
  AO22X1 U1715 ( .IN1(n2189), .IN2(n1766), .IN3(n2244), .IN4(n2269), .Q(
        \fpu_div_frac_dp/n1295 ) );
  AO22X1 U1716 ( .IN1(n2189), .IN2(n1767), .IN3(n2244), .IN4(n2270), .Q(
        \fpu_div_frac_dp/n1294 ) );
  AO22X1 U1717 ( .IN1(n2189), .IN2(n1768), .IN3(n2244), .IN4(n2271), .Q(
        \fpu_div_frac_dp/n1293 ) );
  AO22X1 U1718 ( .IN1(n2189), .IN2(n1769), .IN3(n2244), .IN4(n2272), .Q(
        \fpu_div_frac_dp/n1292 ) );
  AO22X1 U1719 ( .IN1(n2189), .IN2(n1770), .IN3(n2244), .IN4(n2273), .Q(
        \fpu_div_frac_dp/n1291 ) );
  AO22X1 U1720 ( .IN1(n2189), .IN2(n1771), .IN3(n2244), .IN4(n2274), .Q(
        \fpu_div_frac_dp/n1290 ) );
  AO22X1 U1721 ( .IN1(n2189), .IN2(n1772), .IN3(n2244), .IN4(n2275), .Q(
        \fpu_div_frac_dp/n1289 ) );
  AO22X1 U1722 ( .IN1(n2189), .IN2(n1773), .IN3(n2244), .IN4(n2276), .Q(
        \fpu_div_frac_dp/n1288 ) );
  AO22X1 U1723 ( .IN1(n2189), .IN2(n1774), .IN3(n2244), .IN4(n2277), .Q(
        \fpu_div_frac_dp/n1287 ) );
  AO22X1 U1724 ( .IN1(n2189), .IN2(n1775), .IN3(n2244), .IN4(n2278), .Q(
        \fpu_div_frac_dp/n1286 ) );
  AO22X1 U1725 ( .IN1(n2189), .IN2(n1776), .IN3(n2244), .IN4(n2279), .Q(
        \fpu_div_frac_dp/n1285 ) );
  AO22X1 U1726 ( .IN1(n2189), .IN2(n1777), .IN3(n2244), .IN4(n2280), .Q(
        \fpu_div_frac_dp/n1284 ) );
  AO22X1 U1727 ( .IN1(n2189), .IN2(n1778), .IN3(n2244), .IN4(n2281), .Q(
        \fpu_div_frac_dp/n1283 ) );
  AO22X1 U1728 ( .IN1(n2189), .IN2(n1779), .IN3(n2244), .IN4(n2282), .Q(
        \fpu_div_frac_dp/n1282 ) );
  AO22X1 U1729 ( .IN1(n2189), .IN2(n1780), .IN3(n2244), .IN4(n2283), .Q(
        \fpu_div_frac_dp/n1281 ) );
  AO222X1 U1730 ( .IN1(n2238), .IN2(n2284), .IN3(n2285), .IN4(n2240), .IN5(
        n2189), .IN6(n1726), .Q(\fpu_div_frac_dp/n1280 ) );
  AO222X1 U1731 ( .IN1(n2238), .IN2(n2286), .IN3(n2285), .IN4(n2241), .IN5(
        n2189), .IN6(n1727), .Q(\fpu_div_frac_dp/n1279 ) );
  AO222X1 U1732 ( .IN1(n2238), .IN2(n2287), .IN3(n2285), .IN4(n2242), .IN5(
        n2189), .IN6(n1728), .Q(\fpu_div_frac_dp/n1278 ) );
  AO222X1 U1733 ( .IN1(n2238), .IN2(n2288), .IN3(n2285), .IN4(n2243), .IN5(
        n2189), .IN6(n1718), .Q(\fpu_div_frac_dp/n1277 ) );
  NOR2X0 U1734 ( .IN1(n2222), .IN2(\fpu_div_frac_dp/n978 ), .QN(n2285) );
  NOR2X0 U1735 ( .IN1(n2222), .IN2(n1540), .QN(n2238) );
  INVX0 U1736 ( .INP(n2244), .ZN(n2222) );
  NOR2X0 U1737 ( .IN1(n2189), .IN2(se), .QN(n2244) );
  AND2X1 U1738 ( .IN1(n184), .IN2(n1047), .Q(n2189) );
  AO221X1 U1739 ( .IN1(n1883), .IN2(n2289), .IN3(n2290), .IN4(n1683), .IN5(
        n2291), .Q(\fpu_div_frac_dp/n1275 ) );
  AO21X1 U1740 ( .IN1(n2010), .IN2(n1397), .IN3(n2292), .Q(n2291) );
  AO221X1 U1741 ( .IN1(n2293), .IN2(n1883), .IN3(n2290), .IN4(n1437), .IN5(
        n2292), .Q(\fpu_div_frac_dp/n1274 ) );
  INVX0 U1742 ( .INP(n2219), .ZN(n2293) );
  AO221X1 U1743 ( .IN1(n1886), .IN2(n2294), .IN3(n2290), .IN4(n1436), .IN5(
        n2292), .Q(\fpu_div_frac_dp/n1273 ) );
  AO221X1 U1744 ( .IN1(n2295), .IN2(n1886), .IN3(n2290), .IN4(n1435), .IN5(
        n2292), .Q(\fpu_div_frac_dp/n1272 ) );
  AND2X1 U1745 ( .IN1(n1885), .IN2(n2223), .Q(n2292) );
  INVX0 U1746 ( .INP(n2221), .ZN(n2295) );
  AO221X1 U1747 ( .IN1(n1884), .IN2(n2296), .IN3(n2290), .IN4(n1434), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1271 ) );
  AO221X1 U1748 ( .IN1(n2298), .IN2(n1884), .IN3(n2290), .IN4(n1459), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1270 ) );
  AO221X1 U1749 ( .IN1(n2299), .IN2(n1885), .IN3(n2290), .IN4(n1458), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1269 ) );
  AO221X1 U1750 ( .IN1(n2300), .IN2(n1883), .IN3(n2290), .IN4(n1457), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1268 ) );
  AO221X1 U1751 ( .IN1(n2301), .IN2(n1886), .IN3(n2290), .IN4(n1456), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1267 ) );
  AO221X1 U1752 ( .IN1(n2302), .IN2(n1884), .IN3(n2290), .IN4(n1455), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1266 ) );
  AO221X1 U1753 ( .IN1(n2303), .IN2(n1885), .IN3(n2290), .IN4(n1454), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1265 ) );
  AO221X1 U1754 ( .IN1(n2304), .IN2(n1883), .IN3(n2290), .IN4(n1453), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1264 ) );
  AO221X1 U1755 ( .IN1(n2305), .IN2(n1886), .IN3(n2290), .IN4(n1452), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1263 ) );
  AO221X1 U1756 ( .IN1(n2306), .IN2(n1884), .IN3(n2290), .IN4(n1451), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1262 ) );
  AO221X1 U1757 ( .IN1(n2307), .IN2(n1885), .IN3(n2290), .IN4(n1450), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1261 ) );
  AO221X1 U1758 ( .IN1(n2308), .IN2(n1883), .IN3(n2290), .IN4(n1449), .IN5(
        n2297), .Q(\fpu_div_frac_dp/n1260 ) );
  AND2X1 U1759 ( .IN1(n1883), .IN2(n2237), .Q(n2297) );
  AO221X1 U1760 ( .IN1(n2309), .IN2(n1886), .IN3(n2290), .IN4(n1448), .IN5(
        n2310), .Q(\fpu_div_frac_dp/n1259 ) );
  INVX0 U1761 ( .INP(n2239), .ZN(n2309) );
  AO221X1 U1762 ( .IN1(n2311), .IN2(n1884), .IN3(n2290), .IN4(n1447), .IN5(
        n2310), .Q(\fpu_div_frac_dp/n1258 ) );
  AO221X1 U1763 ( .IN1(n2312), .IN2(n1883), .IN3(n2290), .IN4(n1446), .IN5(
        n2310), .Q(\fpu_div_frac_dp/n1257 ) );
  AO221X1 U1764 ( .IN1(n2313), .IN2(n1886), .IN3(n2290), .IN4(n1445), .IN5(
        n2310), .Q(\fpu_div_frac_dp/n1256 ) );
  AO221X1 U1765 ( .IN1(n2314), .IN2(n1884), .IN3(n2290), .IN4(n1444), .IN5(
        n2310), .Q(\fpu_div_frac_dp/n1255 ) );
  AO22X1 U1766 ( .IN1(n2290), .IN2(n1632), .IN3(n2246), .IN4(n1885), .Q(
        \fpu_div_frac_dp/n1254 ) );
  OA22X1 U1767 ( .IN1(n2237), .IN2(n2315), .IN3(n2316), .IN4(n2298), .Q(n2246)
         );
  AO22X1 U1768 ( .IN1(n2290), .IN2(n1631), .IN3(n2248), .IN4(n1883), .Q(
        \fpu_div_frac_dp/n1253 ) );
  OA22X1 U1769 ( .IN1(n2237), .IN2(n2317), .IN3(n2316), .IN4(n2299), .Q(n2248)
         );
  AO22X1 U1770 ( .IN1(n2290), .IN2(n1630), .IN3(n2250), .IN4(n1886), .Q(
        \fpu_div_frac_dp/n1252 ) );
  OA22X1 U1771 ( .IN1(n2237), .IN2(n2318), .IN3(n2316), .IN4(n2300), .Q(n2250)
         );
  AO22X1 U1772 ( .IN1(n2290), .IN2(n1629), .IN3(n2252), .IN4(n1884), .Q(
        \fpu_div_frac_dp/n1251 ) );
  OA22X1 U1773 ( .IN1(n2237), .IN2(n2319), .IN3(n2316), .IN4(n2301), .Q(n2252)
         );
  AO22X1 U1774 ( .IN1(n2290), .IN2(n1628), .IN3(n2254), .IN4(n1885), .Q(
        \fpu_div_frac_dp/n1250 ) );
  OA22X1 U1775 ( .IN1(n2237), .IN2(n2320), .IN3(n2316), .IN4(n2302), .Q(n2254)
         );
  AO22X1 U1776 ( .IN1(n2290), .IN2(n1627), .IN3(n2256), .IN4(n1883), .Q(
        \fpu_div_frac_dp/n1249 ) );
  OA22X1 U1777 ( .IN1(n2237), .IN2(n2321), .IN3(n2316), .IN4(n2303), .Q(n2256)
         );
  AO22X1 U1778 ( .IN1(n2290), .IN2(n1626), .IN3(n2258), .IN4(n1886), .Q(
        \fpu_div_frac_dp/n1248 ) );
  OA22X1 U1779 ( .IN1(n2237), .IN2(n2322), .IN3(n2316), .IN4(n2304), .Q(n2258)
         );
  AO22X1 U1780 ( .IN1(n2290), .IN2(n1625), .IN3(n2260), .IN4(n1884), .Q(
        \fpu_div_frac_dp/n1247 ) );
  OA22X1 U1781 ( .IN1(n2237), .IN2(n2323), .IN3(n2316), .IN4(n2305), .Q(n2260)
         );
  AO222X1 U1782 ( .IN1(n2262), .IN2(n1885), .IN3(n2010), .IN4(d6stg_fdivs), 
        .IN5(n2290), .IN6(n1442), .Q(\fpu_div_frac_dp/n1246 ) );
  OA22X1 U1783 ( .IN1(n2237), .IN2(n2324), .IN3(n2316), .IN4(n2306), .Q(n2262)
         );
  AO22X1 U1784 ( .IN1(n2290), .IN2(n1624), .IN3(n2264), .IN4(n1885), .Q(
        \fpu_div_frac_dp/n1245 ) );
  OA22X1 U1785 ( .IN1(n2237), .IN2(n2325), .IN3(n2316), .IN4(n2307), .Q(n2264)
         );
  AO22X1 U1786 ( .IN1(n2290), .IN2(n1488), .IN3(n2266), .IN4(n1883), .Q(
        \fpu_div_frac_dp/n1244 ) );
  OA22X1 U1787 ( .IN1(n2237), .IN2(n2326), .IN3(n2316), .IN4(n2308), .Q(n2266)
         );
  INVX0 U1788 ( .INP(n2327), .ZN(n2237) );
  AO22X1 U1789 ( .IN1(n2290), .IN2(n1487), .IN3(n2328), .IN4(n1886), .Q(
        \fpu_div_frac_dp/n1243 ) );
  INVX0 U1790 ( .INP(n2267), .ZN(n2328) );
  AO222X1 U1791 ( .IN1(n2329), .IN2(n2330), .IN3(n2331), .IN4(n2218), .IN5(
        n2327), .IN6(n2332), .Q(n2267) );
  AO22X1 U1792 ( .IN1(n2290), .IN2(n1486), .IN3(n2333), .IN4(n1884), .Q(
        \fpu_div_frac_dp/n1242 ) );
  INVX0 U1793 ( .INP(n2268), .ZN(n2333) );
  AO222X1 U1794 ( .IN1(n2329), .IN2(n2334), .IN3(n2331), .IN4(n2219), .IN5(
        n2327), .IN6(n2335), .Q(n2268) );
  AO22X1 U1795 ( .IN1(n2290), .IN2(n1485), .IN3(n2336), .IN4(n1885), .Q(
        \fpu_div_frac_dp/n1241 ) );
  INVX0 U1796 ( .INP(n2269), .ZN(n2336) );
  AO222X1 U1797 ( .IN1(n2329), .IN2(n2337), .IN3(n2331), .IN4(n2220), .IN5(
        n2327), .IN6(n2338), .Q(n2269) );
  AO22X1 U1798 ( .IN1(n2290), .IN2(n1484), .IN3(n2339), .IN4(n1883), .Q(
        \fpu_div_frac_dp/n1240 ) );
  INVX0 U1799 ( .INP(n2270), .ZN(n2339) );
  AO222X1 U1800 ( .IN1(n2329), .IN2(n2340), .IN3(n2331), .IN4(n2221), .IN5(
        n2327), .IN6(n2341), .Q(n2270) );
  AND2X1 U1801 ( .IN1(n2342), .IN2(n1540), .Q(n2331) );
  AO22X1 U1802 ( .IN1(n2290), .IN2(n1483), .IN3(n2343), .IN4(n1886), .Q(
        \fpu_div_frac_dp/n1239 ) );
  INVX0 U1803 ( .INP(n2271), .ZN(n2343) );
  AO222X1 U1804 ( .IN1(n2329), .IN2(n2344), .IN3(n2345), .IN4(n2225), .IN5(
        n2327), .IN6(n2346), .Q(n2271) );
  AO22X1 U1805 ( .IN1(n2290), .IN2(n1482), .IN3(n2347), .IN4(n1884), .Q(
        \fpu_div_frac_dp/n1238 ) );
  INVX0 U1806 ( .INP(n2272), .ZN(n2347) );
  NAND2X0 U1807 ( .IN1(n2348), .IN2(n2349), .QN(n2272) );
  OA222X1 U1808 ( .IN1(n2350), .IN2(n2223), .IN3(n2315), .IN4(n2316), .IN5(
        n2298), .IN6(n2351), .Q(n2349) );
  INVX0 U1809 ( .INP(n2226), .ZN(n2298) );
  AO22X1 U1810 ( .IN1(n2352), .IN2(n2353), .IN3(n2354), .IN4(n2219), .Q(n2226)
         );
  AOI221X1 U1811 ( .IN1(n2354), .IN2(n2355), .IN3(n2356), .IN4(n2357), .IN5(
        n2358), .QN(n2315) );
  AO22X1 U1812 ( .IN1(n2359), .IN2(n2360), .IN3(n2352), .IN4(n2361), .Q(n2358)
         );
  OA222X1 U1813 ( .IN1(n2362), .IN2(n2363), .IN3(n2364), .IN4(n2365), .IN5(
        n2366), .IN6(n2367), .Q(n2348) );
  INVX0 U1814 ( .INP(n2368), .ZN(n2366) );
  AO22X1 U1815 ( .IN1(n2290), .IN2(n1481), .IN3(n2369), .IN4(n1885), .Q(
        \fpu_div_frac_dp/n1237 ) );
  INVX0 U1816 ( .INP(n2273), .ZN(n2369) );
  NAND2X0 U1817 ( .IN1(n2370), .IN2(n2371), .QN(n2273) );
  OA222X1 U1818 ( .IN1(n2372), .IN2(n2223), .IN3(n2299), .IN4(n2351), .IN5(
        n2317), .IN6(n2316), .Q(n2371) );
  AOI221X1 U1819 ( .IN1(n2354), .IN2(n2373), .IN3(n2356), .IN4(n2374), .IN5(
        n2375), .QN(n2317) );
  AO22X1 U1820 ( .IN1(n2359), .IN2(n2376), .IN3(n2352), .IN4(n2377), .Q(n2375)
         );
  INVX0 U1821 ( .INP(n2227), .ZN(n2299) );
  AO22X1 U1822 ( .IN1(n2352), .IN2(n2378), .IN3(n2354), .IN4(n2220), .Q(n2227)
         );
  OA222X1 U1823 ( .IN1(n2379), .IN2(n2363), .IN3(n2380), .IN4(n2365), .IN5(
        n2381), .IN6(n2367), .Q(n2370) );
  INVX0 U1824 ( .INP(n2382), .ZN(n2381) );
  AO22X1 U1825 ( .IN1(n2290), .IN2(n1480), .IN3(n2383), .IN4(n1883), .Q(
        \fpu_div_frac_dp/n1236 ) );
  INVX0 U1826 ( .INP(n2274), .ZN(n2383) );
  NAND2X0 U1827 ( .IN1(n2384), .IN2(n2385), .QN(n2274) );
  OA222X1 U1828 ( .IN1(n2386), .IN2(n2223), .IN3(n2318), .IN4(n2316), .IN5(
        n2300), .IN6(n2351), .Q(n2385) );
  INVX0 U1829 ( .INP(n2228), .ZN(n2300) );
  AO22X1 U1830 ( .IN1(n2352), .IN2(n2387), .IN3(n2354), .IN4(n2221), .Q(n2228)
         );
  AOI221X1 U1831 ( .IN1(n2354), .IN2(n2388), .IN3(n2356), .IN4(n2389), .IN5(
        n2390), .QN(n2318) );
  AO22X1 U1832 ( .IN1(n2359), .IN2(n2391), .IN3(n2352), .IN4(n2392), .Q(n2390)
         );
  OA222X1 U1833 ( .IN1(n2393), .IN2(n2363), .IN3(n2394), .IN4(n2365), .IN5(
        n2395), .IN6(n2367), .Q(n2384) );
  INVX0 U1834 ( .INP(n2396), .ZN(n2395) );
  AO22X1 U1835 ( .IN1(n2290), .IN2(n1479), .IN3(n2397), .IN4(n1886), .Q(
        \fpu_div_frac_dp/n1235 ) );
  INVX0 U1836 ( .INP(n2275), .ZN(n2397) );
  NAND2X0 U1837 ( .IN1(n2398), .IN2(n2399), .QN(n2275) );
  OA222X1 U1838 ( .IN1(n2400), .IN2(n2223), .IN3(n2319), .IN4(n2316), .IN5(
        n2301), .IN6(n2351), .Q(n2399) );
  INVX0 U1839 ( .INP(n2229), .ZN(n2301) );
  AO222X1 U1840 ( .IN1(n2356), .IN2(n2218), .IN3(n2354), .IN4(n2401), .IN5(
        n2352), .IN6(n2402), .Q(n2229) );
  AOI221X1 U1841 ( .IN1(n2352), .IN2(n2403), .IN3(n2356), .IN4(n2404), .IN5(
        n2405), .QN(n2319) );
  AO22X1 U1842 ( .IN1(n2359), .IN2(n2406), .IN3(n2354), .IN4(n2407), .Q(n2405)
         );
  OA222X1 U1843 ( .IN1(n2408), .IN2(n2363), .IN3(n2409), .IN4(n2365), .IN5(
        n2410), .IN6(n2367), .Q(n2398) );
  INVX0 U1844 ( .INP(n2411), .ZN(n2410) );
  AO22X1 U1845 ( .IN1(n2290), .IN2(n1478), .IN3(n2412), .IN4(n1884), .Q(
        \fpu_div_frac_dp/n1234 ) );
  INVX0 U1846 ( .INP(n2276), .ZN(n2412) );
  NAND2X0 U1847 ( .IN1(n2413), .IN2(n2414), .QN(n2276) );
  OA222X1 U1848 ( .IN1(n2415), .IN2(n2223), .IN3(n2320), .IN4(n2316), .IN5(
        n2302), .IN6(n2351), .Q(n2414) );
  INVX0 U1849 ( .INP(n2230), .ZN(n2302) );
  AO222X1 U1850 ( .IN1(n2352), .IN2(n2360), .IN3(n2356), .IN4(n2219), .IN5(
        n2354), .IN6(n2353), .Q(n2230) );
  AOI221X1 U1851 ( .IN1(n2352), .IN2(n2368), .IN3(n2354), .IN4(n2361), .IN5(
        n2416), .QN(n2320) );
  AO22X1 U1852 ( .IN1(n2356), .IN2(n2355), .IN3(n2359), .IN4(n2357), .Q(n2416)
         );
  OA222X1 U1853 ( .IN1(n2350), .IN2(n2363), .IN3(n2362), .IN4(n2365), .IN5(
        n2364), .IN6(n2367), .Q(n2413) );
  INVX0 U1854 ( .INP(n2417), .ZN(n2364) );
  AO22X1 U1855 ( .IN1(n2290), .IN2(n1477), .IN3(n2418), .IN4(n1885), .Q(
        \fpu_div_frac_dp/n1233 ) );
  INVX0 U1856 ( .INP(n2277), .ZN(n2418) );
  NAND2X0 U1857 ( .IN1(n2419), .IN2(n2420), .QN(n2277) );
  OA222X1 U1858 ( .IN1(n2421), .IN2(n2223), .IN3(n2321), .IN4(n2316), .IN5(
        n2303), .IN6(n2351), .Q(n2420) );
  INVX0 U1859 ( .INP(n2231), .ZN(n2303) );
  AO222X1 U1860 ( .IN1(n2352), .IN2(n2376), .IN3(n2356), .IN4(n2220), .IN5(
        n2354), .IN6(n2378), .Q(n2231) );
  AOI221X1 U1861 ( .IN1(n2352), .IN2(n2382), .IN3(n2354), .IN4(n2377), .IN5(
        n2422), .QN(n2321) );
  AO22X1 U1862 ( .IN1(n2356), .IN2(n2373), .IN3(n2359), .IN4(n2374), .Q(n2422)
         );
  OA222X1 U1863 ( .IN1(n2372), .IN2(n2363), .IN3(n2379), .IN4(n2365), .IN5(
        n2380), .IN6(n2367), .Q(n2419) );
  INVX0 U1864 ( .INP(n2423), .ZN(n2380) );
  AO22X1 U1865 ( .IN1(n2290), .IN2(n1476), .IN3(n2424), .IN4(n1883), .Q(
        \fpu_div_frac_dp/n1232 ) );
  INVX0 U1866 ( .INP(n2278), .ZN(n2424) );
  NAND2X0 U1867 ( .IN1(n2425), .IN2(n2426), .QN(n2278) );
  OA222X1 U1868 ( .IN1(n2427), .IN2(n2223), .IN3(n2322), .IN4(n2316), .IN5(
        n2304), .IN6(n2351), .Q(n2426) );
  INVX0 U1869 ( .INP(n2232), .ZN(n2304) );
  AO222X1 U1870 ( .IN1(n2352), .IN2(n2391), .IN3(n2356), .IN4(n2221), .IN5(
        n2354), .IN6(n2387), .Q(n2232) );
  AOI221X1 U1871 ( .IN1(n2352), .IN2(n2396), .IN3(n2354), .IN4(n2392), .IN5(
        n2428), .QN(n2322) );
  AO22X1 U1872 ( .IN1(n2356), .IN2(n2388), .IN3(n2359), .IN4(n2389), .Q(n2428)
         );
  OA222X1 U1873 ( .IN1(n2386), .IN2(n2363), .IN3(n2393), .IN4(n2365), .IN5(
        n2394), .IN6(n2367), .Q(n2425) );
  INVX0 U1874 ( .INP(n2429), .ZN(n2394) );
  AO22X1 U1875 ( .IN1(n2290), .IN2(n1475), .IN3(n2430), .IN4(n1886), .Q(
        \fpu_div_frac_dp/n1231 ) );
  INVX0 U1876 ( .INP(n2279), .ZN(n2430) );
  NAND2X0 U1877 ( .IN1(n2431), .IN2(n2432), .QN(n2279) );
  OA222X1 U1878 ( .IN1(n2433), .IN2(n2223), .IN3(n2305), .IN4(n2351), .IN5(
        n2323), .IN6(n2316), .Q(n2432) );
  AOI221X1 U1879 ( .IN1(n2352), .IN2(n2411), .IN3(n2354), .IN4(n2403), .IN5(
        n2434), .QN(n2323) );
  AO22X1 U1880 ( .IN1(n2359), .IN2(n2404), .IN3(n2356), .IN4(n2407), .Q(n2434)
         );
  INVX0 U1881 ( .INP(n2233), .ZN(n2305) );
  AO221X1 U1882 ( .IN1(n2352), .IN2(n2406), .IN3(n2354), .IN4(n2402), .IN5(
        n2435), .Q(n2233) );
  AO22X1 U1883 ( .IN1(n2359), .IN2(n2218), .IN3(n2356), .IN4(n2401), .Q(n2435)
         );
  OA222X1 U1884 ( .IN1(n2400), .IN2(n2363), .IN3(n2408), .IN4(n2365), .IN5(
        n2409), .IN6(n2367), .Q(n2431) );
  INVX0 U1885 ( .INP(n2436), .ZN(n2409) );
  AO22X1 U1886 ( .IN1(n2290), .IN2(n1474), .IN3(n2437), .IN4(n1884), .Q(
        \fpu_div_frac_dp/n1230 ) );
  INVX0 U1887 ( .INP(n2280), .ZN(n2437) );
  NAND2X0 U1888 ( .IN1(n2438), .IN2(n2439), .QN(n2280) );
  OA222X1 U1889 ( .IN1(n2440), .IN2(n2223), .IN3(n2306), .IN4(n2351), .IN5(
        n2324), .IN6(n2316), .Q(n2439) );
  AOI221X1 U1890 ( .IN1(n2354), .IN2(n2368), .IN3(n2356), .IN4(n2361), .IN5(
        n2441), .QN(n2324) );
  AO22X1 U1891 ( .IN1(n2359), .IN2(n2355), .IN3(n2352), .IN4(n2417), .Q(n2441)
         );
  INVX0 U1892 ( .INP(n2234), .ZN(n2306) );
  AO221X1 U1893 ( .IN1(n2359), .IN2(n2219), .IN3(n2354), .IN4(n2360), .IN5(
        n2442), .Q(n2234) );
  AO22X1 U1894 ( .IN1(n2352), .IN2(n2357), .IN3(n2356), .IN4(n2353), .Q(n2442)
         );
  INVX0 U1895 ( .INP(n2443), .ZN(n2440) );
  OA222X1 U1896 ( .IN1(n2415), .IN2(n2363), .IN3(n2350), .IN4(n2365), .IN5(
        n2362), .IN6(n2367), .Q(n2438) );
  INVX0 U1897 ( .INP(n2444), .ZN(n2362) );
  INVX0 U1898 ( .INP(n2445), .ZN(n2350) );
  INVX0 U1899 ( .INP(n2446), .ZN(n2415) );
  AO22X1 U1900 ( .IN1(n2290), .IN2(n1473), .IN3(n2447), .IN4(n1885), .Q(
        \fpu_div_frac_dp/n1229 ) );
  INVX0 U1901 ( .INP(n2281), .ZN(n2447) );
  NAND2X0 U1902 ( .IN1(n2448), .IN2(n2449), .QN(n2281) );
  OA222X1 U1903 ( .IN1(n2450), .IN2(n2223), .IN3(n2307), .IN4(n2351), .IN5(
        n2325), .IN6(n2316), .Q(n2449) );
  AOI221X1 U1904 ( .IN1(n2354), .IN2(n2382), .IN3(n2356), .IN4(n2377), .IN5(
        n2451), .QN(n2325) );
  AO22X1 U1905 ( .IN1(n2359), .IN2(n2373), .IN3(n2352), .IN4(n2423), .Q(n2451)
         );
  INVX0 U1906 ( .INP(n2235), .ZN(n2307) );
  AO221X1 U1907 ( .IN1(n2359), .IN2(n2220), .IN3(n2354), .IN4(n2376), .IN5(
        n2452), .Q(n2235) );
  AO22X1 U1908 ( .IN1(n2352), .IN2(n2374), .IN3(n2356), .IN4(n2378), .Q(n2452)
         );
  INVX0 U1909 ( .INP(n2453), .ZN(n2450) );
  OA222X1 U1910 ( .IN1(n2421), .IN2(n2363), .IN3(n2372), .IN4(n2365), .IN5(
        n2379), .IN6(n2367), .Q(n2448) );
  INVX0 U1911 ( .INP(n2454), .ZN(n2379) );
  INVX0 U1912 ( .INP(n2455), .ZN(n2372) );
  INVX0 U1913 ( .INP(n2456), .ZN(n2421) );
  AO22X1 U1914 ( .IN1(n2290), .IN2(n1472), .IN3(n2457), .IN4(n1884), .Q(
        \fpu_div_frac_dp/n1228 ) );
  INVX0 U1915 ( .INP(n2282), .ZN(n2457) );
  NAND2X0 U1916 ( .IN1(n2458), .IN2(n2459), .QN(n2282) );
  OA222X1 U1917 ( .IN1(n2460), .IN2(n2223), .IN3(n2308), .IN4(n2351), .IN5(
        n2326), .IN6(n2316), .Q(n2459) );
  INVX0 U1918 ( .INP(n2329), .ZN(n2316) );
  AOI221X1 U1919 ( .IN1(n2354), .IN2(n2396), .IN3(n2356), .IN4(n2392), .IN5(
        n2461), .QN(n2326) );
  AO22X1 U1920 ( .IN1(n2359), .IN2(n2388), .IN3(n2352), .IN4(n2429), .Q(n2461)
         );
  INVX0 U1921 ( .INP(n2345), .ZN(n2351) );
  NOR2X0 U1922 ( .IN1(n1392), .IN2(\fpu_div_frac_dp/n978 ), .QN(n2345) );
  INVX0 U1923 ( .INP(n2236), .ZN(n2308) );
  AO221X1 U1924 ( .IN1(n2359), .IN2(n2221), .IN3(n2354), .IN4(n2391), .IN5(
        n2462), .Q(n2236) );
  AO22X1 U1925 ( .IN1(n2352), .IN2(n2389), .IN3(n2356), .IN4(n2387), .Q(n2462)
         );
  INVX0 U1926 ( .INP(n2463), .ZN(n2460) );
  OA222X1 U1927 ( .IN1(n2427), .IN2(n2363), .IN3(n2386), .IN4(n2365), .IN5(
        n2393), .IN6(n2367), .Q(n2458) );
  INVX0 U1928 ( .INP(n2464), .ZN(n2393) );
  INVX0 U1929 ( .INP(n2465), .ZN(n2386) );
  INVX0 U1930 ( .INP(n2466), .ZN(n2427) );
  AO22X1 U1931 ( .IN1(n2290), .IN2(n1471), .IN3(n2467), .IN4(n1885), .Q(
        \fpu_div_frac_dp/n1227 ) );
  INVX0 U1932 ( .INP(n2283), .ZN(n2467) );
  NAND2X0 U1933 ( .IN1(n2468), .IN2(n2469), .QN(n2283) );
  AOI222X1 U1934 ( .IN1(n1540), .IN2(n2239), .IN3(n2332), .IN4(n2329), .IN5(
        n2470), .IN6(n2471), .QN(n2469) );
  INVX0 U1935 ( .INP(n2223), .ZN(n2471) );
  NAND2X0 U1936 ( .IN1(n2352), .IN2(n2327), .QN(n2223) );
  NOR2X0 U1937 ( .IN1(n1540), .IN2(\fpu_div_frac_dp/n967 ), .QN(n2329) );
  AO221X1 U1938 ( .IN1(n2354), .IN2(n2411), .IN3(n2356), .IN4(n2403), .IN5(
        n2472), .Q(n2332) );
  AO22X1 U1939 ( .IN1(n2359), .IN2(n2407), .IN3(n2352), .IN4(n2436), .Q(n2472)
         );
  AO22X1 U1940 ( .IN1(\fpu_div_frac_dp/n967 ), .IN2(n2330), .IN3(n2473), .IN4(
        n2218), .Q(n2239) );
  AO221X1 U1941 ( .IN1(n2359), .IN2(n2401), .IN3(n2354), .IN4(n2406), .IN5(
        n2474), .Q(n2330) );
  AO22X1 U1942 ( .IN1(n2352), .IN2(n2404), .IN3(n2356), .IN4(n2402), .Q(n2474)
         );
  OA222X1 U1943 ( .IN1(n2433), .IN2(n2363), .IN3(n2400), .IN4(n2365), .IN5(
        n2408), .IN6(n2367), .Q(n2468) );
  NAND2X0 U1944 ( .IN1(n2359), .IN2(n2327), .QN(n2367) );
  INVX0 U1945 ( .INP(n2475), .ZN(n2408) );
  NAND2X0 U1946 ( .IN1(n2356), .IN2(n2327), .QN(n2365) );
  INVX0 U1947 ( .INP(n2476), .ZN(n2400) );
  NAND2X0 U1948 ( .IN1(n2354), .IN2(n2327), .QN(n2363) );
  NOR2X0 U1949 ( .IN1(n1540), .IN2(n1392), .QN(n2327) );
  INVX0 U1950 ( .INP(n2477), .ZN(n2433) );
  AO222X1 U1951 ( .IN1(n2310), .IN2(n2311), .IN3(n2478), .IN4(n2479), .IN5(
        n2290), .IN6(n1441), .Q(\fpu_div_frac_dp/n1226 ) );
  INVX0 U1952 ( .INP(n2284), .ZN(n2479) );
  AO21X1 U1953 ( .IN1(n2342), .IN2(n2480), .IN3(n2481), .Q(n2284) );
  MUX21X1 U1954 ( .IN1(n2482), .IN2(n2335), .S(n1392), .Q(n2481) );
  AO221X1 U1955 ( .IN1(n2354), .IN2(n2417), .IN3(n2352), .IN4(n2444), .IN5(
        n2483), .Q(n2335) );
  AO22X1 U1956 ( .IN1(n2359), .IN2(n2361), .IN3(n2356), .IN4(n2368), .Q(n2483)
         );
  AO221X1 U1957 ( .IN1(n2484), .IN2(n1555), .IN3(n2485), .IN4(n1414), .IN5(
        n2486), .Q(n2368) );
  AO22X1 U1958 ( .IN1(n2487), .IN2(n1413), .IN3(n2488), .IN4(n1554), .Q(n2486)
         );
  AO221X1 U1959 ( .IN1(n2484), .IN2(n1571), .IN3(n2485), .IN4(n1430), .IN5(
        n2489), .Q(n2361) );
  AO22X1 U1960 ( .IN1(n2487), .IN2(n1429), .IN3(n2488), .IN4(n1556), .Q(n2489)
         );
  AO221X1 U1961 ( .IN1(n2484), .IN2(n1559), .IN3(n2485), .IN4(n1418), .IN5(
        n2490), .Q(n2444) );
  AO22X1 U1962 ( .IN1(n2487), .IN2(n1417), .IN3(n2488), .IN4(n1558), .Q(n2490)
         );
  AO221X1 U1963 ( .IN1(n2484), .IN2(n1553), .IN3(n2485), .IN4(n1412), .IN5(
        n2491), .Q(n2417) );
  AO22X1 U1964 ( .IN1(n2487), .IN2(n1411), .IN3(n2488), .IN4(n1560), .Q(n2491)
         );
  AO222X1 U1965 ( .IN1(n2354), .IN2(n2443), .IN3(n2356), .IN4(n2446), .IN5(
        n2359), .IN6(n2445), .Q(n2482) );
  AO221X1 U1966 ( .IN1(n2484), .IN2(n1557), .IN3(n2485), .IN4(n1416), .IN5(
        n2492), .Q(n2445) );
  AO22X1 U1967 ( .IN1(n2487), .IN2(n1415), .IN3(n2488), .IN4(n1562), .Q(n2492)
         );
  AO221X1 U1968 ( .IN1(n2484), .IN2(n1561), .IN3(n2485), .IN4(n1420), .IN5(
        n2493), .Q(n2446) );
  AO22X1 U1969 ( .IN1(n2487), .IN2(n1419), .IN3(n2488), .IN4(n1564), .Q(n2493)
         );
  AO221X1 U1970 ( .IN1(n2484), .IN2(n1563), .IN3(n2485), .IN4(n1422), .IN5(
        n2494), .Q(n2443) );
  AO22X1 U1971 ( .IN1(n2487), .IN2(n1421), .IN3(n2488), .IN4(n1566), .Q(n2494)
         );
  AO221X1 U1972 ( .IN1(n2484), .IN2(n1565), .IN3(n2485), .IN4(n1424), .IN5(
        n2495), .Q(n2480) );
  AO22X1 U1973 ( .IN1(n2487), .IN2(n1423), .IN3(n2488), .IN4(n1567), .Q(n2495)
         );
  INVX0 U1974 ( .INP(n2240), .ZN(n2311) );
  AO22X1 U1975 ( .IN1(\fpu_div_frac_dp/n967 ), .IN2(n2334), .IN3(n2473), .IN4(
        n2219), .Q(n2240) );
  AO22X1 U1976 ( .IN1(n2488), .IN2(n1533), .IN3(n2485), .IN4(n1646), .Q(n2219)
         );
  AO221X1 U1977 ( .IN1(n2354), .IN2(n2357), .IN3(n2352), .IN4(n2355), .IN5(
        n2496), .Q(n2334) );
  AO22X1 U1978 ( .IN1(n2359), .IN2(n2353), .IN3(n2356), .IN4(n2360), .Q(n2496)
         );
  AO221X1 U1979 ( .IN1(n2484), .IN2(n1427), .IN3(n2485), .IN4(n1570), .IN5(
        n2497), .Q(n2360) );
  AO22X1 U1980 ( .IN1(n2487), .IN2(n1569), .IN3(n2488), .IN4(n1426), .Q(n2497)
         );
  AO221X1 U1981 ( .IN1(n2484), .IN2(n1425), .IN3(n2485), .IN4(n1568), .IN5(
        n2498), .Q(n2353) );
  AO22X1 U1982 ( .IN1(n2487), .IN2(n1638), .IN3(n2488), .IN4(n1428), .Q(n2498)
         );
  AO221X1 U1983 ( .IN1(n2484), .IN2(n1573), .IN3(n2485), .IN4(n1432), .IN5(
        n2499), .Q(n2355) );
  AO22X1 U1984 ( .IN1(n2487), .IN2(n1431), .IN3(n2488), .IN4(n1572), .Q(n2499)
         );
  AO221X1 U1985 ( .IN1(n2484), .IN2(n1370), .IN3(n2485), .IN4(n1385), .IN5(
        n2500), .Q(n2357) );
  AO22X1 U1986 ( .IN1(n2487), .IN2(n1384), .IN3(n2488), .IN4(n1574), .Q(n2500)
         );
  AO222X1 U1987 ( .IN1(n2310), .IN2(n2312), .IN3(n2501), .IN4(n2478), .IN5(
        n2290), .IN6(n1440), .Q(\fpu_div_frac_dp/n1225 ) );
  INVX0 U1988 ( .INP(n2286), .ZN(n2501) );
  AO21X1 U1989 ( .IN1(n2342), .IN2(n2502), .IN3(n2503), .Q(n2286) );
  MUX21X1 U1990 ( .IN1(n2504), .IN2(n2338), .S(n1392), .Q(n2503) );
  AO221X1 U1991 ( .IN1(n2354), .IN2(n2423), .IN3(n2352), .IN4(n2454), .IN5(
        n2505), .Q(n2338) );
  AO22X1 U1992 ( .IN1(n2359), .IN2(n2377), .IN3(n2356), .IN4(n2382), .Q(n2505)
         );
  AO221X1 U1993 ( .IN1(n2484), .IN2(n1414), .IN3(n2485), .IN4(n1554), .IN5(
        n2506), .Q(n2382) );
  AO22X1 U1994 ( .IN1(n2487), .IN2(n1555), .IN3(n2488), .IN4(n1411), .Q(n2506)
         );
  AO221X1 U1995 ( .IN1(n2484), .IN2(n1430), .IN3(n2485), .IN4(n1556), .IN5(
        n2507), .Q(n2377) );
  AO22X1 U1996 ( .IN1(n2487), .IN2(n1571), .IN3(n2488), .IN4(n1413), .Q(n2507)
         );
  AO221X1 U1997 ( .IN1(n2484), .IN2(n1418), .IN3(n2485), .IN4(n1558), .IN5(
        n2508), .Q(n2454) );
  AO22X1 U1998 ( .IN1(n2487), .IN2(n1559), .IN3(n2488), .IN4(n1415), .Q(n2508)
         );
  AO221X1 U1999 ( .IN1(n2484), .IN2(n1412), .IN3(n2485), .IN4(n1560), .IN5(
        n2509), .Q(n2423) );
  AO22X1 U2000 ( .IN1(n2487), .IN2(n1553), .IN3(n2488), .IN4(n1417), .Q(n2509)
         );
  AO222X1 U2001 ( .IN1(n2354), .IN2(n2453), .IN3(n2356), .IN4(n2456), .IN5(
        n2359), .IN6(n2455), .Q(n2504) );
  AO221X1 U2002 ( .IN1(n2484), .IN2(n1416), .IN3(n2485), .IN4(n1562), .IN5(
        n2510), .Q(n2455) );
  AO22X1 U2003 ( .IN1(n2487), .IN2(n1557), .IN3(n2488), .IN4(n1419), .Q(n2510)
         );
  AO221X1 U2004 ( .IN1(n2484), .IN2(n1420), .IN3(n2485), .IN4(n1564), .IN5(
        n2511), .Q(n2456) );
  AO22X1 U2005 ( .IN1(n2487), .IN2(n1561), .IN3(n2488), .IN4(n1421), .Q(n2511)
         );
  AO221X1 U2006 ( .IN1(n2484), .IN2(n1422), .IN3(n2485), .IN4(n1566), .IN5(
        n2512), .Q(n2453) );
  AO22X1 U2007 ( .IN1(n2487), .IN2(n1563), .IN3(n2488), .IN4(n1423), .Q(n2512)
         );
  AO221X1 U2008 ( .IN1(n2484), .IN2(n1424), .IN3(n2485), .IN4(n1567), .IN5(
        n2513), .Q(n2502) );
  AO22X1 U2009 ( .IN1(n2487), .IN2(n1565), .IN3(n2488), .IN4(n1530), .Q(n2513)
         );
  INVX0 U2010 ( .INP(n2241), .ZN(n2312) );
  AO22X1 U2011 ( .IN1(\fpu_div_frac_dp/n967 ), .IN2(n2337), .IN3(n2473), .IN4(
        n2220), .Q(n2241) );
  INVX0 U2012 ( .INP(n2294), .ZN(n2220) );
  AO221X1 U2013 ( .IN1(\fpu_div_frac_dp/n325 ), .IN2(n1398), .IN3(
        \fpu_div_frac_dp/n324 ), .IN4(n2488), .IN5(n2514), .Q(n2294) );
  AO21X1 U2014 ( .IN1(\fpu_div_frac_dp/n326 ), .IN2(n1544), .IN3(n2487), .Q(
        n2514) );
  AO221X1 U2015 ( .IN1(n2354), .IN2(n2374), .IN3(n2352), .IN4(n2373), .IN5(
        n2515), .Q(n2337) );
  AO22X1 U2016 ( .IN1(n2359), .IN2(n2378), .IN3(n2356), .IN4(n2376), .Q(n2515)
         );
  AO221X1 U2017 ( .IN1(n2484), .IN2(n1570), .IN3(n2485), .IN4(n1426), .IN5(
        n2516), .Q(n2376) );
  AO22X1 U2018 ( .IN1(n2487), .IN2(n1427), .IN3(n2488), .IN4(n1384), .Q(n2516)
         );
  AO221X1 U2019 ( .IN1(n2484), .IN2(n1568), .IN3(n2485), .IN4(n1428), .IN5(
        n2517), .Q(n2378) );
  AO22X1 U2020 ( .IN1(n2487), .IN2(n1425), .IN3(n2488), .IN4(n1569), .Q(n2517)
         );
  AO221X1 U2021 ( .IN1(n2484), .IN2(n1432), .IN3(n2485), .IN4(n1572), .IN5(
        n2518), .Q(n2373) );
  AO22X1 U2022 ( .IN1(n2487), .IN2(n1573), .IN3(n2488), .IN4(n1429), .Q(n2518)
         );
  AO221X1 U2023 ( .IN1(n2484), .IN2(n1385), .IN3(n2485), .IN4(n1574), .IN5(
        n2519), .Q(n2374) );
  AO22X1 U2024 ( .IN1(n2487), .IN2(n1370), .IN3(n2488), .IN4(n1431), .Q(n2519)
         );
  AO222X1 U2025 ( .IN1(n2310), .IN2(n2313), .IN3(n2520), .IN4(n2478), .IN5(
        n2290), .IN6(n1439), .Q(\fpu_div_frac_dp/n1224 ) );
  INVX0 U2026 ( .INP(n2287), .ZN(n2520) );
  AO21X1 U2027 ( .IN1(n2342), .IN2(n2521), .IN3(n2522), .Q(n2287) );
  MUX21X1 U2028 ( .IN1(n2523), .IN2(n2341), .S(n1392), .Q(n2522) );
  AO221X1 U2029 ( .IN1(n2354), .IN2(n2429), .IN3(n2352), .IN4(n2464), .IN5(
        n2524), .Q(n2341) );
  AO22X1 U2030 ( .IN1(n2359), .IN2(n2392), .IN3(n2356), .IN4(n2396), .Q(n2524)
         );
  AO221X1 U2031 ( .IN1(n2484), .IN2(n1554), .IN3(n2485), .IN4(n1411), .IN5(
        n2525), .Q(n2396) );
  AO22X1 U2032 ( .IN1(n2487), .IN2(n1414), .IN3(n2488), .IN4(n1553), .Q(n2525)
         );
  AO221X1 U2033 ( .IN1(n2484), .IN2(n1556), .IN3(n2485), .IN4(n1413), .IN5(
        n2526), .Q(n2392) );
  AO22X1 U2034 ( .IN1(n2487), .IN2(n1430), .IN3(n2488), .IN4(n1555), .Q(n2526)
         );
  AO221X1 U2035 ( .IN1(n2484), .IN2(n1558), .IN3(n2485), .IN4(n1415), .IN5(
        n2527), .Q(n2464) );
  AO22X1 U2036 ( .IN1(n2487), .IN2(n1418), .IN3(n2488), .IN4(n1557), .Q(n2527)
         );
  AO221X1 U2037 ( .IN1(n2484), .IN2(n1560), .IN3(n2485), .IN4(n1417), .IN5(
        n2528), .Q(n2429) );
  AO22X1 U2038 ( .IN1(n2487), .IN2(n1412), .IN3(n2488), .IN4(n1559), .Q(n2528)
         );
  AO222X1 U2039 ( .IN1(n2354), .IN2(n2463), .IN3(n2356), .IN4(n2466), .IN5(
        n2359), .IN6(n2465), .Q(n2523) );
  AO221X1 U2040 ( .IN1(n2484), .IN2(n1562), .IN3(n2485), .IN4(n1419), .IN5(
        n2529), .Q(n2465) );
  AO22X1 U2041 ( .IN1(n2487), .IN2(n1416), .IN3(n2488), .IN4(n1561), .Q(n2529)
         );
  AO221X1 U2042 ( .IN1(n2484), .IN2(n1564), .IN3(n2485), .IN4(n1421), .IN5(
        n2530), .Q(n2466) );
  AO22X1 U2043 ( .IN1(n2487), .IN2(n1420), .IN3(n2488), .IN4(n1563), .Q(n2530)
         );
  AO221X1 U2044 ( .IN1(n2484), .IN2(n1566), .IN3(n2485), .IN4(n1423), .IN5(
        n2531), .Q(n2463) );
  AO22X1 U2045 ( .IN1(n2487), .IN2(n1422), .IN3(n2488), .IN4(n1565), .Q(n2531)
         );
  AO221X1 U2046 ( .IN1(n2484), .IN2(n1567), .IN3(n2485), .IN4(n1530), .IN5(
        n2532), .Q(n2521) );
  AO22X1 U2047 ( .IN1(n2487), .IN2(n1424), .IN3(n2488), .IN4(n1721), .Q(n2532)
         );
  INVX0 U2048 ( .INP(n2242), .ZN(n2313) );
  AO22X1 U2049 ( .IN1(\fpu_div_frac_dp/n967 ), .IN2(n2340), .IN3(n2473), .IN4(
        n2221), .Q(n2242) );
  AO221X1 U2050 ( .IN1(n2484), .IN2(n1533), .IN3(n2485), .IN4(n1638), .IN5(
        n2533), .Q(n2221) );
  AO22X1 U2051 ( .IN1(n2487), .IN2(n1646), .IN3(n2488), .IN4(n1425), .Q(n2533)
         );
  AND2X1 U2052 ( .IN1(n2352), .IN2(n1392), .Q(n2473) );
  AO221X1 U2053 ( .IN1(n2354), .IN2(n2389), .IN3(n2352), .IN4(n2388), .IN5(
        n2534), .Q(n2340) );
  AO22X1 U2054 ( .IN1(n2359), .IN2(n2387), .IN3(n2356), .IN4(n2391), .Q(n2534)
         );
  AO221X1 U2055 ( .IN1(n2484), .IN2(n1426), .IN3(n2485), .IN4(n1384), .IN5(
        n2535), .Q(n2391) );
  AO22X1 U2056 ( .IN1(n2487), .IN2(n1570), .IN3(n2488), .IN4(n1370), .Q(n2535)
         );
  AO221X1 U2057 ( .IN1(n2484), .IN2(n1428), .IN3(n2485), .IN4(n1569), .IN5(
        n2536), .Q(n2387) );
  AO22X1 U2058 ( .IN1(n2487), .IN2(n1568), .IN3(n2488), .IN4(n1427), .Q(n2536)
         );
  AO221X1 U2059 ( .IN1(n2484), .IN2(n1572), .IN3(n2485), .IN4(n1429), .IN5(
        n2537), .Q(n2388) );
  AO22X1 U2060 ( .IN1(n2487), .IN2(n1432), .IN3(n2488), .IN4(n1571), .Q(n2537)
         );
  AO221X1 U2061 ( .IN1(n2484), .IN2(n1574), .IN3(n2485), .IN4(n1431), .IN5(
        n2538), .Q(n2389) );
  AO22X1 U2062 ( .IN1(n2487), .IN2(n1385), .IN3(n2488), .IN4(n1573), .Q(n2538)
         );
  AO222X1 U2063 ( .IN1(n2310), .IN2(n2314), .IN3(n2539), .IN4(n2478), .IN5(
        n2290), .IN6(n1578), .Q(\fpu_div_frac_dp/n1223 ) );
  AND2X1 U2064 ( .IN1(n1886), .IN2(\fpu_div_frac_dp/n978 ), .Q(n2478) );
  INVX0 U2065 ( .INP(n2288), .ZN(n2539) );
  AO21X1 U2066 ( .IN1(n2342), .IN2(n2540), .IN3(n2541), .Q(n2288) );
  MUX21X1 U2067 ( .IN1(n2542), .IN2(n2346), .S(n1392), .Q(n2541) );
  AO221X1 U2068 ( .IN1(n2354), .IN2(n2436), .IN3(n2352), .IN4(n2475), .IN5(
        n2543), .Q(n2346) );
  AO22X1 U2069 ( .IN1(n2359), .IN2(n2403), .IN3(n2356), .IN4(n2411), .Q(n2543)
         );
  AO221X1 U2070 ( .IN1(n2484), .IN2(n1411), .IN3(n2485), .IN4(n1553), .IN5(
        n2544), .Q(n2411) );
  AO22X1 U2071 ( .IN1(n2487), .IN2(n1554), .IN3(n2488), .IN4(n1412), .Q(n2544)
         );
  AO221X1 U2072 ( .IN1(n2484), .IN2(n1413), .IN3(n2485), .IN4(n1555), .IN5(
        n2545), .Q(n2403) );
  AO22X1 U2073 ( .IN1(n2487), .IN2(n1556), .IN3(n2488), .IN4(n1414), .Q(n2545)
         );
  AO221X1 U2074 ( .IN1(n2484), .IN2(n1415), .IN3(n2485), .IN4(n1557), .IN5(
        n2546), .Q(n2475) );
  AO22X1 U2075 ( .IN1(n2487), .IN2(n1558), .IN3(n2488), .IN4(n1416), .Q(n2546)
         );
  AO221X1 U2076 ( .IN1(n2484), .IN2(n1417), .IN3(n2485), .IN4(n1559), .IN5(
        n2547), .Q(n2436) );
  AO22X1 U2077 ( .IN1(n2487), .IN2(n1560), .IN3(n2488), .IN4(n1418), .Q(n2547)
         );
  AO222X1 U2078 ( .IN1(n2354), .IN2(n2470), .IN3(n2356), .IN4(n2477), .IN5(
        n2359), .IN6(n2476), .Q(n2542) );
  AO221X1 U2079 ( .IN1(n2484), .IN2(n1419), .IN3(n2485), .IN4(n1561), .IN5(
        n2548), .Q(n2476) );
  AO22X1 U2080 ( .IN1(n2487), .IN2(n1562), .IN3(n2488), .IN4(n1420), .Q(n2548)
         );
  AO221X1 U2081 ( .IN1(n2484), .IN2(n1421), .IN3(n2485), .IN4(n1563), .IN5(
        n2549), .Q(n2477) );
  AO22X1 U2082 ( .IN1(n2487), .IN2(n1564), .IN3(n2488), .IN4(n1422), .Q(n2549)
         );
  AO221X1 U2083 ( .IN1(n2484), .IN2(n1423), .IN3(n2485), .IN4(n1565), .IN5(
        n2550), .Q(n2470) );
  AO22X1 U2084 ( .IN1(n2487), .IN2(n1566), .IN3(n2488), .IN4(n1424), .Q(n2550)
         );
  AO221X1 U2085 ( .IN1(n2484), .IN2(n1530), .IN3(n2485), .IN4(n1721), .IN5(
        n2551), .Q(n2540) );
  AO22X1 U2086 ( .IN1(n2487), .IN2(n1567), .IN3(n2488), .IN4(
        \fpu_div_frac_dp/div_shl_data[52] ), .Q(n2551) );
  AND2X1 U2087 ( .IN1(n2352), .IN2(\fpu_div_frac_dp/n967 ), .Q(n2342) );
  INVX0 U2088 ( .INP(n2243), .ZN(n2314) );
  MUX21X1 U2089 ( .IN1(n2344), .IN2(n2225), .S(n1392), .Q(n2243) );
  INVX0 U2090 ( .INP(n2296), .ZN(n2225) );
  NAND2X0 U2091 ( .IN1(n2552), .IN2(\fpu_div_frac_dp/n980 ), .QN(n2296) );
  MUX21X1 U2092 ( .IN1(n2401), .IN2(n2218), .S(n1394), .Q(n2552) );
  INVX0 U2093 ( .INP(n2289), .ZN(n2218) );
  NAND2X0 U2094 ( .IN1(n2488), .IN2(n1646), .QN(n2289) );
  AO221X1 U2095 ( .IN1(n2484), .IN2(n1638), .IN3(n2485), .IN4(n1425), .IN5(
        n2553), .Q(n2401) );
  AO22X1 U2096 ( .IN1(n2487), .IN2(n1533), .IN3(n2488), .IN4(n1568), .Q(n2553)
         );
  AO221X1 U2097 ( .IN1(n2354), .IN2(n2404), .IN3(n2352), .IN4(n2407), .IN5(
        n2554), .Q(n2344) );
  AO22X1 U2098 ( .IN1(n2359), .IN2(n2402), .IN3(n2356), .IN4(n2406), .Q(n2554)
         );
  AO221X1 U2099 ( .IN1(n2484), .IN2(n1384), .IN3(n2485), .IN4(n1370), .IN5(
        n2555), .Q(n2406) );
  AO22X1 U2100 ( .IN1(n2487), .IN2(n1426), .IN3(n2488), .IN4(n1385), .Q(n2555)
         );
  NOR2X0 U2101 ( .IN1(n1394), .IN2(\fpu_div_frac_dp/n980 ), .QN(n2356) );
  AO221X1 U2102 ( .IN1(n2484), .IN2(n1569), .IN3(n2485), .IN4(n1427), .IN5(
        n2556), .Q(n2402) );
  AO22X1 U2103 ( .IN1(n2487), .IN2(n1428), .IN3(n2488), .IN4(n1570), .Q(n2556)
         );
  NOR2X0 U2104 ( .IN1(\fpu_div_frac_dp/n968 ), .IN2(\fpu_div_frac_dp/n980 ), 
        .QN(n2359) );
  AO221X1 U2105 ( .IN1(n2484), .IN2(n1429), .IN3(n2485), .IN4(n1571), .IN5(
        n2557), .Q(n2407) );
  AO22X1 U2106 ( .IN1(n2487), .IN2(n1572), .IN3(n2488), .IN4(n1430), .Q(n2557)
         );
  NOR2X0 U2107 ( .IN1(n1546), .IN2(n1394), .QN(n2352) );
  AO221X1 U2108 ( .IN1(n2484), .IN2(n1431), .IN3(n2485), .IN4(n1573), .IN5(
        n2558), .Q(n2404) );
  AO22X1 U2109 ( .IN1(n2487), .IN2(n1574), .IN3(n2488), .IN4(n1432), .Q(n2558)
         );
  NOR2X0 U2110 ( .IN1(n1544), .IN2(n1398), .QN(n2488) );
  NOR2X0 U2111 ( .IN1(\fpu_div_frac_dp/n960 ), .IN2(\fpu_div_frac_dp/n994 ), 
        .QN(n2487) );
  NOR2X0 U2112 ( .IN1(n1544), .IN2(\fpu_div_frac_dp/n960 ), .QN(n2485) );
  NOR2X0 U2113 ( .IN1(n1398), .IN2(\fpu_div_frac_dp/n994 ), .QN(n2484) );
  NOR2X0 U2114 ( .IN1(n1546), .IN2(\fpu_div_frac_dp/n968 ), .QN(n2354) );
  AND2X1 U2115 ( .IN1(n1884), .IN2(n1540), .Q(n2310) );
  AO21X1 U2116 ( .IN1(n2290), .IN2(n1635), .IN3(n1883), .Q(
        \fpu_div_frac_dp/n1222 ) );
  AO21X1 U2117 ( .IN1(n2290), .IN2(n1866), .IN3(n1886), .Q(
        \fpu_div_frac_dp/n1221 ) );
  AND2X1 U2118 ( .IN1(n2559), .IN2(n1047), .Q(n2290) );
  AO221X1 U2119 ( .IN1(n2560), .IN2(n1529), .IN3(n2561), .IN4(n1637), .IN5(
        n2562), .Q(\fpu_div_frac_dp/n1220 ) );
  AO221X1 U2120 ( .IN1(n2563), .IN2(n2564), .IN3(n2565), .IN4(n1383), .IN5(
        n2566), .Q(n2562) );
  AO221X1 U2121 ( .IN1(n2560), .IN2(div_frac_outa[0]), .IN3(n2561), .IN4(n1362), .IN5(n2567), .Q(\fpu_div_frac_dp/n1219 ) );
  AO221X1 U2122 ( .IN1(n2568), .IN2(n2563), .IN3(n2569), .IN4(n2570), .IN5(
        n2566), .Q(n2567) );
  AO221X1 U2123 ( .IN1(n2560), .IN2(div_frac_outa[1]), .IN3(n2561), .IN4(n1512), .IN5(n2571), .Q(\fpu_div_frac_dp/n1218 ) );
  AO221X1 U2124 ( .IN1(n2572), .IN2(n2563), .IN3(n2569), .IN4(div_frac_outa[0]), .IN5(n2566), .Q(n2571) );
  AO221X1 U2125 ( .IN1(n2560), .IN2(div_frac_outa[2]), .IN3(n2561), .IN4(n1493), .IN5(n2573), .Q(\fpu_div_frac_dp/n1217 ) );
  AO221X1 U2126 ( .IN1(n2574), .IN2(n2563), .IN3(n2569), .IN4(div_frac_outa[1]), .IN5(n2566), .Q(n2573) );
  AO221X1 U2127 ( .IN1(n2560), .IN2(div_frac_outa[3]), .IN3(n2561), .IN4(n1513), .IN5(n2575), .Q(\fpu_div_frac_dp/n1216 ) );
  AO221X1 U2128 ( .IN1(n2576), .IN2(n2563), .IN3(n2569), .IN4(div_frac_outa[2]), .IN5(n2566), .Q(n2575) );
  AO221X1 U2129 ( .IN1(n2560), .IN2(div_frac_outa[4]), .IN3(n2561), .IN4(n1516), .IN5(n2577), .Q(\fpu_div_frac_dp/n1215 ) );
  AO221X1 U2130 ( .IN1(n2578), .IN2(n2563), .IN3(n2569), .IN4(div_frac_outa[3]), .IN5(n2566), .Q(n2577) );
  AO221X1 U2131 ( .IN1(n2560), .IN2(div_frac_outa[5]), .IN3(n2561), .IN4(n1404), .IN5(n2579), .Q(\fpu_div_frac_dp/n1214 ) );
  AO221X1 U2132 ( .IN1(n2580), .IN2(n2563), .IN3(n2569), .IN4(div_frac_outa[4]), .IN5(n2566), .Q(n2579) );
  AO221X1 U2133 ( .IN1(n2560), .IN2(div_frac_outa[6]), .IN3(n2561), .IN4(n1379), .IN5(n2581), .Q(\fpu_div_frac_dp/n1213 ) );
  AO221X1 U2134 ( .IN1(n2582), .IN2(n2563), .IN3(n2569), .IN4(div_frac_outa[5]), .IN5(n2566), .Q(n2581) );
  AO221X1 U2135 ( .IN1(n2560), .IN2(div_frac_outa[7]), .IN3(n2561), .IN4(n1365), .IN5(n2583), .Q(\fpu_div_frac_dp/n1212 ) );
  AO221X1 U2136 ( .IN1(n2584), .IN2(n2563), .IN3(n2569), .IN4(div_frac_outa[6]), .IN5(n2566), .Q(n2583) );
  AO221X1 U2137 ( .IN1(n2560), .IN2(div_frac_outa[8]), .IN3(n2561), .IN4(n1359), .IN5(n2585), .Q(\fpu_div_frac_dp/n1211 ) );
  AO221X1 U2138 ( .IN1(n2586), .IN2(n2563), .IN3(n2569), .IN4(div_frac_outa[7]), .IN5(n2566), .Q(n2585) );
  AO221X1 U2139 ( .IN1(n2560), .IN2(div_frac_outa[9]), .IN3(n2561), .IN4(n1366), .IN5(n2587), .Q(\fpu_div_frac_dp/n1210 ) );
  AO221X1 U2140 ( .IN1(n2588), .IN2(n2563), .IN3(n2569), .IN4(div_frac_outa[8]), .IN5(n2566), .Q(n2587) );
  AO221X1 U2141 ( .IN1(n2560), .IN2(div_frac_outa[10]), .IN3(n2561), .IN4(
        n1380), .IN5(n2589), .Q(\fpu_div_frac_dp/n1209 ) );
  AO221X1 U2142 ( .IN1(n2590), .IN2(n2563), .IN3(n2569), .IN4(div_frac_outa[9]), .IN5(n2566), .Q(n2589) );
  AO221X1 U2143 ( .IN1(n2560), .IN2(div_frac_outa[11]), .IN3(n2561), .IN4(
        n1517), .IN5(n2591), .Q(\fpu_div_frac_dp/n1208 ) );
  AO221X1 U2144 ( .IN1(n2592), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[10]), .IN5(n2566), .Q(n2591) );
  AO221X1 U2145 ( .IN1(n2560), .IN2(div_frac_outa[12]), .IN3(n2561), .IN4(
        n1500), .IN5(n2593), .Q(\fpu_div_frac_dp/n1207 ) );
  AO221X1 U2146 ( .IN1(n2594), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[11]), .IN5(n2566), .Q(n2593) );
  AO221X1 U2147 ( .IN1(n2560), .IN2(div_frac_outa[13]), .IN3(n2561), .IN4(
        n1358), .IN5(n2595), .Q(\fpu_div_frac_dp/n1206 ) );
  AO221X1 U2148 ( .IN1(n2596), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[12]), .IN5(n2566), .Q(n2595) );
  AO221X1 U2149 ( .IN1(n2560), .IN2(div_frac_outa[14]), .IN3(n2561), .IN4(
        n1363), .IN5(n2597), .Q(\fpu_div_frac_dp/n1205 ) );
  AO221X1 U2150 ( .IN1(n2598), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[13]), .IN5(n2566), .Q(n2597) );
  AO221X1 U2151 ( .IN1(n2560), .IN2(div_frac_outa[15]), .IN3(n2561), .IN4(
        n1405), .IN5(n2599), .Q(\fpu_div_frac_dp/n1204 ) );
  AO221X1 U2152 ( .IN1(n2600), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[14]), .IN5(n2566), .Q(n2599) );
  AO221X1 U2153 ( .IN1(n2560), .IN2(div_frac_outa[16]), .IN3(n2561), .IN4(
        n1381), .IN5(n2601), .Q(\fpu_div_frac_dp/n1203 ) );
  AO221X1 U2154 ( .IN1(n2602), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[15]), .IN5(n2566), .Q(n2601) );
  AO221X1 U2155 ( .IN1(n2560), .IN2(div_frac_outa[17]), .IN3(n2561), .IN4(
        n1501), .IN5(n2603), .Q(\fpu_div_frac_dp/n1202 ) );
  AO221X1 U2156 ( .IN1(n2604), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[16]), .IN5(n2566), .Q(n2603) );
  AO221X1 U2157 ( .IN1(n2560), .IN2(div_frac_outa[18]), .IN3(n2561), .IN4(
        n1518), .IN5(n2605), .Q(\fpu_div_frac_dp/n1201 ) );
  AO221X1 U2158 ( .IN1(n2606), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[17]), .IN5(n2566), .Q(n2605) );
  AO221X1 U2159 ( .IN1(n2560), .IN2(div_frac_outa[19]), .IN3(n2561), .IN4(
        n1502), .IN5(n2607), .Q(\fpu_div_frac_dp/n1200 ) );
  AO221X1 U2160 ( .IN1(n2608), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[18]), .IN5(n2566), .Q(n2607) );
  AO221X1 U2161 ( .IN1(n2560), .IN2(div_frac_outa[20]), .IN3(n2561), .IN4(
        n1357), .IN5(n2609), .Q(\fpu_div_frac_dp/n1199 ) );
  AO221X1 U2162 ( .IN1(n2610), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[19]), .IN5(n2566), .Q(n2609) );
  AO221X1 U2163 ( .IN1(n2560), .IN2(div_frac_outa[21]), .IN3(n2561), .IN4(
        n1406), .IN5(n2611), .Q(\fpu_div_frac_dp/n1198 ) );
  AO221X1 U2164 ( .IN1(n2612), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[20]), .IN5(n2566), .Q(n2611) );
  AO221X1 U2165 ( .IN1(n2560), .IN2(div_frac_outa[22]), .IN3(n2561), .IN4(
        n1382), .IN5(n2613), .Q(\fpu_div_frac_dp/n1197 ) );
  AO221X1 U2166 ( .IN1(n2614), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[21]), .IN5(n2566), .Q(n2613) );
  AO221X1 U2167 ( .IN1(n2560), .IN2(div_frac_outa[23]), .IN3(n2561), .IN4(
        n1503), .IN5(n2615), .Q(\fpu_div_frac_dp/n1196 ) );
  AO221X1 U2168 ( .IN1(n2616), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[22]), .IN5(n2566), .Q(n2615) );
  AO221X1 U2169 ( .IN1(n2560), .IN2(div_frac_outa[24]), .IN3(n2561), .IN4(
        n1519), .IN5(n2617), .Q(\fpu_div_frac_dp/n1195 ) );
  AO221X1 U2170 ( .IN1(n2618), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[23]), .IN5(n2566), .Q(n2617) );
  AO221X1 U2171 ( .IN1(n2560), .IN2(div_frac_outa[25]), .IN3(n2561), .IN4(
        n1504), .IN5(n2619), .Q(\fpu_div_frac_dp/n1194 ) );
  AO221X1 U2172 ( .IN1(n2620), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[24]), .IN5(n2566), .Q(n2619) );
  AO221X1 U2173 ( .IN1(n2560), .IN2(div_frac_outa[26]), .IN3(n2561), .IN4(
        n1377), .IN5(n2621), .Q(\fpu_div_frac_dp/n1193 ) );
  AO221X1 U2174 ( .IN1(n2622), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[25]), .IN5(n2566), .Q(n2621) );
  AO221X1 U2175 ( .IN1(n2560), .IN2(div_frac_outa[27]), .IN3(n2561), .IN4(
        n1402), .IN5(n2623), .Q(\fpu_div_frac_dp/n1192 ) );
  AO221X1 U2176 ( .IN1(n2624), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[26]), .IN5(n2566), .Q(n2623) );
  AO221X1 U2177 ( .IN1(n2560), .IN2(div_frac_outa[28]), .IN3(n2561), .IN4(
        n1361), .IN5(n2625), .Q(\fpu_div_frac_dp/n1191 ) );
  AO221X1 U2178 ( .IN1(n2626), .IN2(n2563), .IN3(n2569), .IN4(
        div_frac_outa[27]), .IN5(n2566), .Q(n2625) );
  NAND4X0 U2179 ( .IN1(n2627), .IN2(n2628), .IN3(n2629), .IN4(n2630), .QN(
        \fpu_div_frac_dp/n1190 ) );
  OA222X1 U2180 ( .IN1(\fpu_div_frac_dp/n93 ), .IN2(n2631), .IN3(
        \fpu_div_frac_dp/n993 ), .IN4(n2632), .IN5(\fpu_div_frac_dp/n92 ), 
        .IN6(n2633), .Q(n2630) );
  NAND2X0 U2181 ( .IN1(n2634), .IN2(n2563), .QN(n2629) );
  NAND3X0 U2182 ( .IN1(n2635), .IN2(n1396), .IN3(n2570), .QN(n2627) );
  AO221X1 U2183 ( .IN1(n2560), .IN2(div_frac_outa[30]), .IN3(n2561), .IN4(
        n1520), .IN5(n2636), .Q(\fpu_div_frac_dp/n1189 ) );
  AO221X1 U2184 ( .IN1(n2637), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[29]), .IN5(n2566), .Q(n2636) );
  AO221X1 U2185 ( .IN1(n2560), .IN2(div_frac_outa[31]), .IN3(n2561), .IN4(
        n1505), .IN5(n2638), .Q(\fpu_div_frac_dp/n1188 ) );
  AO221X1 U2186 ( .IN1(n2639), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[30]), .IN5(n2566), .Q(n2638) );
  AO221X1 U2187 ( .IN1(n2560), .IN2(div_frac_outa[32]), .IN3(n2561), .IN4(
        n1506), .IN5(n2640), .Q(\fpu_div_frac_dp/n1187 ) );
  AO221X1 U2188 ( .IN1(n2641), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[31]), .IN5(n2566), .Q(n2640) );
  AO221X1 U2189 ( .IN1(n2560), .IN2(div_frac_outa[33]), .IN3(n2561), .IN4(
        n1507), .IN5(n2642), .Q(\fpu_div_frac_dp/n1186 ) );
  AO221X1 U2190 ( .IN1(n2643), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[32]), .IN5(n2566), .Q(n2642) );
  AO221X1 U2191 ( .IN1(n2560), .IN2(div_frac_outa[34]), .IN3(n2561), .IN4(
        n1521), .IN5(n2644), .Q(\fpu_div_frac_dp/n1185 ) );
  AO221X1 U2192 ( .IN1(n2645), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[33]), .IN5(n2566), .Q(n2644) );
  AO221X1 U2193 ( .IN1(n2560), .IN2(div_frac_outa[35]), .IN3(n2561), .IN4(
        n1494), .IN5(n2646), .Q(\fpu_div_frac_dp/n1184 ) );
  AO221X1 U2194 ( .IN1(n2647), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[34]), .IN5(n2566), .Q(n2646) );
  AO221X1 U2195 ( .IN1(n2560), .IN2(div_frac_outa[36]), .IN3(n2561), .IN4(
        n1497), .IN5(n2648), .Q(\fpu_div_frac_dp/n1183 ) );
  AO221X1 U2196 ( .IN1(n2649), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[35]), .IN5(n2566), .Q(n2648) );
  AO221X1 U2197 ( .IN1(n2560), .IN2(div_frac_outa[37]), .IN3(n2561), .IN4(
        n1495), .IN5(n2650), .Q(\fpu_div_frac_dp/n1182 ) );
  AO221X1 U2198 ( .IN1(n2651), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[36]), .IN5(n2566), .Q(n2650) );
  AO221X1 U2199 ( .IN1(n2560), .IN2(div_frac_outa[38]), .IN3(n2561), .IN4(
        n1514), .IN5(n2652), .Q(\fpu_div_frac_dp/n1181 ) );
  AO221X1 U2200 ( .IN1(n2653), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[37]), .IN5(n2566), .Q(n2652) );
  AO221X1 U2201 ( .IN1(n2560), .IN2(div_frac_outa[39]), .IN3(n2561), .IN4(
        n1508), .IN5(n2654), .Q(\fpu_div_frac_dp/n1180 ) );
  AO221X1 U2202 ( .IN1(n2655), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[38]), .IN5(n2566), .Q(n2654) );
  AO221X1 U2203 ( .IN1(n2560), .IN2(div_frac_outa[40]), .IN3(n2561), .IN4(
        n1509), .IN5(n2656), .Q(\fpu_div_frac_dp/n1179 ) );
  AO221X1 U2204 ( .IN1(n2657), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[39]), .IN5(n2566), .Q(n2656) );
  AO221X1 U2205 ( .IN1(n2560), .IN2(div_frac_outa[41]), .IN3(n2561), .IN4(
        n1522), .IN5(n2658), .Q(\fpu_div_frac_dp/n1178 ) );
  AO221X1 U2206 ( .IN1(n2659), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[40]), .IN5(n2566), .Q(n2658) );
  AO221X1 U2207 ( .IN1(n2560), .IN2(div_frac_outa[42]), .IN3(n2561), .IN4(
        n1498), .IN5(n2660), .Q(\fpu_div_frac_dp/n1177 ) );
  AO221X1 U2208 ( .IN1(n2661), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[41]), .IN5(n2566), .Q(n2660) );
  AO221X1 U2209 ( .IN1(n2560), .IN2(div_frac_outa[43]), .IN3(n2561), .IN4(
        n1496), .IN5(n2662), .Q(\fpu_div_frac_dp/n1176 ) );
  AO221X1 U2210 ( .IN1(n2663), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[42]), .IN5(n2566), .Q(n2662) );
  AO221X1 U2211 ( .IN1(n2560), .IN2(div_frac_outa[44]), .IN3(n2561), .IN4(
        n1515), .IN5(n2664), .Q(\fpu_div_frac_dp/n1175 ) );
  AO221X1 U2212 ( .IN1(n2665), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[43]), .IN5(n2566), .Q(n2664) );
  AO221X1 U2213 ( .IN1(n2560), .IN2(div_frac_outa[45]), .IN3(n2561), .IN4(
        n1510), .IN5(n2666), .Q(\fpu_div_frac_dp/n1174 ) );
  AO221X1 U2214 ( .IN1(n2667), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[44]), .IN5(n2566), .Q(n2666) );
  AO221X1 U2215 ( .IN1(n2560), .IN2(div_frac_outa[46]), .IN3(n2561), .IN4(
        n1511), .IN5(n2668), .Q(\fpu_div_frac_dp/n1173 ) );
  AO221X1 U2216 ( .IN1(n2669), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[45]), .IN5(n2566), .Q(n2668) );
  AO221X1 U2217 ( .IN1(n2560), .IN2(div_frac_outa[47]), .IN3(n2561), .IN4(
        n1523), .IN5(n2670), .Q(\fpu_div_frac_dp/n1172 ) );
  AO221X1 U2218 ( .IN1(n2671), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[46]), .IN5(n2566), .Q(n2670) );
  AO221X1 U2219 ( .IN1(n2560), .IN2(div_frac_outa[48]), .IN3(n2561), .IN4(
        n1378), .IN5(n2672), .Q(\fpu_div_frac_dp/n1171 ) );
  AO221X1 U2220 ( .IN1(n2673), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[47]), .IN5(n2566), .Q(n2672) );
  AO221X1 U2221 ( .IN1(n2560), .IN2(div_frac_outa[49]), .IN3(n2561), .IN4(
        n1407), .IN5(n2674), .Q(\fpu_div_frac_dp/n1170 ) );
  AO221X1 U2222 ( .IN1(n2675), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[48]), .IN5(n2566), .Q(n2674) );
  AO221X1 U2223 ( .IN1(n2560), .IN2(div_frac_outa[50]), .IN3(n2561), .IN4(
        n1364), .IN5(n2676), .Q(\fpu_div_frac_dp/n1169 ) );
  AO221X1 U2224 ( .IN1(n2677), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[49]), .IN5(n2566), .Q(n2676) );
  AO221X1 U2225 ( .IN1(n2560), .IN2(div_frac_outa[51]), .IN3(n2561), .IN4(
        n1526), .IN5(n2678), .Q(\fpu_div_frac_dp/n1168 ) );
  AO221X1 U2226 ( .IN1(n2679), .IN2(n2563), .IN3(n2565), .IN4(
        div_frac_outa[50]), .IN5(n2566), .Q(n2678) );
  AO221X1 U2227 ( .IN1(n2560), .IN2(n1383), .IN3(n2561), .IN4(n1636), .IN5(
        n2680), .Q(\fpu_div_frac_dp/n1167 ) );
  AO221X1 U2228 ( .IN1(n2563), .IN2(n2204), .IN3(n2565), .IN4(
        div_frac_outa[51]), .IN5(n2566), .Q(n2680) );
  AO21X1 U2229 ( .IN1(n2681), .IN2(n1362), .IN3(n2682), .Q(
        \fpu_div_frac_dp/n1166 ) );
  AO21X1 U2230 ( .IN1(n2681), .IN2(n1512), .IN3(n2683), .Q(
        \fpu_div_frac_dp/n1165 ) );
  AO21X1 U2231 ( .IN1(n2681), .IN2(n1493), .IN3(n2684), .Q(
        \fpu_div_frac_dp/n1164 ) );
  AO21X1 U2232 ( .IN1(n2681), .IN2(n1513), .IN3(n2685), .Q(
        \fpu_div_frac_dp/n1163 ) );
  AO21X1 U2233 ( .IN1(n2681), .IN2(n1516), .IN3(n2686), .Q(
        \fpu_div_frac_dp/n1162 ) );
  AO21X1 U2234 ( .IN1(n2681), .IN2(n1404), .IN3(n2687), .Q(
        \fpu_div_frac_dp/n1161 ) );
  AO21X1 U2235 ( .IN1(n2681), .IN2(n1379), .IN3(n2688), .Q(
        \fpu_div_frac_dp/n1160 ) );
  AO21X1 U2236 ( .IN1(n2681), .IN2(n1365), .IN3(n2689), .Q(
        \fpu_div_frac_dp/n1159 ) );
  AO21X1 U2237 ( .IN1(n2681), .IN2(n1359), .IN3(n2690), .Q(
        \fpu_div_frac_dp/n1158 ) );
  AO21X1 U2238 ( .IN1(n2681), .IN2(n1366), .IN3(n2691), .Q(
        \fpu_div_frac_dp/n1157 ) );
  AO21X1 U2239 ( .IN1(n2681), .IN2(n1380), .IN3(n2692), .Q(
        \fpu_div_frac_dp/n1156 ) );
  AO21X1 U2240 ( .IN1(n2681), .IN2(n1517), .IN3(n2693), .Q(
        \fpu_div_frac_dp/n1155 ) );
  AO21X1 U2241 ( .IN1(n2681), .IN2(n1500), .IN3(n2694), .Q(
        \fpu_div_frac_dp/n1154 ) );
  AO21X1 U2242 ( .IN1(n2681), .IN2(n1358), .IN3(n2695), .Q(
        \fpu_div_frac_dp/n1153 ) );
  AO21X1 U2243 ( .IN1(n2681), .IN2(n1363), .IN3(n2696), .Q(
        \fpu_div_frac_dp/n1152 ) );
  AO21X1 U2244 ( .IN1(n2681), .IN2(n1405), .IN3(n2697), .Q(
        \fpu_div_frac_dp/n1151 ) );
  AO21X1 U2245 ( .IN1(n2681), .IN2(n1381), .IN3(n2698), .Q(
        \fpu_div_frac_dp/n1150 ) );
  AO21X1 U2246 ( .IN1(n2681), .IN2(n1501), .IN3(n2699), .Q(
        \fpu_div_frac_dp/n1149 ) );
  AO21X1 U2247 ( .IN1(n2681), .IN2(n1518), .IN3(n2700), .Q(
        \fpu_div_frac_dp/n1148 ) );
  AO21X1 U2248 ( .IN1(n2681), .IN2(n1502), .IN3(n2701), .Q(
        \fpu_div_frac_dp/n1147 ) );
  AO21X1 U2249 ( .IN1(n2681), .IN2(n1357), .IN3(n2702), .Q(
        \fpu_div_frac_dp/n1146 ) );
  AO21X1 U2250 ( .IN1(n2681), .IN2(n1406), .IN3(n2703), .Q(
        \fpu_div_frac_dp/n1145 ) );
  AO21X1 U2251 ( .IN1(n2681), .IN2(n1382), .IN3(n2704), .Q(
        \fpu_div_frac_dp/n1144 ) );
  AO21X1 U2252 ( .IN1(n2681), .IN2(n1503), .IN3(n2705), .Q(
        \fpu_div_frac_dp/n1143 ) );
  AO21X1 U2253 ( .IN1(n2681), .IN2(n1519), .IN3(n2706), .Q(
        \fpu_div_frac_dp/n1142 ) );
  AO21X1 U2254 ( .IN1(n2681), .IN2(n1504), .IN3(n2707), .Q(
        \fpu_div_frac_dp/n1141 ) );
  AO21X1 U2255 ( .IN1(n2681), .IN2(n1377), .IN3(n2708), .Q(
        \fpu_div_frac_dp/n1140 ) );
  AO21X1 U2256 ( .IN1(n2681), .IN2(n1402), .IN3(n2709), .Q(
        \fpu_div_frac_dp/n1139 ) );
  AO21X1 U2257 ( .IN1(n2681), .IN2(n1361), .IN3(n2710), .Q(
        \fpu_div_frac_dp/n1138 ) );
  AO21X1 U2258 ( .IN1(n2681), .IN2(n1537), .IN3(n2711), .Q(
        \fpu_div_frac_dp/n1137 ) );
  AO21X1 U2259 ( .IN1(n2681), .IN2(n1520), .IN3(n2712), .Q(
        \fpu_div_frac_dp/n1136 ) );
  AO21X1 U2260 ( .IN1(n2681), .IN2(n1505), .IN3(n2713), .Q(
        \fpu_div_frac_dp/n1135 ) );
  AO21X1 U2261 ( .IN1(n2681), .IN2(n1506), .IN3(n2714), .Q(
        \fpu_div_frac_dp/n1134 ) );
  AO21X1 U2262 ( .IN1(n2681), .IN2(n1507), .IN3(n2715), .Q(
        \fpu_div_frac_dp/n1133 ) );
  AO21X1 U2263 ( .IN1(n2681), .IN2(n1521), .IN3(n2716), .Q(
        \fpu_div_frac_dp/n1132 ) );
  AO21X1 U2264 ( .IN1(n2681), .IN2(n1494), .IN3(n2717), .Q(
        \fpu_div_frac_dp/n1131 ) );
  AO21X1 U2265 ( .IN1(n2681), .IN2(n1497), .IN3(n2718), .Q(
        \fpu_div_frac_dp/n1130 ) );
  AO21X1 U2266 ( .IN1(n2681), .IN2(n1495), .IN3(n2719), .Q(
        \fpu_div_frac_dp/n1129 ) );
  AO21X1 U2267 ( .IN1(n2681), .IN2(n1514), .IN3(n2720), .Q(
        \fpu_div_frac_dp/n1128 ) );
  AO21X1 U2268 ( .IN1(n2681), .IN2(n1508), .IN3(n2721), .Q(
        \fpu_div_frac_dp/n1127 ) );
  AO21X1 U2269 ( .IN1(n2681), .IN2(n1509), .IN3(n2722), .Q(
        \fpu_div_frac_dp/n1126 ) );
  AO21X1 U2270 ( .IN1(n2681), .IN2(n1522), .IN3(n2723), .Q(
        \fpu_div_frac_dp/n1125 ) );
  AO21X1 U2271 ( .IN1(n2681), .IN2(n1498), .IN3(n2724), .Q(
        \fpu_div_frac_dp/n1124 ) );
  AO21X1 U2272 ( .IN1(n2681), .IN2(n1496), .IN3(n2725), .Q(
        \fpu_div_frac_dp/n1123 ) );
  AO21X1 U2273 ( .IN1(n2681), .IN2(n1515), .IN3(n2726), .Q(
        \fpu_div_frac_dp/n1122 ) );
  AO21X1 U2274 ( .IN1(n2681), .IN2(n1510), .IN3(n2727), .Q(
        \fpu_div_frac_dp/n1121 ) );
  AO21X1 U2275 ( .IN1(n2681), .IN2(n1511), .IN3(n2728), .Q(
        \fpu_div_frac_dp/n1120 ) );
  AO21X1 U2276 ( .IN1(n2681), .IN2(n1523), .IN3(n2729), .Q(
        \fpu_div_frac_dp/n1119 ) );
  AO21X1 U2277 ( .IN1(n2681), .IN2(n1378), .IN3(n2730), .Q(
        \fpu_div_frac_dp/n1118 ) );
  AO21X1 U2278 ( .IN1(n2681), .IN2(n1407), .IN3(n2731), .Q(
        \fpu_div_frac_dp/n1117 ) );
  AO21X1 U2279 ( .IN1(n2681), .IN2(n1364), .IN3(n2732), .Q(
        \fpu_div_frac_dp/n1116 ) );
  AO21X1 U2280 ( .IN1(n2681), .IN2(n1526), .IN3(n2733), .Q(
        \fpu_div_frac_dp/n1115 ) );
  AO21X1 U2281 ( .IN1(n2681), .IN2(n1636), .IN3(n2734), .Q(
        \fpu_div_frac_dp/n1114 ) );
  AO21X1 U2282 ( .IN1(n2681), .IN2(n1637), .IN3(n2735), .Q(
        \fpu_div_frac_dp/n1113 ) );
  AO21X1 U2283 ( .IN1(n2681), .IN2(n1527), .IN3(n2682), .Q(
        \fpu_div_frac_dp/n1112 ) );
  AO222X1 U2284 ( .IN1(n2736), .IN2(div_frac_outa[1]), .IN3(n2737), .IN4(
        div_frac_outa[2]), .IN5(n1885), .IN6(n1729), .Q(n2682) );
  AO21X1 U2285 ( .IN1(n2681), .IN2(n1623), .IN3(n2683), .Q(
        \fpu_div_frac_dp/n1111 ) );
  AO221X1 U2286 ( .IN1(n1885), .IN2(n1733), .IN3(n2738), .IN4(n1362), .IN5(
        n2739), .Q(n2683) );
  AO222X1 U2287 ( .IN1(n2737), .IN2(div_frac_outa[3]), .IN3(n2740), .IN4(n2568), .IN5(n2736), .IN6(div_frac_outa[2]), .Q(n2739) );
  XNOR3X1 U2288 ( .IN1(n1373), .IN2(\fpu_div_frac_dp/n997 ), .IN3(n1527), .Q(
        n2568) );
  AO21X1 U2289 ( .IN1(n2681), .IN2(n1622), .IN3(n2684), .Q(
        \fpu_div_frac_dp/n1110 ) );
  AO221X1 U2290 ( .IN1(n1883), .IN2(n1734), .IN3(n2738), .IN4(n1512), .IN5(
        n2741), .Q(n2684) );
  AO222X1 U2291 ( .IN1(n2737), .IN2(div_frac_outa[4]), .IN3(n2740), .IN4(n2572), .IN5(n2736), .IN6(div_frac_outa[3]), .Q(n2741) );
  XNOR3X1 U2292 ( .IN1(n1437), .IN2(\fpu_div_frac_dp/n11 ), .IN3(n2742), .Q(
        n2572) );
  AO21X1 U2293 ( .IN1(n2681), .IN2(n1621), .IN3(n2685), .Q(
        \fpu_div_frac_dp/n1109 ) );
  AO221X1 U2294 ( .IN1(n1886), .IN2(n1735), .IN3(n2738), .IN4(n1493), .IN5(
        n2743), .Q(n2685) );
  AO222X1 U2295 ( .IN1(n2737), .IN2(div_frac_outa[5]), .IN3(n2740), .IN4(n2574), .IN5(n2736), .IN6(div_frac_outa[4]), .Q(n2743) );
  XNOR3X1 U2296 ( .IN1(n1436), .IN2(\fpu_div_frac_dp/n14 ), .IN3(n2744), .Q(
        n2574) );
  AO21X1 U2297 ( .IN1(n2681), .IN2(n1620), .IN3(n2686), .Q(
        \fpu_div_frac_dp/n1108 ) );
  AO221X1 U2298 ( .IN1(n1884), .IN2(n1736), .IN3(n2738), .IN4(n1513), .IN5(
        n2745), .Q(n2686) );
  AO222X1 U2299 ( .IN1(n2737), .IN2(div_frac_outa[6]), .IN3(n2740), .IN4(n2576), .IN5(n2736), .IN6(div_frac_outa[5]), .Q(n2745) );
  XNOR3X1 U2300 ( .IN1(n1435), .IN2(\fpu_div_frac_dp/n17 ), .IN3(n2746), .Q(
        n2576) );
  AO21X1 U2301 ( .IN1(n2681), .IN2(n1596), .IN3(n2687), .Q(
        \fpu_div_frac_dp/n1107 ) );
  AO221X1 U2302 ( .IN1(n1885), .IN2(n1737), .IN3(n2738), .IN4(n1516), .IN5(
        n2747), .Q(n2687) );
  AO222X1 U2303 ( .IN1(n2737), .IN2(div_frac_outa[7]), .IN3(n2740), .IN4(n2578), .IN5(n2736), .IN6(div_frac_outa[6]), .Q(n2747) );
  XNOR3X1 U2304 ( .IN1(n1434), .IN2(\fpu_div_frac_dp/n20 ), .IN3(n2748), .Q(
        n2578) );
  AO21X1 U2305 ( .IN1(n2681), .IN2(n1595), .IN3(n2688), .Q(
        \fpu_div_frac_dp/n1106 ) );
  AO221X1 U2306 ( .IN1(n1883), .IN2(n1738), .IN3(n2738), .IN4(n1404), .IN5(
        n2749), .Q(n2688) );
  AO222X1 U2307 ( .IN1(n2737), .IN2(div_frac_outa[8]), .IN3(n2740), .IN4(n2580), .IN5(n2736), .IN6(div_frac_outa[7]), .Q(n2749) );
  XNOR3X1 U2308 ( .IN1(n1596), .IN2(\fpu_div_frac_dp/n214 ), .IN3(n2750), .Q(
        n2580) );
  AO21X1 U2309 ( .IN1(n2681), .IN2(n1594), .IN3(n2689), .Q(
        \fpu_div_frac_dp/n1105 ) );
  AO221X1 U2310 ( .IN1(n1886), .IN2(n1739), .IN3(n2738), .IN4(n1379), .IN5(
        n2751), .Q(n2689) );
  AO222X1 U2311 ( .IN1(n2737), .IN2(div_frac_outa[9]), .IN3(n2740), .IN4(n2582), .IN5(n2736), .IN6(div_frac_outa[8]), .Q(n2751) );
  XNOR3X1 U2312 ( .IN1(n1595), .IN2(\fpu_div_frac_dp/n213 ), .IN3(n2752), .Q(
        n2582) );
  AO21X1 U2313 ( .IN1(n2681), .IN2(n1593), .IN3(n2690), .Q(
        \fpu_div_frac_dp/n1104 ) );
  AO221X1 U2314 ( .IN1(n1884), .IN2(n1740), .IN3(n2738), .IN4(n1365), .IN5(
        n2753), .Q(n2690) );
  AO222X1 U2315 ( .IN1(n2737), .IN2(div_frac_outa[10]), .IN3(n2740), .IN4(
        n2584), .IN5(n2736), .IN6(div_frac_outa[9]), .Q(n2753) );
  XNOR3X1 U2316 ( .IN1(n1594), .IN2(\fpu_div_frac_dp/n212 ), .IN3(n2754), .Q(
        n2584) );
  AO21X1 U2317 ( .IN1(n2681), .IN2(n1592), .IN3(n2691), .Q(
        \fpu_div_frac_dp/n1103 ) );
  AO221X1 U2318 ( .IN1(n1885), .IN2(n1741), .IN3(n2738), .IN4(n1359), .IN5(
        n2755), .Q(n2691) );
  AO222X1 U2319 ( .IN1(n2737), .IN2(div_frac_outa[11]), .IN3(n2740), .IN4(
        n2586), .IN5(n2736), .IN6(div_frac_outa[10]), .Q(n2755) );
  XNOR3X1 U2320 ( .IN1(n1593), .IN2(\fpu_div_frac_dp/n211 ), .IN3(n2756), .Q(
        n2586) );
  AO21X1 U2321 ( .IN1(n2681), .IN2(n1591), .IN3(n2692), .Q(
        \fpu_div_frac_dp/n1102 ) );
  AO221X1 U2322 ( .IN1(n1883), .IN2(n1742), .IN3(n2738), .IN4(n1366), .IN5(
        n2757), .Q(n2692) );
  AO222X1 U2323 ( .IN1(n2737), .IN2(div_frac_outa[12]), .IN3(n2740), .IN4(
        n2588), .IN5(n2736), .IN6(div_frac_outa[11]), .Q(n2757) );
  XNOR3X1 U2324 ( .IN1(n1592), .IN2(\fpu_div_frac_dp/n210 ), .IN3(n2758), .Q(
        n2588) );
  AO21X1 U2325 ( .IN1(n2681), .IN2(n1590), .IN3(n2693), .Q(
        \fpu_div_frac_dp/n1101 ) );
  AO221X1 U2326 ( .IN1(n1886), .IN2(n1743), .IN3(n2738), .IN4(n1380), .IN5(
        n2759), .Q(n2693) );
  AO222X1 U2327 ( .IN1(n2737), .IN2(div_frac_outa[13]), .IN3(n2740), .IN4(
        n2590), .IN5(n2736), .IN6(div_frac_outa[12]), .Q(n2759) );
  XNOR3X1 U2328 ( .IN1(n1591), .IN2(\fpu_div_frac_dp/n209 ), .IN3(n2760), .Q(
        n2590) );
  AO21X1 U2329 ( .IN1(n2681), .IN2(n1586), .IN3(n2694), .Q(
        \fpu_div_frac_dp/n1100 ) );
  AO221X1 U2330 ( .IN1(n1884), .IN2(n1744), .IN3(n2738), .IN4(n1517), .IN5(
        n2761), .Q(n2694) );
  AO222X1 U2331 ( .IN1(n2737), .IN2(div_frac_outa[14]), .IN3(n2740), .IN4(
        n2592), .IN5(n2736), .IN6(div_frac_outa[13]), .Q(n2761) );
  XNOR3X1 U2332 ( .IN1(n1590), .IN2(\fpu_div_frac_dp/n208 ), .IN3(n2762), .Q(
        n2592) );
  AO21X1 U2333 ( .IN1(n2681), .IN2(n1589), .IN3(n2695), .Q(
        \fpu_div_frac_dp/n1099 ) );
  AO221X1 U2334 ( .IN1(n1885), .IN2(n1745), .IN3(n2738), .IN4(n1500), .IN5(
        n2763), .Q(n2695) );
  AO222X1 U2335 ( .IN1(n2737), .IN2(div_frac_outa[15]), .IN3(n2740), .IN4(
        n2594), .IN5(n2736), .IN6(div_frac_outa[14]), .Q(n2763) );
  XNOR3X1 U2336 ( .IN1(n1586), .IN2(\fpu_div_frac_dp/n207 ), .IN3(n2764), .Q(
        n2594) );
  AO21X1 U2337 ( .IN1(n2681), .IN2(n1585), .IN3(n2696), .Q(
        \fpu_div_frac_dp/n1098 ) );
  AO221X1 U2338 ( .IN1(n1883), .IN2(n1746), .IN3(n2738), .IN4(n1358), .IN5(
        n2765), .Q(n2696) );
  AO222X1 U2339 ( .IN1(n2737), .IN2(div_frac_outa[16]), .IN3(n2740), .IN4(
        n2596), .IN5(n2736), .IN6(div_frac_outa[15]), .Q(n2765) );
  XNOR3X1 U2340 ( .IN1(n1589), .IN2(\fpu_div_frac_dp/n206 ), .IN3(n2766), .Q(
        n2596) );
  AO21X1 U2341 ( .IN1(n2681), .IN2(n1584), .IN3(n2697), .Q(
        \fpu_div_frac_dp/n1097 ) );
  AO221X1 U2342 ( .IN1(n1886), .IN2(n1747), .IN3(n2738), .IN4(n1363), .IN5(
        n2767), .Q(n2697) );
  AO222X1 U2343 ( .IN1(n2737), .IN2(div_frac_outa[17]), .IN3(n2740), .IN4(
        n2598), .IN5(n2736), .IN6(div_frac_outa[16]), .Q(n2767) );
  XNOR3X1 U2344 ( .IN1(n1585), .IN2(\fpu_div_frac_dp/n205 ), .IN3(n2768), .Q(
        n2598) );
  AO21X1 U2345 ( .IN1(n2681), .IN2(n1588), .IN3(n2698), .Q(
        \fpu_div_frac_dp/n1096 ) );
  AO221X1 U2346 ( .IN1(n1884), .IN2(n1748), .IN3(n2738), .IN4(n1405), .IN5(
        n2769), .Q(n2698) );
  AO222X1 U2347 ( .IN1(n2737), .IN2(div_frac_outa[18]), .IN3(n2740), .IN4(
        n2600), .IN5(n2736), .IN6(div_frac_outa[17]), .Q(n2769) );
  XNOR3X1 U2348 ( .IN1(n1584), .IN2(\fpu_div_frac_dp/n204 ), .IN3(n2770), .Q(
        n2600) );
  AO21X1 U2349 ( .IN1(n2681), .IN2(n1583), .IN3(n2699), .Q(
        \fpu_div_frac_dp/n1095 ) );
  AO221X1 U2350 ( .IN1(n1885), .IN2(n1749), .IN3(n2738), .IN4(n1381), .IN5(
        n2771), .Q(n2699) );
  AO222X1 U2351 ( .IN1(n2737), .IN2(div_frac_outa[19]), .IN3(n2740), .IN4(
        n2602), .IN5(n2736), .IN6(div_frac_outa[18]), .Q(n2771) );
  XNOR3X1 U2352 ( .IN1(n1588), .IN2(\fpu_div_frac_dp/n203 ), .IN3(n2772), .Q(
        n2602) );
  AO21X1 U2353 ( .IN1(n2681), .IN2(n1582), .IN3(n2700), .Q(
        \fpu_div_frac_dp/n1094 ) );
  AO221X1 U2354 ( .IN1(n1883), .IN2(n1750), .IN3(n2738), .IN4(n1501), .IN5(
        n2773), .Q(n2700) );
  AO222X1 U2355 ( .IN1(n2737), .IN2(div_frac_outa[20]), .IN3(n2740), .IN4(
        n2604), .IN5(n2736), .IN6(div_frac_outa[19]), .Q(n2773) );
  XNOR3X1 U2356 ( .IN1(n1583), .IN2(\fpu_div_frac_dp/n202 ), .IN3(n2774), .Q(
        n2604) );
  AO21X1 U2357 ( .IN1(n2681), .IN2(n1587), .IN3(n2701), .Q(
        \fpu_div_frac_dp/n1093 ) );
  AO221X1 U2358 ( .IN1(n1886), .IN2(n1751), .IN3(n2738), .IN4(n1518), .IN5(
        n2775), .Q(n2701) );
  AO222X1 U2359 ( .IN1(n2737), .IN2(div_frac_outa[21]), .IN3(n2740), .IN4(
        n2606), .IN5(n2736), .IN6(div_frac_outa[20]), .Q(n2775) );
  XNOR3X1 U2360 ( .IN1(n1582), .IN2(\fpu_div_frac_dp/n201 ), .IN3(n2776), .Q(
        n2606) );
  AO21X1 U2361 ( .IN1(n2681), .IN2(n1581), .IN3(n2702), .Q(
        \fpu_div_frac_dp/n1092 ) );
  AO221X1 U2362 ( .IN1(n1884), .IN2(n1752), .IN3(n2738), .IN4(n1502), .IN5(
        n2777), .Q(n2702) );
  AO222X1 U2363 ( .IN1(n2737), .IN2(div_frac_outa[22]), .IN3(n2740), .IN4(
        n2608), .IN5(n2736), .IN6(div_frac_outa[21]), .Q(n2777) );
  XNOR3X1 U2364 ( .IN1(n1587), .IN2(\fpu_div_frac_dp/n200 ), .IN3(n2778), .Q(
        n2608) );
  AO21X1 U2365 ( .IN1(n2681), .IN2(n1470), .IN3(n2703), .Q(
        \fpu_div_frac_dp/n1091 ) );
  AO221X1 U2366 ( .IN1(n1885), .IN2(n1753), .IN3(n2738), .IN4(n1357), .IN5(
        n2779), .Q(n2703) );
  AO222X1 U2367 ( .IN1(n2737), .IN2(div_frac_outa[23]), .IN3(n2740), .IN4(
        n2610), .IN5(n2736), .IN6(div_frac_outa[22]), .Q(n2779) );
  XNOR3X1 U2368 ( .IN1(n1581), .IN2(\fpu_div_frac_dp/n199 ), .IN3(n2780), .Q(
        n2610) );
  AO21X1 U2369 ( .IN1(n2681), .IN2(n1469), .IN3(n2704), .Q(
        \fpu_div_frac_dp/n1090 ) );
  AO221X1 U2370 ( .IN1(n1883), .IN2(n1754), .IN3(n2738), .IN4(n1406), .IN5(
        n2781), .Q(n2704) );
  AO222X1 U2371 ( .IN1(n2737), .IN2(div_frac_outa[24]), .IN3(n2740), .IN4(
        n2612), .IN5(n2736), .IN6(div_frac_outa[23]), .Q(n2781) );
  XNOR3X1 U2372 ( .IN1(n1470), .IN2(\fpu_div_frac_dp/n198 ), .IN3(n2782), .Q(
        n2612) );
  AO21X1 U2373 ( .IN1(n2681), .IN2(n1468), .IN3(n2705), .Q(
        \fpu_div_frac_dp/n1089 ) );
  AO221X1 U2374 ( .IN1(n1886), .IN2(n1755), .IN3(n2738), .IN4(n1382), .IN5(
        n2783), .Q(n2705) );
  AO222X1 U2375 ( .IN1(n2737), .IN2(div_frac_outa[25]), .IN3(n2740), .IN4(
        n2614), .IN5(n2736), .IN6(div_frac_outa[24]), .Q(n2783) );
  XNOR3X1 U2376 ( .IN1(n1469), .IN2(\fpu_div_frac_dp/n197 ), .IN3(n2784), .Q(
        n2614) );
  AO21X1 U2377 ( .IN1(n2681), .IN2(n1467), .IN3(n2706), .Q(
        \fpu_div_frac_dp/n1088 ) );
  AO221X1 U2378 ( .IN1(n1884), .IN2(n1756), .IN3(n2738), .IN4(n1503), .IN5(
        n2785), .Q(n2706) );
  AO222X1 U2379 ( .IN1(n2737), .IN2(div_frac_outa[26]), .IN3(n2740), .IN4(
        n2616), .IN5(n2736), .IN6(div_frac_outa[25]), .Q(n2785) );
  XNOR3X1 U2380 ( .IN1(n1468), .IN2(\fpu_div_frac_dp/n196 ), .IN3(n2786), .Q(
        n2616) );
  AO21X1 U2381 ( .IN1(n2681), .IN2(n1466), .IN3(n2707), .Q(
        \fpu_div_frac_dp/n1087 ) );
  AO221X1 U2382 ( .IN1(n1885), .IN2(n1757), .IN3(n2738), .IN4(n1519), .IN5(
        n2787), .Q(n2707) );
  AO222X1 U2383 ( .IN1(n2737), .IN2(div_frac_outa[27]), .IN3(n2740), .IN4(
        n2618), .IN5(n2736), .IN6(div_frac_outa[26]), .Q(n2787) );
  XNOR3X1 U2384 ( .IN1(n1467), .IN2(\fpu_div_frac_dp/n195 ), .IN3(n2788), .Q(
        n2618) );
  AO21X1 U2385 ( .IN1(n2681), .IN2(n1465), .IN3(n2708), .Q(
        \fpu_div_frac_dp/n1086 ) );
  AO221X1 U2386 ( .IN1(n1883), .IN2(n1758), .IN3(n2738), .IN4(n1504), .IN5(
        n2789), .Q(n2708) );
  AO222X1 U2387 ( .IN1(n2736), .IN2(div_frac_outa[27]), .IN3(n2737), .IN4(
        div_frac_outa[28]), .IN5(n2740), .IN6(n2620), .Q(n2789) );
  XNOR3X1 U2388 ( .IN1(n1466), .IN2(\fpu_div_frac_dp/n194 ), .IN3(n2790), .Q(
        n2620) );
  AO21X1 U2389 ( .IN1(n2681), .IN2(n1464), .IN3(n2709), .Q(
        \fpu_div_frac_dp/n1085 ) );
  AO221X1 U2390 ( .IN1(n1886), .IN2(n1759), .IN3(n2738), .IN4(n1377), .IN5(
        n2791), .Q(n2709) );
  AO222X1 U2391 ( .IN1(n2736), .IN2(div_frac_outa[28]), .IN3(n2737), .IN4(
        div_frac_outa[29]), .IN5(n2740), .IN6(n2622), .Q(n2791) );
  XNOR3X1 U2392 ( .IN1(n1465), .IN2(\fpu_div_frac_dp/n193 ), .IN3(n2792), .Q(
        n2622) );
  AO21X1 U2393 ( .IN1(n2681), .IN2(n1463), .IN3(n2710), .Q(
        \fpu_div_frac_dp/n1084 ) );
  AO221X1 U2394 ( .IN1(n1884), .IN2(n1760), .IN3(n2738), .IN4(n1402), .IN5(
        n2793), .Q(n2710) );
  AO222X1 U2395 ( .IN1(n2736), .IN2(div_frac_outa[29]), .IN3(n2737), .IN4(
        div_frac_outa[30]), .IN5(n2740), .IN6(n2624), .Q(n2793) );
  XNOR3X1 U2396 ( .IN1(n1464), .IN2(\fpu_div_frac_dp/n192 ), .IN3(n2794), .Q(
        n2624) );
  AND2X1 U2397 ( .IN1(n2795), .IN2(n2017), .Q(n2737) );
  AND2X1 U2398 ( .IN1(n2795), .IN2(n2796), .Q(n2736) );
  AND2X1 U2399 ( .IN1(n2010), .IN2(n1397), .Q(n2795) );
  AO21X1 U2400 ( .IN1(n2681), .IN2(n1612), .IN3(n2711), .Q(
        \fpu_div_frac_dp/n1083 ) );
  AO221X1 U2401 ( .IN1(n1885), .IN2(n1761), .IN3(n2738), .IN4(n1361), .IN5(
        n2797), .Q(n2711) );
  AO222X1 U2402 ( .IN1(n2798), .IN2(div_frac_outa[30]), .IN3(n2740), .IN4(
        n2626), .IN5(n2799), .IN6(div_frac_outa[31]), .Q(n2797) );
  XNOR3X1 U2403 ( .IN1(n1463), .IN2(\fpu_div_frac_dp/n191 ), .IN3(n2800), .Q(
        n2626) );
  AO21X1 U2404 ( .IN1(n2681), .IN2(n1462), .IN3(n2712), .Q(
        \fpu_div_frac_dp/n1082 ) );
  AO221X1 U2405 ( .IN1(n1883), .IN2(n1762), .IN3(n2738), .IN4(n1537), .IN5(
        n2801), .Q(n2712) );
  AO222X1 U2406 ( .IN1(n2798), .IN2(div_frac_outa[31]), .IN3(n2740), .IN4(
        n2634), .IN5(n2799), .IN6(div_frac_outa[32]), .Q(n2801) );
  XNOR3X1 U2407 ( .IN1(n1442), .IN2(\fpu_div_frac_dp/n94 ), .IN3(n2802), .Q(
        n2634) );
  AO21X1 U2408 ( .IN1(n2681), .IN2(n1619), .IN3(n2713), .Q(
        \fpu_div_frac_dp/n1081 ) );
  AO221X1 U2409 ( .IN1(n1886), .IN2(n1763), .IN3(n2738), .IN4(n1520), .IN5(
        n2803), .Q(n2713) );
  AO222X1 U2410 ( .IN1(n2798), .IN2(div_frac_outa[32]), .IN3(n2740), .IN4(
        n2637), .IN5(n2799), .IN6(div_frac_outa[33]), .Q(n2803) );
  XNOR3X1 U2411 ( .IN1(n1462), .IN2(\fpu_div_frac_dp/n189 ), .IN3(n2804), .Q(
        n2637) );
  AO21X1 U2412 ( .IN1(n2681), .IN2(n1611), .IN3(n2714), .Q(
        \fpu_div_frac_dp/n1080 ) );
  AO221X1 U2413 ( .IN1(n1884), .IN2(n1764), .IN3(n2738), .IN4(n1505), .IN5(
        n2805), .Q(n2714) );
  AO222X1 U2414 ( .IN1(n2798), .IN2(div_frac_outa[33]), .IN3(n2740), .IN4(
        n2639), .IN5(n2799), .IN6(div_frac_outa[34]), .Q(n2805) );
  XNOR3X1 U2415 ( .IN1(n1488), .IN2(\fpu_div_frac_dp/n100 ), .IN3(n2806), .Q(
        n2639) );
  AO21X1 U2416 ( .IN1(n2681), .IN2(n1610), .IN3(n2715), .Q(
        \fpu_div_frac_dp/n1079 ) );
  AO221X1 U2417 ( .IN1(n1885), .IN2(n1765), .IN3(n2738), .IN4(n1506), .IN5(
        n2807), .Q(n2715) );
  AO222X1 U2418 ( .IN1(n2798), .IN2(div_frac_outa[34]), .IN3(n2740), .IN4(
        n2641), .IN5(n2799), .IN6(div_frac_outa[35]), .Q(n2807) );
  XNOR3X1 U2419 ( .IN1(n1487), .IN2(\fpu_div_frac_dp/n103 ), .IN3(n2808), .Q(
        n2641) );
  AO21X1 U2420 ( .IN1(n2681), .IN2(n1618), .IN3(n2716), .Q(
        \fpu_div_frac_dp/n1078 ) );
  AO221X1 U2421 ( .IN1(n1883), .IN2(n1766), .IN3(n2738), .IN4(n1507), .IN5(
        n2809), .Q(n2716) );
  AO222X1 U2422 ( .IN1(n2798), .IN2(div_frac_outa[35]), .IN3(n2740), .IN4(
        n2643), .IN5(n2799), .IN6(div_frac_outa[36]), .Q(n2809) );
  XNOR3X1 U2423 ( .IN1(n1486), .IN2(\fpu_div_frac_dp/n106 ), .IN3(n2810), .Q(
        n2643) );
  AO21X1 U2424 ( .IN1(n2681), .IN2(n1609), .IN3(n2717), .Q(
        \fpu_div_frac_dp/n1077 ) );
  AO221X1 U2425 ( .IN1(n1886), .IN2(n1767), .IN3(n2738), .IN4(n1521), .IN5(
        n2811), .Q(n2717) );
  AO222X1 U2426 ( .IN1(n2798), .IN2(div_frac_outa[36]), .IN3(n2740), .IN4(
        n2645), .IN5(n2799), .IN6(div_frac_outa[37]), .Q(n2811) );
  XNOR3X1 U2427 ( .IN1(n1485), .IN2(\fpu_div_frac_dp/n109 ), .IN3(n2812), .Q(
        n2645) );
  AO21X1 U2428 ( .IN1(n2681), .IN2(n1608), .IN3(n2718), .Q(
        \fpu_div_frac_dp/n1076 ) );
  AO221X1 U2429 ( .IN1(n1884), .IN2(n1768), .IN3(n2738), .IN4(n1494), .IN5(
        n2813), .Q(n2718) );
  AO222X1 U2430 ( .IN1(n2798), .IN2(div_frac_outa[37]), .IN3(n2740), .IN4(
        n2647), .IN5(n2799), .IN6(div_frac_outa[38]), .Q(n2813) );
  XNOR3X1 U2431 ( .IN1(n1484), .IN2(\fpu_div_frac_dp/n112 ), .IN3(n2814), .Q(
        n2647) );
  AO21X1 U2432 ( .IN1(n2681), .IN2(n1617), .IN3(n2719), .Q(
        \fpu_div_frac_dp/n1075 ) );
  AO221X1 U2433 ( .IN1(n1885), .IN2(n1769), .IN3(n2738), .IN4(n1497), .IN5(
        n2815), .Q(n2719) );
  AO222X1 U2434 ( .IN1(n2798), .IN2(div_frac_outa[38]), .IN3(n2740), .IN4(
        n2649), .IN5(n2799), .IN6(div_frac_outa[39]), .Q(n2815) );
  XNOR3X1 U2435 ( .IN1(n1483), .IN2(\fpu_div_frac_dp/n115 ), .IN3(n2816), .Q(
        n2649) );
  AO21X1 U2436 ( .IN1(n2681), .IN2(n1607), .IN3(n2720), .Q(
        \fpu_div_frac_dp/n1074 ) );
  AO221X1 U2437 ( .IN1(n1883), .IN2(n1770), .IN3(n2738), .IN4(n1495), .IN5(
        n2817), .Q(n2720) );
  AO222X1 U2438 ( .IN1(n2798), .IN2(div_frac_outa[39]), .IN3(n2740), .IN4(
        n2651), .IN5(n2799), .IN6(div_frac_outa[40]), .Q(n2817) );
  XNOR3X1 U2439 ( .IN1(n1482), .IN2(\fpu_div_frac_dp/n118 ), .IN3(n2818), .Q(
        n2651) );
  AO21X1 U2440 ( .IN1(n2681), .IN2(n1606), .IN3(n2721), .Q(
        \fpu_div_frac_dp/n1073 ) );
  AO221X1 U2441 ( .IN1(n1886), .IN2(n1771), .IN3(n2738), .IN4(n1514), .IN5(
        n2819), .Q(n2721) );
  AO222X1 U2442 ( .IN1(n2798), .IN2(div_frac_outa[40]), .IN3(n2740), .IN4(
        n2653), .IN5(n2799), .IN6(div_frac_outa[41]), .Q(n2819) );
  XNOR3X1 U2443 ( .IN1(n1481), .IN2(\fpu_div_frac_dp/n121 ), .IN3(n2820), .Q(
        n2653) );
  AO21X1 U2444 ( .IN1(n2681), .IN2(n1616), .IN3(n2722), .Q(
        \fpu_div_frac_dp/n1072 ) );
  AO221X1 U2445 ( .IN1(n1884), .IN2(n1772), .IN3(n2738), .IN4(n1508), .IN5(
        n2821), .Q(n2722) );
  AO222X1 U2446 ( .IN1(n2798), .IN2(div_frac_outa[41]), .IN3(n2740), .IN4(
        n2655), .IN5(n2799), .IN6(div_frac_outa[42]), .Q(n2821) );
  XNOR3X1 U2447 ( .IN1(n1480), .IN2(\fpu_div_frac_dp/n124 ), .IN3(n2822), .Q(
        n2655) );
  AO21X1 U2448 ( .IN1(n2681), .IN2(n1605), .IN3(n2723), .Q(
        \fpu_div_frac_dp/n1071 ) );
  AO221X1 U2449 ( .IN1(n1885), .IN2(n1773), .IN3(n2738), .IN4(n1509), .IN5(
        n2823), .Q(n2723) );
  AO222X1 U2450 ( .IN1(n2798), .IN2(div_frac_outa[42]), .IN3(n2740), .IN4(
        n2657), .IN5(n2799), .IN6(div_frac_outa[43]), .Q(n2823) );
  XNOR3X1 U2451 ( .IN1(n1479), .IN2(\fpu_div_frac_dp/n127 ), .IN3(n2824), .Q(
        n2657) );
  AO21X1 U2452 ( .IN1(n2681), .IN2(n1604), .IN3(n2724), .Q(
        \fpu_div_frac_dp/n1070 ) );
  AO221X1 U2453 ( .IN1(n1883), .IN2(n1774), .IN3(n2738), .IN4(n1522), .IN5(
        n2825), .Q(n2724) );
  AO222X1 U2454 ( .IN1(n2798), .IN2(div_frac_outa[43]), .IN3(n2740), .IN4(
        n2659), .IN5(n2799), .IN6(div_frac_outa[44]), .Q(n2825) );
  XNOR3X1 U2455 ( .IN1(n1478), .IN2(\fpu_div_frac_dp/n130 ), .IN3(n2826), .Q(
        n2659) );
  AO21X1 U2456 ( .IN1(n2681), .IN2(n1615), .IN3(n2725), .Q(
        \fpu_div_frac_dp/n1069 ) );
  AO221X1 U2457 ( .IN1(n1886), .IN2(n1775), .IN3(n2738), .IN4(n1498), .IN5(
        n2827), .Q(n2725) );
  AO222X1 U2458 ( .IN1(n2798), .IN2(div_frac_outa[44]), .IN3(n2740), .IN4(
        n2661), .IN5(n2799), .IN6(div_frac_outa[45]), .Q(n2827) );
  XNOR3X1 U2459 ( .IN1(n1477), .IN2(\fpu_div_frac_dp/n133 ), .IN3(n2828), .Q(
        n2661) );
  AO21X1 U2460 ( .IN1(n2681), .IN2(n1603), .IN3(n2726), .Q(
        \fpu_div_frac_dp/n1068 ) );
  AO221X1 U2461 ( .IN1(n1884), .IN2(n1776), .IN3(n2738), .IN4(n1496), .IN5(
        n2829), .Q(n2726) );
  AO222X1 U2462 ( .IN1(n2798), .IN2(div_frac_outa[45]), .IN3(n2740), .IN4(
        n2663), .IN5(n2799), .IN6(div_frac_outa[46]), .Q(n2829) );
  XNOR3X1 U2463 ( .IN1(n1476), .IN2(\fpu_div_frac_dp/n136 ), .IN3(n2830), .Q(
        n2663) );
  AO21X1 U2464 ( .IN1(n2681), .IN2(n1602), .IN3(n2727), .Q(
        \fpu_div_frac_dp/n1067 ) );
  AO221X1 U2465 ( .IN1(n1885), .IN2(n1777), .IN3(n2738), .IN4(n1515), .IN5(
        n2831), .Q(n2727) );
  AO222X1 U2466 ( .IN1(n2798), .IN2(div_frac_outa[46]), .IN3(n2740), .IN4(
        n2665), .IN5(n2799), .IN6(div_frac_outa[47]), .Q(n2831) );
  XNOR3X1 U2467 ( .IN1(n1475), .IN2(\fpu_div_frac_dp/n139 ), .IN3(n2832), .Q(
        n2665) );
  AO21X1 U2468 ( .IN1(n2681), .IN2(n1614), .IN3(n2728), .Q(
        \fpu_div_frac_dp/n1066 ) );
  AO221X1 U2469 ( .IN1(n1883), .IN2(n1778), .IN3(n2738), .IN4(n1510), .IN5(
        n2833), .Q(n2728) );
  AO222X1 U2470 ( .IN1(n2798), .IN2(div_frac_outa[47]), .IN3(n2740), .IN4(
        n2667), .IN5(n2799), .IN6(div_frac_outa[48]), .Q(n2833) );
  XNOR3X1 U2471 ( .IN1(n1474), .IN2(\fpu_div_frac_dp/n142 ), .IN3(n2834), .Q(
        n2667) );
  AO21X1 U2472 ( .IN1(n2681), .IN2(n1601), .IN3(n2729), .Q(
        \fpu_div_frac_dp/n1065 ) );
  AO221X1 U2473 ( .IN1(n1886), .IN2(n1779), .IN3(n2738), .IN4(n1511), .IN5(
        n2835), .Q(n2729) );
  AO222X1 U2474 ( .IN1(n2798), .IN2(div_frac_outa[48]), .IN3(n2740), .IN4(
        n2669), .IN5(n2799), .IN6(div_frac_outa[49]), .Q(n2835) );
  XNOR3X1 U2475 ( .IN1(n1473), .IN2(\fpu_div_frac_dp/n145 ), .IN3(n2836), .Q(
        n2669) );
  AO21X1 U2476 ( .IN1(n2681), .IN2(n1600), .IN3(n2730), .Q(
        \fpu_div_frac_dp/n1064 ) );
  AO221X1 U2477 ( .IN1(n1884), .IN2(n1780), .IN3(n2738), .IN4(n1523), .IN5(
        n2837), .Q(n2730) );
  AO222X1 U2478 ( .IN1(n2798), .IN2(div_frac_outa[49]), .IN3(n2740), .IN4(
        n2671), .IN5(n2799), .IN6(div_frac_outa[50]), .Q(n2837) );
  XNOR3X1 U2479 ( .IN1(n1472), .IN2(\fpu_div_frac_dp/n148 ), .IN3(n2838), .Q(
        n2671) );
  AO21X1 U2480 ( .IN1(n2681), .IN2(n1613), .IN3(n2731), .Q(
        \fpu_div_frac_dp/n1063 ) );
  AO221X1 U2481 ( .IN1(n1885), .IN2(n1726), .IN3(n2738), .IN4(n1378), .IN5(
        n2839), .Q(n2731) );
  AO222X1 U2482 ( .IN1(n2798), .IN2(div_frac_outa[50]), .IN3(n2740), .IN4(
        n2673), .IN5(n2799), .IN6(div_frac_outa[51]), .Q(n2839) );
  XNOR3X1 U2483 ( .IN1(n1471), .IN2(\fpu_div_frac_dp/n151 ), .IN3(n2840), .Q(
        n2673) );
  AO21X1 U2484 ( .IN1(n2681), .IN2(n1599), .IN3(n2732), .Q(
        \fpu_div_frac_dp/n1062 ) );
  AO221X1 U2485 ( .IN1(n1883), .IN2(n1727), .IN3(n2738), .IN4(n1407), .IN5(
        n2841), .Q(n2732) );
  AO222X1 U2486 ( .IN1(n2798), .IN2(div_frac_outa[51]), .IN3(n2740), .IN4(
        n2675), .IN5(n2799), .IN6(n1383), .Q(n2841) );
  XNOR3X1 U2487 ( .IN1(n1441), .IN2(\fpu_div_frac_dp/n154 ), .IN3(n2842), .Q(
        n2675) );
  AO21X1 U2488 ( .IN1(n2681), .IN2(n1598), .IN3(n2733), .Q(
        \fpu_div_frac_dp/n1061 ) );
  AO221X1 U2489 ( .IN1(n1886), .IN2(n1728), .IN3(n2738), .IN4(n1364), .IN5(
        n2843), .Q(n2733) );
  AO222X1 U2490 ( .IN1(n2799), .IN2(n1529), .IN3(n2798), .IN4(n1383), .IN5(
        n2740), .IN6(n2677), .Q(n2843) );
  XNOR3X1 U2491 ( .IN1(n1440), .IN2(\fpu_div_frac_dp/n158 ), .IN3(n2844), .Q(
        n2677) );
  AND2X1 U2492 ( .IN1(n2010), .IN2(n2796), .Q(n2798) );
  INVX0 U2493 ( .INP(n2017), .ZN(n2796) );
  AND2X1 U2494 ( .IN1(n2010), .IN2(n2017), .Q(n2799) );
  NAND3X0 U2495 ( .IN1(n613), .IN2(n2130), .IN3(\fpu_div_frac_dp/n1 ), .QN(
        n2017) );
  NAND4X0 U2496 ( .IN1(n614), .IN2(n603), .IN3(n2845), .IN4(n2846), .QN(n2130)
         );
  NOR4X0 U2497 ( .IN1(n2847), .IN2(div_exp_out[2]), .IN3(div_exp_out[3]), 
        .IN4(div_exp_out[4]), .QN(n2846) );
  NOR2X0 U2498 ( .IN1(div_exp_out[1]), .IN2(div_exp_out[7]), .QN(n2845) );
  NOR2X0 U2499 ( .IN1(n193), .IN2(se), .QN(n2010) );
  AO21X1 U2500 ( .IN1(n2681), .IN2(n1399), .IN3(n2734), .Q(
        \fpu_div_frac_dp/n1060 ) );
  AO222X1 U2501 ( .IN1(n2740), .IN2(n2679), .IN3(n1884), .IN4(n1718), .IN5(
        n2738), .IN6(n1526), .Q(n2734) );
  XNOR3X1 U2502 ( .IN1(n1439), .IN2(\fpu_div_frac_dp/n163 ), .IN3(n2848), .Q(
        n2679) );
  AO21X1 U2503 ( .IN1(n2681), .IN2(n1443), .IN3(n2735), .Q(
        \fpu_div_frac_dp/n1059 ) );
  AO22X1 U2504 ( .IN1(n2738), .IN2(n1636), .IN3(n2740), .IN4(n2204), .Q(n2735)
         );
  INVX0 U2505 ( .INP(n2009), .ZN(n2204) );
  XNOR3X1 U2506 ( .IN1(n1578), .IN2(n1399), .IN3(n2849), .Q(n2009) );
  AO21X1 U2507 ( .IN1(n2681), .IN2(n1644), .IN3(n2850), .Q(
        \fpu_div_frac_dp/n1058 ) );
  AO21X1 U2508 ( .IN1(n2681), .IN2(n1460), .IN3(n2850), .Q(
        \fpu_div_frac_dp/n1057 ) );
  AO22X1 U2509 ( .IN1(n2738), .IN2(n1637), .IN3(n2740), .IN4(n2564), .Q(n2850)
         );
  XNOR3X1 U2510 ( .IN1(n1443), .IN2(\fpu_div_frac_dp/n166 ), .IN3(n2851), .Q(
        n2564) );
  AND2X1 U2511 ( .IN1(n2852), .IN2(n2570), .Q(n2740) );
  INVX0 U2512 ( .INP(n2853), .ZN(n2570) );
  AND2X1 U2513 ( .IN1(n2852), .IN2(n2853), .Q(n2738) );
  AND3X1 U2514 ( .IN1(n2854), .IN2(n1047), .IN3(n607), .Q(n2852) );
  AND3X1 U2515 ( .IN1(n2855), .IN2(n1047), .IN3(n2559), .Q(n2681) );
  NAND2X0 U2516 ( .IN1(n607), .IN2(n2854), .QN(n2855) );
  AO221X1 U2517 ( .IN1(n2560), .IN2(n1864), .IN3(n2561), .IN4(n1460), .IN5(
        n2856), .Q(\fpu_div_frac_dp/n1056 ) );
  AO221X1 U2518 ( .IN1(n2563), .IN2(n2853), .IN3(n2565), .IN4(n1529), .IN5(
        n2566), .Q(n2856) );
  NAND4X0 U2519 ( .IN1(n2857), .IN2(n2216), .IN3(n613), .IN4(n2105), .QN(n2628) );
  AND3X1 U2520 ( .IN1(n1393), .IN2(n1047), .IN3(n1719), .Q(n2105) );
  AO21X1 U2521 ( .IN1(n2635), .IN2(n1396), .IN3(n2569), .Q(n2565) );
  INVX0 U2522 ( .INP(n2632), .ZN(n2569) );
  NAND2X0 U2523 ( .IN1(n2635), .IN2(n1461), .QN(n2632) );
  AND3X1 U2524 ( .IN1(n939), .IN2(n1047), .IN3(n607), .Q(n2635) );
  XNOR3X1 U2525 ( .IN1(n2858), .IN2(n1644), .IN3(\fpu_div_frac_dp/n165 ), .Q(
        n2853) );
  OA22X1 U2526 ( .IN1(n2859), .IN2(n1443), .IN3(n1635), .IN4(n2851), .Q(n2858)
         );
  AND2X1 U2527 ( .IN1(n2851), .IN2(n1635), .Q(n2859) );
  AO22X1 U2528 ( .IN1(n2849), .IN2(n1399), .IN3(n2860), .IN4(n1578), .Q(n2851)
         );
  OR2X1 U2529 ( .IN1(n2849), .IN2(n1399), .Q(n2860) );
  AO22X1 U2530 ( .IN1(n2848), .IN2(n1598), .IN3(n2861), .IN4(n1439), .Q(n2849)
         );
  OR2X1 U2531 ( .IN1(n1598), .IN2(n2848), .Q(n2861) );
  AO22X1 U2532 ( .IN1(n2844), .IN2(n1599), .IN3(n2862), .IN4(n1440), .Q(n2848)
         );
  OR2X1 U2533 ( .IN1(n1599), .IN2(n2844), .Q(n2862) );
  AO22X1 U2534 ( .IN1(n2842), .IN2(n1613), .IN3(n2863), .IN4(n1441), .Q(n2844)
         );
  OR2X1 U2535 ( .IN1(n1613), .IN2(n2842), .Q(n2863) );
  AO22X1 U2536 ( .IN1(n2840), .IN2(n1600), .IN3(n2864), .IN4(n1471), .Q(n2842)
         );
  OR2X1 U2537 ( .IN1(n1600), .IN2(n2840), .Q(n2864) );
  AO22X1 U2538 ( .IN1(n2838), .IN2(n1601), .IN3(n2865), .IN4(n1472), .Q(n2840)
         );
  OR2X1 U2539 ( .IN1(n1601), .IN2(n2838), .Q(n2865) );
  AO22X1 U2540 ( .IN1(n2836), .IN2(n1614), .IN3(n2866), .IN4(n1473), .Q(n2838)
         );
  OR2X1 U2541 ( .IN1(n1614), .IN2(n2836), .Q(n2866) );
  AO22X1 U2542 ( .IN1(n2834), .IN2(n1602), .IN3(n2867), .IN4(n1474), .Q(n2836)
         );
  OR2X1 U2543 ( .IN1(n1602), .IN2(n2834), .Q(n2867) );
  AO22X1 U2544 ( .IN1(n2832), .IN2(n1603), .IN3(n2868), .IN4(n1475), .Q(n2834)
         );
  OR2X1 U2545 ( .IN1(n1603), .IN2(n2832), .Q(n2868) );
  AO22X1 U2546 ( .IN1(n2830), .IN2(n1615), .IN3(n2869), .IN4(n1476), .Q(n2832)
         );
  OR2X1 U2547 ( .IN1(n1615), .IN2(n2830), .Q(n2869) );
  AO22X1 U2548 ( .IN1(n2828), .IN2(n1604), .IN3(n2870), .IN4(n1477), .Q(n2830)
         );
  OR2X1 U2549 ( .IN1(n1604), .IN2(n2828), .Q(n2870) );
  AO22X1 U2550 ( .IN1(n2826), .IN2(n1605), .IN3(n2871), .IN4(n1478), .Q(n2828)
         );
  OR2X1 U2551 ( .IN1(n1605), .IN2(n2826), .Q(n2871) );
  AO22X1 U2552 ( .IN1(n2824), .IN2(n1616), .IN3(n2872), .IN4(n1479), .Q(n2826)
         );
  OR2X1 U2553 ( .IN1(n1616), .IN2(n2824), .Q(n2872) );
  AO22X1 U2554 ( .IN1(n2822), .IN2(n1606), .IN3(n2873), .IN4(n1480), .Q(n2824)
         );
  OR2X1 U2555 ( .IN1(n1606), .IN2(n2822), .Q(n2873) );
  AO22X1 U2556 ( .IN1(n2820), .IN2(n1607), .IN3(n2874), .IN4(n1481), .Q(n2822)
         );
  OR2X1 U2557 ( .IN1(n1607), .IN2(n2820), .Q(n2874) );
  AO22X1 U2558 ( .IN1(n2818), .IN2(n1617), .IN3(n2875), .IN4(n1482), .Q(n2820)
         );
  OR2X1 U2559 ( .IN1(n1617), .IN2(n2818), .Q(n2875) );
  AO22X1 U2560 ( .IN1(n2816), .IN2(n1608), .IN3(n2876), .IN4(n1483), .Q(n2818)
         );
  OR2X1 U2561 ( .IN1(n1608), .IN2(n2816), .Q(n2876) );
  AO22X1 U2562 ( .IN1(n2814), .IN2(n1609), .IN3(n2877), .IN4(n1484), .Q(n2816)
         );
  OR2X1 U2563 ( .IN1(n1609), .IN2(n2814), .Q(n2877) );
  AO22X1 U2564 ( .IN1(n2812), .IN2(n1618), .IN3(n2878), .IN4(n1485), .Q(n2814)
         );
  OR2X1 U2565 ( .IN1(n1618), .IN2(n2812), .Q(n2878) );
  AO22X1 U2566 ( .IN1(n2810), .IN2(n1610), .IN3(n2879), .IN4(n1486), .Q(n2812)
         );
  OR2X1 U2567 ( .IN1(n1610), .IN2(n2810), .Q(n2879) );
  AO22X1 U2568 ( .IN1(n2808), .IN2(n1611), .IN3(n2880), .IN4(n1487), .Q(n2810)
         );
  OR2X1 U2569 ( .IN1(n1611), .IN2(n2808), .Q(n2880) );
  AO22X1 U2570 ( .IN1(n2806), .IN2(n1619), .IN3(n2881), .IN4(n1488), .Q(n2808)
         );
  OR2X1 U2571 ( .IN1(n1619), .IN2(n2806), .Q(n2881) );
  AO22X1 U2572 ( .IN1(n2804), .IN2(n1624), .IN3(n2882), .IN4(n1462), .Q(n2806)
         );
  OR2X1 U2573 ( .IN1(n1624), .IN2(n2804), .Q(n2882) );
  AO22X1 U2574 ( .IN1(n2802), .IN2(n1612), .IN3(n2883), .IN4(n1442), .Q(n2804)
         );
  OR2X1 U2575 ( .IN1(n1612), .IN2(n2802), .Q(n2883) );
  AO22X1 U2576 ( .IN1(n2800), .IN2(n1625), .IN3(n2884), .IN4(n1463), .Q(n2802)
         );
  OR2X1 U2577 ( .IN1(n1625), .IN2(n2800), .Q(n2884) );
  AO22X1 U2578 ( .IN1(n2794), .IN2(n1626), .IN3(n2885), .IN4(n1464), .Q(n2800)
         );
  OR2X1 U2579 ( .IN1(n1626), .IN2(n2794), .Q(n2885) );
  AO22X1 U2580 ( .IN1(n2792), .IN2(n1627), .IN3(n2886), .IN4(n1465), .Q(n2794)
         );
  OR2X1 U2581 ( .IN1(n1627), .IN2(n2792), .Q(n2886) );
  AO22X1 U2582 ( .IN1(n2790), .IN2(n1628), .IN3(n2887), .IN4(n1466), .Q(n2792)
         );
  OR2X1 U2583 ( .IN1(n1628), .IN2(n2790), .Q(n2887) );
  AO22X1 U2584 ( .IN1(n2788), .IN2(n1629), .IN3(n2888), .IN4(n1467), .Q(n2790)
         );
  OR2X1 U2585 ( .IN1(n1629), .IN2(n2788), .Q(n2888) );
  AO22X1 U2586 ( .IN1(n2786), .IN2(n1630), .IN3(n2889), .IN4(n1468), .Q(n2788)
         );
  OR2X1 U2587 ( .IN1(n1630), .IN2(n2786), .Q(n2889) );
  AO22X1 U2588 ( .IN1(n2784), .IN2(n1631), .IN3(n2890), .IN4(n1469), .Q(n2786)
         );
  OR2X1 U2589 ( .IN1(n1631), .IN2(n2784), .Q(n2890) );
  AO22X1 U2590 ( .IN1(n2782), .IN2(n1632), .IN3(n2891), .IN4(n1470), .Q(n2784)
         );
  OR2X1 U2591 ( .IN1(n1632), .IN2(n2782), .Q(n2891) );
  AO22X1 U2592 ( .IN1(n2780), .IN2(n1444), .IN3(n2892), .IN4(n1581), .Q(n2782)
         );
  OR2X1 U2593 ( .IN1(n1444), .IN2(n2780), .Q(n2892) );
  AO22X1 U2594 ( .IN1(n2778), .IN2(n1445), .IN3(n2893), .IN4(n1587), .Q(n2780)
         );
  OR2X1 U2595 ( .IN1(n1445), .IN2(n2778), .Q(n2893) );
  AO22X1 U2596 ( .IN1(n2776), .IN2(n1446), .IN3(n2894), .IN4(n1582), .Q(n2778)
         );
  OR2X1 U2597 ( .IN1(n1446), .IN2(n2776), .Q(n2894) );
  AO22X1 U2598 ( .IN1(n2774), .IN2(n1447), .IN3(n2895), .IN4(n1583), .Q(n2776)
         );
  OR2X1 U2599 ( .IN1(n1447), .IN2(n2774), .Q(n2895) );
  AO22X1 U2600 ( .IN1(n2772), .IN2(n1448), .IN3(n2896), .IN4(n1588), .Q(n2774)
         );
  OR2X1 U2601 ( .IN1(n1448), .IN2(n2772), .Q(n2896) );
  AO22X1 U2602 ( .IN1(n2770), .IN2(n1449), .IN3(n2897), .IN4(n1584), .Q(n2772)
         );
  OR2X1 U2603 ( .IN1(n1449), .IN2(n2770), .Q(n2897) );
  AO22X1 U2604 ( .IN1(n2768), .IN2(n1450), .IN3(n2898), .IN4(n1585), .Q(n2770)
         );
  OR2X1 U2605 ( .IN1(n1450), .IN2(n2768), .Q(n2898) );
  AO22X1 U2606 ( .IN1(n2766), .IN2(n1451), .IN3(n2899), .IN4(n1589), .Q(n2768)
         );
  OR2X1 U2607 ( .IN1(n1451), .IN2(n2766), .Q(n2899) );
  AO22X1 U2608 ( .IN1(n2764), .IN2(n1452), .IN3(n2900), .IN4(n1586), .Q(n2766)
         );
  OR2X1 U2609 ( .IN1(n1452), .IN2(n2764), .Q(n2900) );
  AO22X1 U2610 ( .IN1(n2762), .IN2(n1453), .IN3(n2901), .IN4(n1590), .Q(n2764)
         );
  OR2X1 U2611 ( .IN1(n1453), .IN2(n2762), .Q(n2901) );
  AO22X1 U2612 ( .IN1(n2760), .IN2(n1454), .IN3(n2902), .IN4(n1591), .Q(n2762)
         );
  OR2X1 U2613 ( .IN1(n1454), .IN2(n2760), .Q(n2902) );
  AO22X1 U2614 ( .IN1(n2758), .IN2(n1455), .IN3(n2903), .IN4(n1592), .Q(n2760)
         );
  OR2X1 U2615 ( .IN1(n1455), .IN2(n2758), .Q(n2903) );
  AO22X1 U2616 ( .IN1(n2756), .IN2(n1456), .IN3(n2904), .IN4(n1593), .Q(n2758)
         );
  OR2X1 U2617 ( .IN1(n1456), .IN2(n2756), .Q(n2904) );
  AO22X1 U2618 ( .IN1(n2754), .IN2(n1457), .IN3(n2905), .IN4(n1594), .Q(n2756)
         );
  OR2X1 U2619 ( .IN1(n1457), .IN2(n2754), .Q(n2905) );
  AO22X1 U2620 ( .IN1(n2752), .IN2(n1458), .IN3(n2906), .IN4(n1595), .Q(n2754)
         );
  OR2X1 U2621 ( .IN1(n1458), .IN2(n2752), .Q(n2906) );
  AO22X1 U2622 ( .IN1(n2750), .IN2(n1459), .IN3(n2907), .IN4(n1596), .Q(n2752)
         );
  OR2X1 U2623 ( .IN1(n1459), .IN2(n2750), .Q(n2907) );
  AO22X1 U2624 ( .IN1(n2748), .IN2(n1620), .IN3(n2908), .IN4(n1434), .Q(n2750)
         );
  OR2X1 U2625 ( .IN1(n1620), .IN2(n2748), .Q(n2908) );
  AO22X1 U2626 ( .IN1(n2746), .IN2(n1621), .IN3(n2909), .IN4(n1435), .Q(n2748)
         );
  OR2X1 U2627 ( .IN1(n1621), .IN2(n2746), .Q(n2909) );
  AO22X1 U2628 ( .IN1(n2744), .IN2(n1622), .IN3(n2910), .IN4(n1436), .Q(n2746)
         );
  OR2X1 U2629 ( .IN1(n1622), .IN2(n2744), .Q(n2910) );
  AO22X1 U2630 ( .IN1(n2742), .IN2(n1623), .IN3(n2911), .IN4(n1437), .Q(n2744)
         );
  OR2X1 U2631 ( .IN1(n1623), .IN2(n2742), .Q(n2911) );
  AO22X1 U2632 ( .IN1(n1527), .IN2(n1683), .IN3(n2912), .IN4(n1373), .Q(n2742)
         );
  NAND2X0 U2633 ( .IN1(\fpu_div_frac_dp/n997 ), .IN2(\fpu_div_frac_dp/n8 ), 
        .QN(n2912) );
  AND3X1 U2634 ( .IN1(n2106), .IN2(n1047), .IN3(n2200), .Q(n2563) );
  INVX0 U2635 ( .INP(n2913), .ZN(n2106) );
  INVX0 U2636 ( .INP(n2631), .ZN(n2561) );
  NAND3X0 U2637 ( .IN1(n2913), .IN2(n1047), .IN3(n2200), .QN(n2631) );
  INVX0 U2638 ( .INP(n2203), .ZN(n2200) );
  NAND2X0 U2639 ( .IN1(n1393), .IN2(n2914), .QN(n2203) );
  NAND3X0 U2640 ( .IN1(n2216), .IN2(n1719), .IN3(n613), .QN(n2914) );
  AO222X1 U2641 ( .IN1(n2107), .IN2(div_exp_out[0]), .IN3(n2847), .IN4(n1391), 
        .IN5(d7stg_fdivd), .IN6(n1371), .Q(n2216) );
  NAND4X0 U2642 ( .IN1(n618), .IN2(n599), .IN3(n584), .IN4(n580), .QN(n2847)
         );
  AND4X1 U2643 ( .IN1(div_exp_out[3]), .IN2(div_exp_out[4]), .IN3(n2915), 
        .IN4(n2916), .Q(n2107) );
  NOR4X0 U2644 ( .IN1(n614), .IN2(n603), .IN3(n598), .IN4(n595), .QN(n2916) );
  OA21X1 U2645 ( .IN1(n2917), .IN2(n1391), .IN3(div_exp_out[2]), .Q(n2915) );
  NOR4X0 U2646 ( .IN1(n599), .IN2(n584), .IN3(n580), .IN4(n22), .QN(n2917) );
  NAND3X0 U2647 ( .IN1(n2918), .IN2(n2919), .IN3(n2058), .QN(n2913) );
  INVX0 U2648 ( .INP(n2857), .ZN(n2058) );
  XOR2X1 U2649 ( .IN1(n593), .IN2(n2920), .Q(n2857) );
  NOR2X0 U2650 ( .IN1(n58), .IN2(n625), .QN(n2920) );
  INVX0 U2651 ( .INP(n2022), .ZN(n2919) );
  NOR2X0 U2652 ( .IN1(n1717), .IN2(n1536), .QN(n2022) );
  NAND2X0 U2653 ( .IN1(n58), .IN2(n2921), .QN(n2918) );
  AO21X1 U2654 ( .IN1(n17), .IN2(n15), .IN3(n16), .Q(n2921) );
  NAND4X0 U2655 ( .IN1(n185), .IN2(n194), .IN3(n2922), .IN4(n1047), .QN(n2633)
         );
  NAND3X0 U2656 ( .IN1(n2923), .IN2(n939), .IN3(n607), .QN(n2922) );
  INVX0 U2657 ( .INP(n2033), .ZN(n939) );
  NAND2X0 U2658 ( .IN1(n611), .IN2(n581), .QN(n2923) );
  AO222X1 U2659 ( .IN1(n2924), .IN2(n2925), .IN3(n2926), .IN4(
        \fpu_div_frac_dp/n602 ), .IN5(n2927), .IN6(n2928), .Q(
        \fpu_div_frac_dp/i_dstg_xtra_regs/N9 ) );
  NAND4X0 U2660 ( .IN1(n2929), .IN2(n2930), .IN3(n2931), .IN4(n2932), .QN(
        n2927) );
  NAND3X0 U2661 ( .IN1(n2933), .IN2(n1403), .IN3(n2934), .QN(n2932) );
  AO21X1 U2662 ( .IN1(n1684), .IN2(n1047), .IN3(
        \fpu_div_frac_dp/i_div_shl_data/N50 ), .Q(n2933) );
  NAND3X0 U2663 ( .IN1(n2935), .IN2(n1410), .IN3(n2936), .QN(n2931) );
  AO21X1 U2664 ( .IN1(\fpu_div_frac_dp/i_div_shl_data/N44 ), .IN2(n1633), 
        .IN3(\fpu_div_frac_dp/i_div_shl_data/N46 ), .Q(n2935) );
  NAND3X0 U2665 ( .IN1(n2937), .IN2(n1368), .IN3(n2938), .QN(n2930) );
  AO21X1 U2666 ( .IN1(n1389), .IN2(n1047), .IN3(
        \fpu_div_frac_dp/i_div_shl_data/N54 ), .Q(n2938) );
  NAND3X0 U2667 ( .IN1(n2939), .IN2(n1400), .IN3(n2940), .QN(n2929) );
  AO21X1 U2668 ( .IN1(n1685), .IN2(n1047), .IN3(
        \fpu_div_frac_dp/i_div_shl_data/N42 ), .Q(n2939) );
  NOR2X0 U2669 ( .IN1(n2941), .IN2(n2942), .QN(n2926) );
  OA221X1 U2670 ( .IN1(\fpu_div_frac_dp/n377 ), .IN2(n2943), .IN3(
        \fpu_div_frac_dp/n2333 ), .IN4(n2944), .IN5(n2945), .Q(n2942) );
  OA21X1 U2671 ( .IN1(\fpu_div_frac_dp/n996 ), .IN2(n1499), .IN3(n1369), .Q(
        n2944) );
  OA221X1 U2672 ( .IN1(n2946), .IN2(n2947), .IN3(n2948), .IN4(n2949), .IN5(
        n2950), .Q(n2941) );
  AO221X1 U2673 ( .IN1(n2951), .IN2(n2952), .IN3(\fpu_div_frac_dp/n364 ), 
        .IN4(n1360), .IN5(\fpu_div_frac_dp/n363 ), .Q(n2950) );
  NAND3X0 U2674 ( .IN1(n2953), .IN2(n1408), .IN3(n2954), .QN(n2952) );
  NAND2X0 U2675 ( .IN1(\fpu_div_frac_dp/n367 ), .IN2(n1580), .QN(n2954) );
  NOR2X0 U2676 ( .IN1(\fpu_div_frac_dp/n988 ), .IN2(n1374), .QN(n2948) );
  AO21X1 U2677 ( .IN1(\fpu_div_frac_dp/n373 ), .IN2(n1528), .IN3(
        \fpu_div_frac_dp/n372 ), .Q(n2947) );
  NAND4X0 U2678 ( .IN1(n2955), .IN2(n2956), .IN3(n2957), .IN4(n2958), .QN(
        n2925) );
  NAND4X0 U2679 ( .IN1(n2959), .IN2(n2960), .IN3(n2961), .IN4(n1649), .QN(
        n2958) );
  AO21X1 U2680 ( .IN1(n1681), .IN2(n1047), .IN3(
        \fpu_div_frac_dp/i_div_shl_data/N26 ), .Q(n2961) );
  NAND4X0 U2681 ( .IN1(n1438), .IN2(n1047), .IN3(n2962), .IN4(n2963), .QN(
        n2957) );
  OA21X1 U2682 ( .IN1(\fpu_div_frac_dp/n981 ), .IN2(n2964), .IN3(n2965), .Q(
        n2963) );
  NAND2X0 U2683 ( .IN1(\fpu_div_frac_dp/n358 ), .IN2(n1597), .QN(n2962) );
  NAND3X0 U2684 ( .IN1(n2966), .IN2(n1367), .IN3(n2967), .QN(n2956) );
  AO21X1 U2685 ( .IN1(n1390), .IN2(n1047), .IN3(
        \fpu_div_frac_dp/i_div_shl_data/N38 ), .Q(n2967) );
  NAND2X0 U2686 ( .IN1(n2968), .IN2(n2969), .QN(n2955) );
  AO21X1 U2687 ( .IN1(\fpu_div_frac_dp/i_div_shl_data/N32 ), .IN2(n1492), 
        .IN3(\fpu_div_frac_dp/i_div_shl_data/N34 ), .Q(n2969) );
  AO22X1 U2688 ( .IN1(\fpu_div_frac_dp/n602 ), .IN2(n2945), .IN3(n2924), .IN4(
        n1047), .Q(\fpu_div_frac_dp/i_dstg_xtra_regs/N7 ) );
  AO22X1 U2689 ( .IN1(n2970), .IN2(n1047), .IN3(n2971), .IN4(
        \fpu_div_frac_dp/n602 ), .Q(\fpu_div_frac_dp/i_dstg_xtra_regs/N6 ) );
  NOR2X0 U2690 ( .IN1(n2945), .IN2(n2953), .QN(n2971) );
  AO22X1 U2691 ( .IN1(n2936), .IN2(n2928), .IN3(n2924), .IN4(n2965), .Q(n2970)
         );
  INVX0 U2692 ( .INP(n2972), .ZN(n2924) );
  OAI22X1 U2693 ( .IN1(n2973), .IN2(n2974), .IN3(n2975), .IN4(n2976), .QN(
        \fpu_div_frac_dp/i_dstg_xtra_regs/N5 ) );
  NAND2X0 U2694 ( .IN1(n2977), .IN2(n1047), .QN(n2976) );
  OA21X1 U2695 ( .IN1(n2978), .IN2(n2979), .IN3(n2980), .Q(n2975) );
  INVX0 U2696 ( .INP(n2934), .ZN(n2980) );
  OA221X1 U2697 ( .IN1(n2965), .IN2(n2966), .IN3(n2964), .IN4(n2981), .IN5(
        n2982), .Q(n2978) );
  INVX0 U2698 ( .INP(n2960), .ZN(n2964) );
  OA22X1 U2699 ( .IN1(n2983), .IN2(n2946), .IN3(n2984), .IN4(n2985), .Q(n2973)
         );
  AND2X1 U2700 ( .IN1(n2943), .IN2(n2945), .Q(n2983) );
  OAI221X1 U2701 ( .IN1(n2974), .IN2(n2986), .IN3(se), .IN4(n2987), .IN5(n2988), .QN(\fpu_div_frac_dp/i_dstg_xtra_regs/N4 ) );
  NAND4X0 U2702 ( .IN1(n2936), .IN2(n2989), .IN3(n2990), .IN4(n2928), .QN(
        n2988) );
  NOR2X0 U2703 ( .IN1(\fpu_div_frac_dp/n984 ), .IN2(\fpu_div_frac_dp/n345 ), 
        .QN(n2990) );
  NAND3X0 U2704 ( .IN1(n2991), .IN2(n2992), .IN3(n2993), .QN(n2989) );
  NAND3X0 U2705 ( .IN1(n1400), .IN2(n1047), .IN3(n1577), .QN(n2993) );
  INVX0 U2706 ( .INP(\fpu_div_frac_dp/i_div_shl_data/N45 ), .ZN(n2992) );
  OA221X1 U2707 ( .IN1(n2994), .IN2(n2972), .IN3(n2995), .IN4(n2996), .IN5(
        n2997), .Q(n2987) );
  NAND3X0 U2708 ( .IN1(n1634), .IN2(n1403), .IN3(n2934), .QN(n2997) );
  NOR2X0 U2709 ( .IN1(n2937), .IN2(n2936), .QN(n2934) );
  NAND2X0 U2710 ( .IN1(n1524), .IN2(n1368), .QN(n2996) );
  NAND2X0 U2711 ( .IN1(n2982), .IN2(n2977), .QN(n2972) );
  OA221X1 U2712 ( .IN1(n2998), .IN2(n2981), .IN3(n2999), .IN4(n3000), .IN5(
        n3001), .Q(n2994) );
  NAND3X0 U2713 ( .IN1(n3002), .IN2(n1388), .IN3(n2968), .QN(n3001) );
  NAND2X0 U2714 ( .IN1(n1525), .IN2(n1367), .QN(n3000) );
  INVX0 U2715 ( .INP(n2966), .ZN(n2999) );
  OA21X1 U2716 ( .IN1(\fpu_div_frac_dp/n360 ), .IN2(\fpu_div_frac_dp/n2330 ), 
        .IN3(n2960), .Q(n2998) );
  AO21X1 U2717 ( .IN1(n2945), .IN2(n3003), .IN3(n3004), .Q(n2986) );
  OA221X1 U2718 ( .IN1(\fpu_div_frac_dp/n988 ), .IN2(n2949), .IN3(n2946), 
        .IN4(n3005), .IN5(n3006), .Q(n3004) );
  NAND3X0 U2719 ( .IN1(n1386), .IN2(n1360), .IN3(n3007), .QN(n3006) );
  NAND2X0 U2720 ( .IN1(n2951), .IN2(n3008), .QN(n3007) );
  NAND3X0 U2721 ( .IN1(n1408), .IN2(n1580), .IN3(n2953), .QN(n3008) );
  NAND2X0 U2722 ( .IN1(n1674), .IN2(n1528), .QN(n3005) );
  NAND3X0 U2723 ( .IN1(n3009), .IN2(n1576), .IN3(n3010), .QN(n2949) );
  NAND3X0 U2724 ( .IN1(n1650), .IN2(n1531), .IN3(n1374), .QN(n3009) );
  NAND3X0 U2725 ( .IN1(n1387), .IN2(n1369), .IN3(n2943), .QN(n3003) );
  NAND4X0 U2726 ( .IN1(n1387), .IN2(n1369), .IN3(n1499), .IN4(n1673), .QN(
        n2943) );
  NOR4X0 U2727 ( .IN1(n2946), .IN2(\fpu_div_frac_dp/n372 ), .IN3(n3011), .IN4(
        \fpu_div_frac_dp/n373 ), .QN(n2945) );
  OR2X1 U2728 ( .IN1(\fpu_div_frac_dp/n983 ), .IN2(\fpu_div_frac_dp/n374 ), 
        .Q(n3011) );
  NAND4X0 U2729 ( .IN1(n3010), .IN2(n1576), .IN3(n3012), .IN4(n1374), .QN(
        n2946) );
  NOR2X0 U2730 ( .IN1(\fpu_div_frac_dp/n988 ), .IN2(\fpu_div_frac_dp/n371 ), 
        .QN(n3012) );
  INVX0 U2731 ( .INP(n2953), .ZN(n3010) );
  NAND2X0 U2732 ( .IN1(n2984), .IN2(n2951), .QN(n2953) );
  INVX0 U2733 ( .INP(n2985), .ZN(n2951) );
  NAND4X0 U2734 ( .IN1(n1386), .IN2(n1535), .IN3(n1675), .IN4(n1360), .QN(
        n2985) );
  NOR4X0 U2735 ( .IN1(\fpu_div_frac_dp/n366 ), .IN2(\fpu_div_frac_dp/n367 ), 
        .IN3(\fpu_div_frac_dp/n368 ), .IN4(\fpu_div_frac_dp/n982 ), .QN(n2984)
         );
  INVX0 U2736 ( .INP(\fpu_div_frac_dp/n602 ), .ZN(n2974) );
  NOR2X0 U2737 ( .IN1(n2977), .IN2(se), .QN(\fpu_div_frac_dp/n602 ) );
  NAND4X0 U2738 ( .IN1(n2960), .IN2(n2982), .IN3(n2959), .IN4(n3013), .QN(
        n2977) );
  NOR4X0 U2739 ( .IN1(\fpu_div_frac_dp/n362 ), .IN2(\fpu_div_frac_dp/n361 ), 
        .IN3(\fpu_div_frac_dp/n360 ), .IN4(\fpu_div_frac_dp/n2330 ), .QN(n3013) );
  INVX0 U2740 ( .INP(n2981), .ZN(n2959) );
  NAND3X0 U2741 ( .IN1(n1438), .IN2(n1597), .IN3(n2965), .QN(n2981) );
  INVX0 U2742 ( .INP(n3002), .ZN(n2965) );
  NAND4X0 U2743 ( .IN1(n2968), .IN2(n1388), .IN3(n1492), .IN4(n1680), .QN(
        n3002) );
  NOR2X0 U2744 ( .IN1(n2966), .IN2(\fpu_div_frac_dp/n354 ), .QN(n2968) );
  NAND4X0 U2745 ( .IN1(n1525), .IN2(n1367), .IN3(n1390), .IN4(n1678), .QN(
        n2966) );
  INVX0 U2746 ( .INP(n2928), .ZN(n2982) );
  NAND4X0 U2747 ( .IN1(n2940), .IN2(n1577), .IN3(n3014), .IN4(n1400), .QN(
        n2928) );
  NOR2X0 U2748 ( .IN1(\fpu_div_frac_dp/n350 ), .IN2(\fpu_div_frac_dp/n349 ), 
        .QN(n3014) );
  INVX0 U2749 ( .INP(n2979), .ZN(n2940) );
  NAND4X0 U2750 ( .IN1(n2936), .IN2(n1410), .IN3(n3015), .IN4(n1633), .QN(
        n2979) );
  NOR2X0 U2751 ( .IN1(\fpu_div_frac_dp/n984 ), .IN2(\fpu_div_frac_dp/n347 ), 
        .QN(n3015) );
  AND4X1 U2752 ( .IN1(n2995), .IN2(n1634), .IN3(n3016), .IN4(n1403), .Q(n2936)
         );
  NOR2X0 U2753 ( .IN1(\fpu_div_frac_dp/n344 ), .IN2(\fpu_div_frac_dp/n343 ), 
        .QN(n3016) );
  INVX0 U2754 ( .INP(n2937), .ZN(n2995) );
  NAND4X0 U2755 ( .IN1(n1524), .IN2(n1368), .IN3(n1389), .IN4(n1677), .QN(
        n2937) );
  NOR2X0 U2756 ( .IN1(\fpu_div_frac_dp/n358 ), .IN2(\fpu_div_frac_dp/n359 ), 
        .QN(n2960) );
  AND2X1 U2757 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n373 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N9 ) );
  AND2X1 U2758 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n374 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N8 ) );
  NOR2X0 U2759 ( .IN1(se), .IN2(n1387), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N7 ) );
  NOR2X0 U2760 ( .IN1(se), .IN2(n1369), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N6 ) );
  NOR2X0 U2761 ( .IN1(se), .IN2(n1368), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N55 ) );
  NOR2X0 U2762 ( .IN1(n1524), .IN2(se), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N54 ) );
  NOR2X0 U2763 ( .IN1(se), .IN2(n1389), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N53 ) );
  NOR2X0 U2764 ( .IN1(se), .IN2(n1677), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N52 ) );
  NOR2X0 U2765 ( .IN1(se), .IN2(n1403), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N51 ) );
  NOR2X0 U2766 ( .IN1(n1634), .IN2(se), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N50 ) );
  NOR2X0 U2767 ( .IN1(se), .IN2(n1673), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N5 ) );
  NOR2X0 U2768 ( .IN1(se), .IN2(n1684), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N49 ) );
  AND2X1 U2769 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n344 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N48 ) );
  NOR2X0 U2770 ( .IN1(se), .IN2(n1410), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N47 ) );
  AND2X1 U2771 ( .IN1(\fpu_div_frac_dp/n984 ), .IN2(n1047), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N46 ) );
  NOR2X0 U2772 ( .IN1(n1633), .IN2(se), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N45 ) );
  INVX0 U2773 ( .INP(n2991), .ZN(\fpu_div_frac_dp/i_div_shl_data/N44 ) );
  NAND2X0 U2774 ( .IN1(\fpu_div_frac_dp/n347 ), .IN2(n1047), .QN(n2991) );
  NOR2X0 U2775 ( .IN1(se), .IN2(n1400), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N43 ) );
  NOR2X0 U2776 ( .IN1(n1577), .IN2(se), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N42 ) );
  NOR2X0 U2777 ( .IN1(se), .IN2(n1685), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N41 ) );
  AND2X1 U2778 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n350 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N40 ) );
  NOR2X0 U2779 ( .IN1(se), .IN2(n1499), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N4 ) );
  NOR2X0 U2780 ( .IN1(se), .IN2(n1367), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N39 ) );
  NOR2X0 U2781 ( .IN1(n1525), .IN2(se), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N38 ) );
  NOR2X0 U2782 ( .IN1(se), .IN2(n1390), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N37 ) );
  NOR2X0 U2783 ( .IN1(se), .IN2(n1678), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N36 ) );
  AND2X1 U2784 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n354 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N35 ) );
  NOR2X0 U2785 ( .IN1(n1388), .IN2(se), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N34 ) );
  NOR2X0 U2786 ( .IN1(se), .IN2(n1492), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N33 ) );
  NOR2X0 U2787 ( .IN1(n1680), .IN2(se), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N32 ) );
  NOR2X0 U2788 ( .IN1(se), .IN2(n1438), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N31 ) );
  AND2X1 U2789 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n377 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N3 ) );
  AND2X1 U2790 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n358 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N29 ) );
  AND2X1 U2791 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n359 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N28 ) );
  NOR2X0 U2792 ( .IN1(se), .IN2(n1649), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N27 ) );
  AND2X1 U2793 ( .IN1(\fpu_div_frac_dp/n2330 ), .IN2(n1047), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N26 ) );
  NOR2X0 U2794 ( .IN1(se), .IN2(n1681), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N25 ) );
  AND2X1 U2795 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n362 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N24 ) );
  NOR2X0 U2796 ( .IN1(se), .IN2(n1386), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N23 ) );
  NOR2X0 U2797 ( .IN1(se), .IN2(n1360), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N22 ) );
  NOR2X0 U2798 ( .IN1(se), .IN2(n1535), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N21 ) );
  NOR2X0 U2799 ( .IN1(se), .IN2(n1675), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N20 ) );
  NOR2X0 U2800 ( .IN1(se), .IN2(n1408), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N19 ) );
  NOR2X0 U2801 ( .IN1(se), .IN2(n1580), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N18 ) );
  AND2X1 U2802 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n367 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N17 ) );
  AND2X1 U2803 ( .IN1(n1047), .IN2(\fpu_div_frac_dp/n368 ), .Q(
        \fpu_div_frac_dp/i_div_shl_data/N16 ) );
  NOR2X0 U2804 ( .IN1(se), .IN2(n1576), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N15 ) );
  NOR2X0 U2805 ( .IN1(se), .IN2(n1531), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N14 ) );
  NOR2X0 U2806 ( .IN1(se), .IN2(n1374), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N13 ) );
  NOR2X0 U2807 ( .IN1(se), .IN2(n1650), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N12 ) );
  NOR2X0 U2808 ( .IN1(se), .IN2(n1674), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N11 ) );
  NOR2X0 U2809 ( .IN1(se), .IN2(n1528), .QN(
        \fpu_div_frac_dp/i_div_shl_data/N10 ) );
  OA221X1 U2810 ( .IN1(n3017), .IN2(n3018), .IN3(\fpu_div_frac_dp/n481 ), 
        .IN4(n3019), .IN5(n3020), .Q(\fpu_div_frac_dp/i_div_norm_inv/N9 ) );
  OA22X1 U2811 ( .IN1(\fpu_div_frac_dp/n427 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n482 ), .IN4(n3022), .Q(n3020) );
  NOR2X0 U2812 ( .IN1(n3023), .IN2(n1686), .QN(n3017) );
  OA221X1 U2813 ( .IN1(n3024), .IN2(n3018), .IN3(\fpu_div_frac_dp/n482 ), 
        .IN4(n3019), .IN5(n3025), .Q(\fpu_div_frac_dp/i_div_norm_inv/N8 ) );
  OA22X1 U2814 ( .IN1(\fpu_div_frac_dp/n428 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n483 ), .IN4(n3022), .Q(n3025) );
  NOR2X0 U2815 ( .IN1(n3023), .IN2(n1687), .QN(n3024) );
  OA221X1 U2816 ( .IN1(n3026), .IN2(n3018), .IN3(\fpu_div_frac_dp/n483 ), 
        .IN4(n3019), .IN5(n3027), .Q(\fpu_div_frac_dp/i_div_norm_inv/N7 ) );
  OA22X1 U2817 ( .IN1(\fpu_div_frac_dp/n429 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n484 ), .IN4(n3022), .Q(n3027) );
  NOR2X0 U2818 ( .IN1(n3023), .IN2(n1688), .QN(n3026) );
  OA221X1 U2819 ( .IN1(n3028), .IN2(n3018), .IN3(\fpu_div_frac_dp/n484 ), 
        .IN4(n3019), .IN5(n3029), .Q(\fpu_div_frac_dp/i_div_norm_inv/N6 ) );
  OA22X1 U2820 ( .IN1(\fpu_div_frac_dp/n430 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n485 ), .IN4(n3022), .Q(n3029) );
  NOR2X0 U2821 ( .IN1(n3023), .IN2(n1689), .QN(n3028) );
  NOR4X0 U2822 ( .IN1(n3030), .IN2(n3031), .IN3(n3032), .IN4(n3033), .QN(
        \fpu_div_frac_dp/i_div_norm_inv/N55 ) );
  OAI221X1 U2823 ( .IN1(n3021), .IN2(\fpu_div_frac_dp/n381 ), .IN3(n3022), 
        .IN4(\fpu_div_frac_dp/n436 ), .IN5(n3034), .QN(n3031) );
  NAND4X0 U2824 ( .IN1(n3035), .IN2(n3019), .IN3(n3036), .IN4(n3037), .QN(
        n3030) );
  OA222X1 U2825 ( .IN1(\fpu_div_frac_dp/n433 ), .IN2(n3038), .IN3(n2187), 
        .IN4(n3039), .IN5(n3040), .IN6(n1549), .Q(n3037) );
  OA22X1 U2826 ( .IN1(n253), .IN2(n2043), .IN3(n2054), .IN4(n3041), .Q(n3039)
         );
  OA21X1 U2827 ( .IN1(n1731), .IN2(n1538), .IN3(n585), .Q(n2054) );
  NAND2X0 U2828 ( .IN1(n35), .IN2(n1356), .QN(n2043) );
  AO21X1 U2829 ( .IN1(n52), .IN2(n37), .IN3(n1543), .Q(n35) );
  OR2X1 U2830 ( .IN1(n3042), .IN2(\fpu_div_frac_dp/n378 ), .Q(n3036) );
  AND4X1 U2831 ( .IN1(n3043), .IN2(n3044), .IN3(n3045), .IN4(n3046), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N54 ) );
  OA222X1 U2832 ( .IN1(\fpu_div_frac_dp/n437 ), .IN2(n3022), .IN3(n370), .IN4(
        n3047), .IN5(n3035), .IN6(n3048), .Q(n3046) );
  OA222X1 U2833 ( .IN1(\fpu_div_frac_dp/n434 ), .IN2(n3038), .IN3(n3034), 
        .IN4(n3049), .IN5(n3050), .IN6(n3019), .Q(n3045) );
  NOR2X0 U2834 ( .IN1(n3051), .IN2(n1670), .QN(n3050) );
  NOR2X0 U2835 ( .IN1(n3052), .IN2(n1671), .QN(n3049) );
  OA222X1 U2836 ( .IN1(\fpu_div_frac_dp/n379 ), .IN2(n3042), .IN3(
        \fpu_div_frac_dp/n433 ), .IN4(n3035), .IN5(\fpu_div_frac_dp/n382 ), 
        .IN6(n3021), .Q(n3044) );
  OA21X1 U2837 ( .IN1(\fpu_div_frac_dp/n378 ), .IN2(n3047), .IN3(n3053), .Q(
        n3043) );
  AND3X1 U2838 ( .IN1(n3054), .IN2(n3055), .IN3(n3056), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N53 ) );
  OA221X1 U2839 ( .IN1(\fpu_div_frac_dp/n437 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n379 ), .IN5(n3057), .Q(n3056) );
  OA22X1 U2840 ( .IN1(\fpu_div_frac_dp/n435 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n380 ), .IN4(n3042), .Q(n3057) );
  OA22X1 U2841 ( .IN1(\fpu_div_frac_dp/n438 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n382 ), .Q(n3055) );
  OA22X1 U2842 ( .IN1(n3058), .IN2(n3059), .IN3(\fpu_div_frac_dp/n434 ), .IN4(
        n3035), .Q(n3054) );
  NOR2X0 U2843 ( .IN1(n3033), .IN2(n1653), .QN(n3058) );
  AND3X1 U2844 ( .IN1(n3060), .IN2(n3061), .IN3(n3062), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N52 ) );
  OA221X1 U2845 ( .IN1(\fpu_div_frac_dp/n438 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n380 ), .IN5(n3063), .Q(n3062) );
  OA22X1 U2846 ( .IN1(\fpu_div_frac_dp/n436 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n381 ), .IN4(n3042), .Q(n3063) );
  OA22X1 U2847 ( .IN1(\fpu_div_frac_dp/n439 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n383 ), .Q(n3061) );
  OA22X1 U2848 ( .IN1(n3064), .IN2(n3059), .IN3(\fpu_div_frac_dp/n435 ), .IN4(
        n3035), .Q(n3060) );
  NOR2X0 U2849 ( .IN1(n3033), .IN2(n1654), .QN(n3064) );
  AND3X1 U2850 ( .IN1(n3065), .IN2(n3066), .IN3(n3067), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N51 ) );
  OA221X1 U2851 ( .IN1(\fpu_div_frac_dp/n439 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n381 ), .IN5(n3068), .Q(n3067) );
  OA22X1 U2852 ( .IN1(\fpu_div_frac_dp/n437 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n382 ), .IN4(n3042), .Q(n3068) );
  OA22X1 U2853 ( .IN1(\fpu_div_frac_dp/n440 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n384 ), .Q(n3066) );
  OA22X1 U2854 ( .IN1(n3069), .IN2(n3059), .IN3(\fpu_div_frac_dp/n436 ), .IN4(
        n3035), .Q(n3065) );
  NOR2X0 U2855 ( .IN1(n3033), .IN2(n1655), .QN(n3069) );
  AND3X1 U2856 ( .IN1(n3070), .IN2(n3071), .IN3(n3072), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N50 ) );
  OA221X1 U2857 ( .IN1(\fpu_div_frac_dp/n440 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n382 ), .IN5(n3073), .Q(n3072) );
  OA22X1 U2858 ( .IN1(\fpu_div_frac_dp/n438 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n383 ), .IN4(n3042), .Q(n3073) );
  OA22X1 U2859 ( .IN1(\fpu_div_frac_dp/n441 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n385 ), .Q(n3071) );
  OA22X1 U2860 ( .IN1(n3074), .IN2(n3059), .IN3(\fpu_div_frac_dp/n437 ), .IN4(
        n3035), .Q(n3070) );
  NOR2X0 U2861 ( .IN1(n3033), .IN2(n1656), .QN(n3074) );
  OA221X1 U2862 ( .IN1(n3075), .IN2(n3018), .IN3(\fpu_div_frac_dp/n485 ), 
        .IN4(n3019), .IN5(n3076), .Q(\fpu_div_frac_dp/i_div_norm_inv/N5 ) );
  OA22X1 U2863 ( .IN1(\fpu_div_frac_dp/n431 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n486 ), .IN4(n3022), .Q(n3076) );
  NOR2X0 U2864 ( .IN1(n3023), .IN2(n1690), .QN(n3075) );
  AND3X1 U2865 ( .IN1(n3077), .IN2(n3078), .IN3(n3079), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N49 ) );
  OA221X1 U2866 ( .IN1(\fpu_div_frac_dp/n441 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n383 ), .IN5(n3080), .Q(n3079) );
  OA22X1 U2867 ( .IN1(\fpu_div_frac_dp/n439 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n384 ), .IN4(n3042), .Q(n3080) );
  OA22X1 U2868 ( .IN1(\fpu_div_frac_dp/n442 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n386 ), .Q(n3078) );
  OA22X1 U2869 ( .IN1(n3081), .IN2(n3059), .IN3(\fpu_div_frac_dp/n438 ), .IN4(
        n3035), .Q(n3077) );
  NOR2X0 U2870 ( .IN1(n3033), .IN2(n1657), .QN(n3081) );
  AND3X1 U2871 ( .IN1(n3082), .IN2(n3083), .IN3(n3084), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N48 ) );
  OA221X1 U2872 ( .IN1(\fpu_div_frac_dp/n442 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n384 ), .IN5(n3085), .Q(n3084) );
  OA22X1 U2873 ( .IN1(\fpu_div_frac_dp/n440 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n385 ), .IN4(n3042), .Q(n3085) );
  OA22X1 U2874 ( .IN1(\fpu_div_frac_dp/n443 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n387 ), .Q(n3083) );
  OA22X1 U2875 ( .IN1(n3086), .IN2(n3059), .IN3(\fpu_div_frac_dp/n439 ), .IN4(
        n3035), .Q(n3082) );
  NOR2X0 U2876 ( .IN1(n3033), .IN2(n1658), .QN(n3086) );
  AND3X1 U2877 ( .IN1(n3087), .IN2(n3088), .IN3(n3089), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N47 ) );
  OA221X1 U2878 ( .IN1(\fpu_div_frac_dp/n443 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n385 ), .IN5(n3090), .Q(n3089) );
  OA22X1 U2879 ( .IN1(\fpu_div_frac_dp/n441 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n386 ), .IN4(n3042), .Q(n3090) );
  OA22X1 U2880 ( .IN1(\fpu_div_frac_dp/n444 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n388 ), .Q(n3088) );
  OA22X1 U2881 ( .IN1(n3091), .IN2(n3059), .IN3(\fpu_div_frac_dp/n440 ), .IN4(
        n3035), .Q(n3087) );
  NOR2X0 U2882 ( .IN1(n3033), .IN2(n1659), .QN(n3091) );
  AND3X1 U2883 ( .IN1(n3092), .IN2(n3093), .IN3(n3094), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N46 ) );
  OA221X1 U2884 ( .IN1(\fpu_div_frac_dp/n444 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n386 ), .IN5(n3095), .Q(n3094) );
  OA22X1 U2885 ( .IN1(\fpu_div_frac_dp/n442 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n387 ), .IN4(n3042), .Q(n3095) );
  OA22X1 U2886 ( .IN1(\fpu_div_frac_dp/n445 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n389 ), .Q(n3093) );
  OA22X1 U2887 ( .IN1(n3096), .IN2(n3059), .IN3(\fpu_div_frac_dp/n441 ), .IN4(
        n3035), .Q(n3092) );
  NOR2X0 U2888 ( .IN1(n3033), .IN2(n1660), .QN(n3096) );
  AND3X1 U2889 ( .IN1(n3097), .IN2(n3098), .IN3(n3099), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N45 ) );
  OA221X1 U2890 ( .IN1(\fpu_div_frac_dp/n445 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n387 ), .IN5(n3100), .Q(n3099) );
  OA22X1 U2891 ( .IN1(\fpu_div_frac_dp/n443 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n388 ), .IN4(n3042), .Q(n3100) );
  OA22X1 U2892 ( .IN1(\fpu_div_frac_dp/n446 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n390 ), .Q(n3098) );
  OA22X1 U2893 ( .IN1(n3101), .IN2(n3059), .IN3(\fpu_div_frac_dp/n442 ), .IN4(
        n3035), .Q(n3097) );
  NOR2X0 U2894 ( .IN1(n3033), .IN2(n1661), .QN(n3101) );
  AND3X1 U2895 ( .IN1(n3102), .IN2(n3103), .IN3(n3104), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N44 ) );
  OA221X1 U2896 ( .IN1(\fpu_div_frac_dp/n446 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n388 ), .IN5(n3105), .Q(n3104) );
  OA22X1 U2897 ( .IN1(\fpu_div_frac_dp/n444 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n389 ), .IN4(n3042), .Q(n3105) );
  OA22X1 U2898 ( .IN1(\fpu_div_frac_dp/n447 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n391 ), .Q(n3103) );
  OA22X1 U2899 ( .IN1(n3106), .IN2(n3059), .IN3(\fpu_div_frac_dp/n443 ), .IN4(
        n3035), .Q(n3102) );
  NOR2X0 U2900 ( .IN1(n3033), .IN2(n1662), .QN(n3106) );
  AND3X1 U2901 ( .IN1(n3107), .IN2(n3108), .IN3(n3109), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N43 ) );
  OA221X1 U2902 ( .IN1(\fpu_div_frac_dp/n447 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n389 ), .IN5(n3110), .Q(n3109) );
  OA22X1 U2903 ( .IN1(\fpu_div_frac_dp/n445 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n390 ), .IN4(n3042), .Q(n3110) );
  OA22X1 U2904 ( .IN1(\fpu_div_frac_dp/n448 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n392 ), .Q(n3108) );
  OA22X1 U2905 ( .IN1(n3111), .IN2(n3059), .IN3(\fpu_div_frac_dp/n444 ), .IN4(
        n3035), .Q(n3107) );
  NOR2X0 U2906 ( .IN1(n3033), .IN2(n1663), .QN(n3111) );
  AND3X1 U2907 ( .IN1(n3112), .IN2(n3113), .IN3(n3114), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N42 ) );
  OA221X1 U2908 ( .IN1(\fpu_div_frac_dp/n448 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n390 ), .IN5(n3115), .Q(n3114) );
  OA22X1 U2909 ( .IN1(\fpu_div_frac_dp/n446 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n391 ), .IN4(n3042), .Q(n3115) );
  OA22X1 U2910 ( .IN1(\fpu_div_frac_dp/n449 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n393 ), .Q(n3113) );
  OA22X1 U2911 ( .IN1(n3116), .IN2(n3059), .IN3(\fpu_div_frac_dp/n445 ), .IN4(
        n3035), .Q(n3112) );
  NOR2X0 U2912 ( .IN1(n3033), .IN2(n1664), .QN(n3116) );
  AND3X1 U2913 ( .IN1(n3117), .IN2(n3118), .IN3(n3119), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N41 ) );
  OA221X1 U2914 ( .IN1(\fpu_div_frac_dp/n449 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n391 ), .IN5(n3120), .Q(n3119) );
  OA22X1 U2915 ( .IN1(\fpu_div_frac_dp/n447 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n392 ), .IN4(n3042), .Q(n3120) );
  OA22X1 U2916 ( .IN1(\fpu_div_frac_dp/n450 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n394 ), .Q(n3118) );
  OA22X1 U2917 ( .IN1(n3121), .IN2(n3059), .IN3(\fpu_div_frac_dp/n446 ), .IN4(
        n3035), .Q(n3117) );
  NOR2X0 U2918 ( .IN1(n3033), .IN2(n1665), .QN(n3121) );
  AND3X1 U2919 ( .IN1(n3122), .IN2(n3123), .IN3(n3124), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N40 ) );
  OA221X1 U2920 ( .IN1(\fpu_div_frac_dp/n450 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n392 ), .IN5(n3125), .Q(n3124) );
  OA22X1 U2921 ( .IN1(\fpu_div_frac_dp/n448 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n393 ), .IN4(n3042), .Q(n3125) );
  OA22X1 U2922 ( .IN1(\fpu_div_frac_dp/n451 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n395 ), .Q(n3123) );
  OA22X1 U2923 ( .IN1(n3126), .IN2(n3059), .IN3(\fpu_div_frac_dp/n447 ), .IN4(
        n3035), .Q(n3122) );
  NOR2X0 U2924 ( .IN1(n3033), .IN2(n1666), .QN(n3126) );
  OA221X1 U2925 ( .IN1(n3127), .IN2(n3018), .IN3(\fpu_div_frac_dp/n486 ), 
        .IN4(n3019), .IN5(n3128), .Q(\fpu_div_frac_dp/i_div_norm_inv/N4 ) );
  OA22X1 U2926 ( .IN1(\fpu_div_frac_dp/n432 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n487 ), .IN4(n3022), .Q(n3128) );
  NOR2X0 U2927 ( .IN1(n3023), .IN2(n1691), .QN(n3127) );
  AND3X1 U2928 ( .IN1(n3129), .IN2(n3130), .IN3(n3131), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N39 ) );
  OA221X1 U2929 ( .IN1(\fpu_div_frac_dp/n451 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n393 ), .IN5(n3132), .Q(n3131) );
  OA22X1 U2930 ( .IN1(\fpu_div_frac_dp/n449 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n394 ), .IN4(n3042), .Q(n3132) );
  OA22X1 U2931 ( .IN1(\fpu_div_frac_dp/n452 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n396 ), .Q(n3130) );
  OA22X1 U2932 ( .IN1(n3133), .IN2(n3059), .IN3(\fpu_div_frac_dp/n448 ), .IN4(
        n3035), .Q(n3129) );
  NOR2X0 U2933 ( .IN1(n3033), .IN2(n1667), .QN(n3133) );
  AND3X1 U2934 ( .IN1(n3134), .IN2(n3135), .IN3(n3136), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N38 ) );
  OA221X1 U2935 ( .IN1(\fpu_div_frac_dp/n452 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n394 ), .IN5(n3137), .Q(n3136) );
  OA22X1 U2936 ( .IN1(\fpu_div_frac_dp/n450 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n395 ), .IN4(n3042), .Q(n3137) );
  OA22X1 U2937 ( .IN1(\fpu_div_frac_dp/n453 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n397 ), .Q(n3135) );
  OA22X1 U2938 ( .IN1(n3138), .IN2(n3059), .IN3(\fpu_div_frac_dp/n449 ), .IN4(
        n3035), .Q(n3134) );
  NOR2X0 U2939 ( .IN1(n3033), .IN2(n1668), .QN(n3138) );
  AND3X1 U2940 ( .IN1(n3139), .IN2(n3140), .IN3(n3141), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N37 ) );
  OA221X1 U2941 ( .IN1(\fpu_div_frac_dp/n453 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n395 ), .IN5(n3142), .Q(n3141) );
  OA22X1 U2942 ( .IN1(\fpu_div_frac_dp/n451 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n396 ), .IN4(n3042), .Q(n3142) );
  OA22X1 U2943 ( .IN1(\fpu_div_frac_dp/n454 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n398 ), .Q(n3140) );
  OA22X1 U2944 ( .IN1(n3143), .IN2(n3059), .IN3(\fpu_div_frac_dp/n450 ), .IN4(
        n3035), .Q(n3139) );
  NOR2X0 U2945 ( .IN1(n3033), .IN2(n1669), .QN(n3143) );
  AND3X1 U2946 ( .IN1(n3144), .IN2(n3145), .IN3(n3146), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N36 ) );
  OA221X1 U2947 ( .IN1(\fpu_div_frac_dp/n454 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n396 ), .IN5(n3147), .Q(n3146) );
  OA22X1 U2948 ( .IN1(\fpu_div_frac_dp/n452 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n397 ), .IN4(n3042), .Q(n3147) );
  OA22X1 U2949 ( .IN1(\fpu_div_frac_dp/n455 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n399 ), .Q(n3145) );
  OA22X1 U2950 ( .IN1(n3148), .IN2(n3059), .IN3(\fpu_div_frac_dp/n451 ), .IN4(
        n3035), .Q(n3144) );
  NOR2X0 U2951 ( .IN1(n3033), .IN2(n1652), .QN(n3148) );
  AND3X1 U2952 ( .IN1(n3149), .IN2(n3150), .IN3(n3151), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N35 ) );
  OA221X1 U2953 ( .IN1(\fpu_div_frac_dp/n455 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n397 ), .IN5(n3152), .Q(n3151) );
  OA22X1 U2954 ( .IN1(\fpu_div_frac_dp/n453 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n398 ), .IN4(n3042), .Q(n3152) );
  OA22X1 U2955 ( .IN1(\fpu_div_frac_dp/n456 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n400 ), .Q(n3150) );
  OA22X1 U2956 ( .IN1(n3153), .IN2(n3059), .IN3(\fpu_div_frac_dp/n452 ), .IN4(
        n3035), .Q(n3149) );
  NOR2X0 U2957 ( .IN1(n3033), .IN2(n1711), .QN(n3153) );
  AND3X1 U2958 ( .IN1(n3154), .IN2(n3155), .IN3(n3156), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N34 ) );
  OA221X1 U2959 ( .IN1(\fpu_div_frac_dp/n456 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n398 ), .IN5(n3157), .Q(n3156) );
  OA22X1 U2960 ( .IN1(\fpu_div_frac_dp/n454 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n399 ), .IN4(n3042), .Q(n3157) );
  OA22X1 U2961 ( .IN1(\fpu_div_frac_dp/n457 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n401 ), .Q(n3155) );
  OA22X1 U2962 ( .IN1(n3158), .IN2(n3059), .IN3(\fpu_div_frac_dp/n453 ), .IN4(
        n3035), .Q(n3154) );
  NOR2X0 U2963 ( .IN1(n3033), .IN2(n1712), .QN(n3158) );
  AND3X1 U2964 ( .IN1(n3159), .IN2(n3160), .IN3(n3161), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N33 ) );
  OA221X1 U2965 ( .IN1(\fpu_div_frac_dp/n457 ), .IN2(n3019), .IN3(n3047), 
        .IN4(\fpu_div_frac_dp/n399 ), .IN5(n3162), .Q(n3161) );
  OA22X1 U2966 ( .IN1(\fpu_div_frac_dp/n455 ), .IN2(n3038), .IN3(
        \fpu_div_frac_dp/n400 ), .IN4(n3042), .Q(n3162) );
  NAND2X0 U2967 ( .IN1(n3163), .IN2(\fpu_div_ctl/d2stg_denorm_sng_in2 ), .QN(
        n3042) );
  NAND4X0 U2968 ( .IN1(n3164), .IN2(n604), .IN3(n3165), .IN4(n352), .QN(n3038)
         );
  AND2X1 U2969 ( .IN1(n1643), .IN2(n370), .Q(n3165) );
  OA22X1 U2970 ( .IN1(\fpu_div_frac_dp/n458 ), .IN2(n3022), .IN3(n3034), .IN4(
        \fpu_div_frac_dp/n402 ), .Q(n3160) );
  OA22X1 U2971 ( .IN1(n3166), .IN2(n3059), .IN3(\fpu_div_frac_dp/n454 ), .IN4(
        n3035), .Q(n3159) );
  NOR2X0 U2972 ( .IN1(n3033), .IN2(n3167), .QN(n3059) );
  NOR2X0 U2973 ( .IN1(n3033), .IN2(n1714), .QN(n3166) );
  AND3X1 U2974 ( .IN1(n3168), .IN2(n3053), .IN3(n3169), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N32 ) );
  OA221X1 U2975 ( .IN1(\fpu_div_frac_dp/n455 ), .IN2(n3035), .IN3(n3034), 
        .IN4(\fpu_div_frac_dp/n403 ), .IN5(n3170), .Q(n3169) );
  OA22X1 U2976 ( .IN1(n3047), .IN2(\fpu_div_frac_dp/n400 ), .IN3(
        \fpu_div_frac_dp/n404 ), .IN4(n3021), .Q(n3170) );
  INVX0 U2977 ( .INP(n3032), .ZN(n3047) );
  AO22X1 U2978 ( .IN1(n3163), .IN2(\fpu_div_ctl/d2stg_norm_sng_in2 ), .IN3(
        n3171), .IN4(n3172), .Q(n3032) );
  NAND2X0 U2979 ( .IN1(n370), .IN2(n3173), .QN(n3171) );
  NAND4X0 U2980 ( .IN1(n3164), .IN2(n3173), .IN3(n3174), .IN4(n370), .QN(n3035) );
  NAND4X0 U2981 ( .IN1(n621), .IN2(n585), .IN3(n1679), .IN4(n1376), .QN(n370)
         );
  NOR2X0 U2982 ( .IN1(n604), .IN2(n50), .QN(n3174) );
  NAND2X0 U2983 ( .IN1(n3048), .IN2(n3175), .QN(n3173) );
  INVX0 U2984 ( .INP(n352), .ZN(n3175) );
  NAND3X0 U2985 ( .IN1(n1376), .IN2(n1645), .IN3(n585), .QN(n352) );
  INVX0 U2986 ( .INP(n3033), .ZN(n3053) );
  NAND2X0 U2987 ( .IN1(n3176), .IN2(n1047), .QN(n3033) );
  OA22X1 U2988 ( .IN1(\fpu_div_frac_dp/n459 ), .IN2(n3022), .IN3(
        \fpu_div_frac_dp/n458 ), .IN4(n3019), .Q(n3168) );
  OA221X1 U2989 ( .IN1(n3177), .IN2(n3018), .IN3(\fpu_div_frac_dp/n459 ), 
        .IN4(n3019), .IN5(n3178), .Q(\fpu_div_frac_dp/i_div_norm_inv/N31 ) );
  OA22X1 U2990 ( .IN1(\fpu_div_frac_dp/n405 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n460 ), .IN4(n3022), .Q(n3178) );
  NOR2X0 U2991 ( .IN1(n3023), .IN2(n1713), .QN(n3177) );
  OA221X1 U2992 ( .IN1(n3179), .IN2(n3018), .IN3(\fpu_div_frac_dp/n460 ), 
        .IN4(n3019), .IN5(n3180), .Q(\fpu_div_frac_dp/i_div_norm_inv/N30 ) );
  OA22X1 U2993 ( .IN1(\fpu_div_frac_dp/n406 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n461 ), .IN4(n3022), .Q(n3180) );
  NOR2X0 U2994 ( .IN1(n3023), .IN2(n1692), .QN(n3179) );
  OA221X1 U2995 ( .IN1(n3034), .IN2(\fpu_div_frac_dp/n432 ), .IN3(
        \fpu_div_frac_dp/n487 ), .IN4(n3019), .IN5(n3181), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N3 ) );
  OA221X1 U2996 ( .IN1(n3182), .IN2(n3018), .IN3(\fpu_div_frac_dp/n461 ), 
        .IN4(n3019), .IN5(n3183), .Q(\fpu_div_frac_dp/i_div_norm_inv/N29 ) );
  OA22X1 U2997 ( .IN1(\fpu_div_frac_dp/n407 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n462 ), .IN4(n3022), .Q(n3183) );
  NOR2X0 U2998 ( .IN1(n3023), .IN2(n1693), .QN(n3182) );
  OA221X1 U2999 ( .IN1(n3184), .IN2(n3018), .IN3(\fpu_div_frac_dp/n462 ), 
        .IN4(n3019), .IN5(n3185), .Q(\fpu_div_frac_dp/i_div_norm_inv/N28 ) );
  OA22X1 U3000 ( .IN1(\fpu_div_frac_dp/n408 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n463 ), .IN4(n3022), .Q(n3185) );
  NOR2X0 U3001 ( .IN1(n3023), .IN2(n1694), .QN(n3184) );
  OA221X1 U3002 ( .IN1(n3186), .IN2(n3018), .IN3(\fpu_div_frac_dp/n463 ), 
        .IN4(n3019), .IN5(n3187), .Q(\fpu_div_frac_dp/i_div_norm_inv/N27 ) );
  OA22X1 U3003 ( .IN1(\fpu_div_frac_dp/n409 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n464 ), .IN4(n3022), .Q(n3187) );
  NOR2X0 U3004 ( .IN1(n3023), .IN2(n1695), .QN(n3186) );
  OA221X1 U3005 ( .IN1(n3188), .IN2(n3018), .IN3(\fpu_div_frac_dp/n464 ), 
        .IN4(n3019), .IN5(n3189), .Q(\fpu_div_frac_dp/i_div_norm_inv/N26 ) );
  OA22X1 U3006 ( .IN1(\fpu_div_frac_dp/n410 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n465 ), .IN4(n3022), .Q(n3189) );
  NOR2X0 U3007 ( .IN1(n3023), .IN2(n1696), .QN(n3188) );
  OA221X1 U3008 ( .IN1(n3190), .IN2(n3018), .IN3(\fpu_div_frac_dp/n465 ), 
        .IN4(n3019), .IN5(n3191), .Q(\fpu_div_frac_dp/i_div_norm_inv/N25 ) );
  OA22X1 U3009 ( .IN1(\fpu_div_frac_dp/n411 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n466 ), .IN4(n3022), .Q(n3191) );
  NOR2X0 U3010 ( .IN1(n3023), .IN2(n1697), .QN(n3190) );
  OA221X1 U3011 ( .IN1(n3192), .IN2(n3018), .IN3(\fpu_div_frac_dp/n466 ), 
        .IN4(n3019), .IN5(n3193), .Q(\fpu_div_frac_dp/i_div_norm_inv/N24 ) );
  OA22X1 U3012 ( .IN1(\fpu_div_frac_dp/n412 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n467 ), .IN4(n3022), .Q(n3193) );
  NOR2X0 U3013 ( .IN1(n3023), .IN2(n1698), .QN(n3192) );
  OA221X1 U3014 ( .IN1(n3194), .IN2(n3018), .IN3(\fpu_div_frac_dp/n467 ), 
        .IN4(n3019), .IN5(n3195), .Q(\fpu_div_frac_dp/i_div_norm_inv/N23 ) );
  OA22X1 U3015 ( .IN1(\fpu_div_frac_dp/n413 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n468 ), .IN4(n3022), .Q(n3195) );
  NOR2X0 U3016 ( .IN1(n3023), .IN2(n1699), .QN(n3194) );
  OA221X1 U3017 ( .IN1(n3196), .IN2(n3018), .IN3(\fpu_div_frac_dp/n468 ), 
        .IN4(n3019), .IN5(n3197), .Q(\fpu_div_frac_dp/i_div_norm_inv/N22 ) );
  OA22X1 U3018 ( .IN1(\fpu_div_frac_dp/n414 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n469 ), .IN4(n3022), .Q(n3197) );
  NOR2X0 U3019 ( .IN1(n3023), .IN2(n1700), .QN(n3196) );
  OA221X1 U3020 ( .IN1(n3198), .IN2(n3018), .IN3(\fpu_div_frac_dp/n469 ), 
        .IN4(n3019), .IN5(n3199), .Q(\fpu_div_frac_dp/i_div_norm_inv/N21 ) );
  OA22X1 U3021 ( .IN1(\fpu_div_frac_dp/n415 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n470 ), .IN4(n3022), .Q(n3199) );
  NOR2X0 U3022 ( .IN1(n3023), .IN2(n1701), .QN(n3198) );
  OA221X1 U3023 ( .IN1(n3200), .IN2(n3018), .IN3(\fpu_div_frac_dp/n470 ), 
        .IN4(n3019), .IN5(n3201), .Q(\fpu_div_frac_dp/i_div_norm_inv/N20 ) );
  OA22X1 U3024 ( .IN1(\fpu_div_frac_dp/n416 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n471 ), .IN4(n3022), .Q(n3201) );
  NOR2X0 U3025 ( .IN1(n3023), .IN2(n1702), .QN(n3200) );
  OA221X1 U3026 ( .IN1(n3202), .IN2(n3018), .IN3(\fpu_div_frac_dp/n471 ), 
        .IN4(n3019), .IN5(n3203), .Q(\fpu_div_frac_dp/i_div_norm_inv/N19 ) );
  OA22X1 U3027 ( .IN1(\fpu_div_frac_dp/n417 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n472 ), .IN4(n3022), .Q(n3203) );
  NOR2X0 U3028 ( .IN1(n3023), .IN2(n1703), .QN(n3202) );
  OA221X1 U3029 ( .IN1(n3204), .IN2(n3018), .IN3(\fpu_div_frac_dp/n472 ), 
        .IN4(n3019), .IN5(n3205), .Q(\fpu_div_frac_dp/i_div_norm_inv/N18 ) );
  OA22X1 U3030 ( .IN1(\fpu_div_frac_dp/n418 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n473 ), .IN4(n3022), .Q(n3205) );
  NOR2X0 U3031 ( .IN1(n3023), .IN2(n1704), .QN(n3204) );
  OA221X1 U3032 ( .IN1(n3206), .IN2(n3018), .IN3(\fpu_div_frac_dp/n473 ), 
        .IN4(n3019), .IN5(n3207), .Q(\fpu_div_frac_dp/i_div_norm_inv/N17 ) );
  OA22X1 U3033 ( .IN1(\fpu_div_frac_dp/n419 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n474 ), .IN4(n3022), .Q(n3207) );
  NOR2X0 U3034 ( .IN1(n3023), .IN2(n1705), .QN(n3206) );
  OA221X1 U3035 ( .IN1(n3208), .IN2(n3018), .IN3(\fpu_div_frac_dp/n474 ), 
        .IN4(n3019), .IN5(n3209), .Q(\fpu_div_frac_dp/i_div_norm_inv/N16 ) );
  OA22X1 U3036 ( .IN1(\fpu_div_frac_dp/n420 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n475 ), .IN4(n3022), .Q(n3209) );
  NOR2X0 U3037 ( .IN1(n3023), .IN2(n1706), .QN(n3208) );
  OA221X1 U3038 ( .IN1(n3210), .IN2(n3018), .IN3(\fpu_div_frac_dp/n475 ), 
        .IN4(n3019), .IN5(n3211), .Q(\fpu_div_frac_dp/i_div_norm_inv/N15 ) );
  OA22X1 U3039 ( .IN1(\fpu_div_frac_dp/n421 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n476 ), .IN4(n3022), .Q(n3211) );
  NOR2X0 U3040 ( .IN1(n3023), .IN2(n1707), .QN(n3210) );
  OA221X1 U3041 ( .IN1(n3212), .IN2(n3018), .IN3(\fpu_div_frac_dp/n476 ), 
        .IN4(n3019), .IN5(n3213), .Q(\fpu_div_frac_dp/i_div_norm_inv/N14 ) );
  OA22X1 U3042 ( .IN1(\fpu_div_frac_dp/n422 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n477 ), .IN4(n3022), .Q(n3213) );
  NOR2X0 U3043 ( .IN1(n3023), .IN2(n1708), .QN(n3212) );
  AND3X1 U3044 ( .IN1(n3181), .IN2(n3214), .IN3(n3215), .Q(
        \fpu_div_frac_dp/i_div_norm_inv/N13 ) );
  OA222X1 U3045 ( .IN1(\fpu_div_frac_dp/n477 ), .IN2(n3019), .IN3(
        \fpu_div_frac_dp/n422 ), .IN4(n3034), .IN5(\fpu_div_frac_dp/n478 ), 
        .IN6(n3022), .Q(n3215) );
  INVX0 U3046 ( .INP(n3216), .ZN(n3034) );
  NAND2X0 U3047 ( .IN1(n3167), .IN2(n1639), .QN(n3214) );
  INVX0 U3048 ( .INP(n3021), .ZN(n3167) );
  OA221X1 U3049 ( .IN1(n3217), .IN2(n3018), .IN3(\fpu_div_frac_dp/n478 ), 
        .IN4(n3019), .IN5(n3218), .Q(\fpu_div_frac_dp/i_div_norm_inv/N12 ) );
  OA22X1 U3050 ( .IN1(\fpu_div_frac_dp/n424 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n479 ), .IN4(n3022), .Q(n3218) );
  NOR2X0 U3051 ( .IN1(n3023), .IN2(n1639), .QN(n3217) );
  OA221X1 U3052 ( .IN1(n3219), .IN2(n3018), .IN3(\fpu_div_frac_dp/n479 ), 
        .IN4(n3019), .IN5(n3220), .Q(\fpu_div_frac_dp/i_div_norm_inv/N11 ) );
  OA22X1 U3053 ( .IN1(\fpu_div_frac_dp/n425 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n480 ), .IN4(n3022), .Q(n3220) );
  NOR2X0 U3054 ( .IN1(n3023), .IN2(n1709), .QN(n3219) );
  OA221X1 U3055 ( .IN1(n3221), .IN2(n3018), .IN3(\fpu_div_frac_dp/n480 ), 
        .IN4(n3019), .IN5(n3222), .Q(\fpu_div_frac_dp/i_div_norm_inv/N10 ) );
  OA22X1 U3056 ( .IN1(\fpu_div_frac_dp/n426 ), .IN2(n3021), .IN3(
        \fpu_div_frac_dp/n481 ), .IN4(n3022), .Q(n3222) );
  NAND4X0 U3057 ( .IN1(n3164), .IN2(n604), .IN3(n3223), .IN4(n351), .QN(n3022)
         );
  NOR2X0 U3058 ( .IN1(n520), .IN2(n3052), .QN(n3223) );
  INVX0 U3059 ( .INP(n373), .ZN(n3052) );
  NAND2X0 U3060 ( .IN1(n3163), .IN2(\fpu_div_ctl/d2stg_denorm_dbl_in2 ), .QN(
        n3021) );
  NAND4X0 U3061 ( .IN1(n3164), .IN2(n3224), .IN3(n3225), .IN4(n373), .QN(n3019) );
  NOR2X0 U3062 ( .IN1(n604), .IN2(n520), .QN(n3225) );
  AOI21X1 U3063 ( .IN1(n3226), .IN2(n3227), .IN3(n2187), .QN(n3164) );
  NAND4X0 U3064 ( .IN1(n3228), .IN2(n3041), .IN3(n1356), .IN4(n253), .QN(n3227) );
  NOR2X0 U3065 ( .IN1(n3216), .IN2(n3023), .QN(n3018) );
  AO22X1 U3066 ( .IN1(n3163), .IN2(\fpu_div_ctl/d2stg_norm_dbl_in2 ), .IN3(
        n3229), .IN4(n3172), .Q(n3216) );
  NAND2X0 U3067 ( .IN1(n373), .IN2(n3224), .QN(n3229) );
  OR2X1 U3068 ( .IN1(n3051), .IN2(n351), .Q(n3224) );
  NAND3X0 U3069 ( .IN1(n1375), .IN2(n1651), .IN3(n585), .QN(n351) );
  INVX0 U3070 ( .INP(n3230), .ZN(n3051) );
  NAND4X0 U3071 ( .IN1(n624), .IN2(n585), .IN3(n1375), .IN4(n1682), .QN(n373)
         );
  INVX0 U3072 ( .INP(n2188), .ZN(n3163) );
  NAND2X0 U3073 ( .IN1(n619), .IN2(n3040), .QN(n2188) );
  AND2X1 U3074 ( .IN1(n86), .IN2(n36), .Q(n3040) );
  NOR2X0 U3075 ( .IN1(n3023), .IN2(n1710), .QN(n3221) );
  INVX0 U3076 ( .INP(n3181), .ZN(n3023) );
  OA21X1 U3077 ( .IN1(n3176), .IN2(n25), .IN3(n1047), .Q(n3181) );
  NAND2X0 U3078 ( .IN1(n3231), .IN2(n3172), .QN(n3176) );
  INVX0 U3079 ( .INP(n2187), .ZN(n3172) );
  OAI22X1 U3080 ( .IN1(n1356), .IN2(n253), .IN3(n3228), .IN4(n3041), .QN(n3231) );
  INVX0 U3081 ( .INP(n2131), .ZN(\fpu_div_frac_dp/d1stg_step ) );
  NAND4X0 U3082 ( .IN1(n127), .IN2(n125), .IN3(n149), .IN4(n117), .QN(n2131)
         );
  NAND2X0 U3083 ( .IN1(fdiv_clken_l), .IN2(n1047), .QN(
        \fpu_div_frac_dp/ckbuf_div_frac_dp/N1 ) );
  NAND2X0 U3084 ( .IN1(fdiv_clken_l_div_exp_buf1), .IN2(n1047), .QN(
        \fpu_div_exp_dp/ckbuf_div_exp_dp/N1 ) );
  OR4X1 U3085 ( .IN1(n3232), .IN2(\fpu_div_ctl/i_d2stg_opdec/N11 ), .IN3(
        \fpu_div_ctl/i_d3stg_opdec/N11 ), .IN4(\fpu_div_ctl/i_d4stg_opdec/N11 ), .Q(\fpu_div_ctl/i_div_pipe_active/N7 ) );
  AND2X1 U3086 ( .IN1(n1354), .IN2(n3233), .Q(n3232) );
  NAND3X0 U3087 ( .IN1(n2559), .IN2(n2060), .IN3(n196), .QN(n3233) );
  NOR2X0 U3088 ( .IN1(n1373), .IN2(n1393), .QN(n2060) );
  NOR2X0 U3089 ( .IN1(n1433), .IN2(n1552), .QN(n2559) );
  OR2X1 U3090 ( .IN1(\fpu_div_ctl/i_d7stg_opdec/N11 ), .IN2(
        \fpu_div_ctl/i_d6stg_opdec/N11 ), .Q(
        \fpu_div_ctl/i_div_expadd2_in1_exp_out/N7 ) );
  AND2X1 U3091 ( .IN1(n512), .IN2(n3234), .Q(
        \fpu_div_ctl/i_div_expadd1_in1_sng/N3 ) );
  AO21X1 U3092 ( .IN1(n1956), .IN2(\fpu_div_ctl/d1stg_sngopa[4] ), .IN3(n1957), 
        .Q(n512) );
  AND2X1 U3093 ( .IN1(inq_op[0]), .IN2(n1959), .Q(n1957) );
  AND2X1 U3094 ( .IN1(n506), .IN2(n3234), .Q(
        \fpu_div_ctl/i_div_expadd1_in1_dbl/N3 ) );
  AO21X1 U3095 ( .IN1(n1956), .IN2(\fpu_div_ctl/d1stg_dblopa[4] ), .IN3(n1958), 
        .Q(n506) );
  AND2X1 U3096 ( .IN1(inq_op[1]), .IN2(n1959), .Q(n1958) );
  NOR2X0 U3097 ( .IN1(n3235), .IN2(se), .QN(n1959) );
  NOR2X0 U3098 ( .IN1(n3236), .IN2(se), .QN(n1956) );
  NOR2X0 U3099 ( .IN1(n192), .IN2(n1999), .QN(\fpu_div_ctl/i_d7stg_opdec/N9 )
         );
  NOR2X0 U3100 ( .IN1(n1999), .IN2(n193), .QN(\fpu_div_ctl/i_d7stg_opdec/N11 )
         );
  NOR2X0 U3101 ( .IN1(n611), .IN2(n3237), .QN(\fpu_div_ctl/i_d6stg_opdec/N9 )
         );
  NOR2X0 U3102 ( .IN1(n3237), .IN2(n191), .QN(\fpu_div_ctl/i_d6stg_opdec/N11 )
         );
  NOR2X0 U3103 ( .IN1(n581), .IN2(n3237), .QN(\fpu_div_ctl/i_d6stg_opdec/N10 )
         );
  NAND2X0 U3104 ( .IN1(n1354), .IN2(n2190), .QN(n3237) );
  NAND2X0 U3105 ( .IN1(n3238), .IN2(n3239), .QN(n2190) );
  NAND3X0 U3106 ( .IN1(n3240), .IN2(n1541), .IN3(n3241), .QN(n3239) );
  MUX21X1 U3107 ( .IN1(n3242), .IN2(n3243), .S(n1395), .Q(n3241) );
  NOR2X0 U3108 ( .IN1(n581), .IN2(n1545), .QN(n3243) );
  NOR2X0 U3109 ( .IN1(n611), .IN2(n594), .QN(n3242) );
  MUX21X1 U3110 ( .IN1(n3244), .IN2(n3245), .S(n616), .Q(n3240) );
  NOR2X0 U3111 ( .IN1(n620), .IN2(n612), .QN(n3245) );
  NOR2X0 U3112 ( .IN1(n1372), .IN2(n1542), .QN(n3244) );
  AO22X1 U3113 ( .IN1(n2000), .IN2(n3246), .IN3(n607), .IN4(n3247), .Q(n3238)
         );
  NAND3X0 U3114 ( .IN1(n3248), .IN2(n1373), .IN3(n3249), .QN(n3246) );
  INVX0 U3115 ( .INP(n3247), .ZN(n3249) );
  NAND4X0 U3116 ( .IN1(n607), .IN2(n3250), .IN3(n3251), .IN4(n3252), .QN(n3247) );
  NOR4X0 U3117 ( .IN1(n3253), .IN2(n3254), .IN3(n3255), .IN4(n3256), .QN(n3252) );
  XOR2X1 U3118 ( .IN1(n616), .IN2(n605), .Q(n3256) );
  XNOR2X1 U3119 ( .IN1(n1542), .IN2(n596), .Q(n3255) );
  XNOR2X1 U3120 ( .IN1(n1575), .IN2(n594), .Q(n3254) );
  XNOR2X1 U3121 ( .IN1(n1541), .IN2(n592), .Q(n3253) );
  NOR2X0 U3122 ( .IN1(n3257), .IN2(n3258), .QN(n3251) );
  XNOR2X1 U3123 ( .IN1(n1545), .IN2(n590), .Q(n3258) );
  XNOR2X1 U3124 ( .IN1(n610), .IN2(n1395), .Q(n3257) );
  INVX0 U3125 ( .INP(n2094), .ZN(n3250) );
  NAND4X0 U3126 ( .IN1(n33), .IN2(n32), .IN3(n34), .IN4(n3259), .QN(n2094) );
  AND3X1 U3127 ( .IN1(n30), .IN2(n29), .IN3(n31), .Q(n3259) );
  NAND4X0 U3128 ( .IN1(n3260), .IN2(n605), .IN3(n3261), .IN4(n596), .QN(n3248)
         );
  NOR2X0 U3129 ( .IN1(n1409), .IN2(n1575), .QN(n3261) );
  INVX0 U3130 ( .INP(n2092), .ZN(n3260) );
  NAND2X0 U3131 ( .IN1(n590), .IN2(n610), .QN(n2092) );
  NOR2X0 U3132 ( .IN1(n1999), .IN2(n184), .QN(\fpu_div_ctl/i_d4stg_opdec/N11 )
         );
  NOR2X0 U3133 ( .IN1(n181), .IN2(n1999), .QN(\fpu_div_ctl/i_d3stg_opdec/N9 )
         );
  NOR2X0 U3134 ( .IN1(n1999), .IN2(n1549), .QN(\fpu_div_ctl/i_d3stg_opdec/N11 ) );
  NOR2X0 U3135 ( .IN1(n182), .IN2(n1999), .QN(\fpu_div_ctl/i_d3stg_opdec/N10 )
         );
  AOI21X1 U3136 ( .IN1(n3048), .IN2(n3230), .IN3(se), .QN(
        \fpu_div_ctl/i_d2stg_snan_in1/N3 ) );
  NAND4X0 U3137 ( .IN1(n628), .IN2(n591), .IN3(n1375), .IN4(n1489), .QN(n3230)
         );
  NAND4X0 U3138 ( .IN1(n591), .IN2(n627), .IN3(n1376), .IN4(n1490), .QN(n3048)
         );
  NOR3X0 U3139 ( .IN1(n1543), .IN2(se), .IN3(n3262), .QN(
        \fpu_div_ctl/i_d2stg_qnan_in1/N3 ) );
  OA22X1 U3140 ( .IN1(n627), .IN2(n47), .IN3(n628), .IN4(n54), .Q(n3262) );
  NOR2X0 U3141 ( .IN1(n1999), .IN2(n2187), .QN(\fpu_div_ctl/i_d2stg_opdec/N11 ) );
  INVX0 U3142 ( .INP(n1354), .ZN(n1999) );
  NOR3X0 U3143 ( .IN1(n50), .IN2(se), .IN3(n606), .QN(
        \fpu_div_ctl/i_d2stg_norm_sng_in2/N3 ) );
  NOR3X0 U3144 ( .IN1(n520), .IN2(se), .IN3(n606), .QN(
        \fpu_div_ctl/i_d2stg_norm_dbl_in2/N3 ) );
  NOR2X0 U3145 ( .IN1(se), .IN2(n3263), .QN(\fpu_div_ctl/i_d2stg_nan_in2/N3 )
         );
  NOR2X0 U3146 ( .IN1(se), .IN2(n3226), .QN(\fpu_div_ctl/i_d2stg_nan_in/N3 )
         );
  OA21X1 U3147 ( .IN1(n3264), .IN2(n1543), .IN3(n3263), .Q(n3226) );
  NAND2X0 U3148 ( .IN1(n585), .IN2(n3265), .QN(n3263) );
  AO22X1 U3149 ( .IN1(n1547), .IN2(n3266), .IN3(n1401), .IN4(n3267), .Q(n3265)
         );
  NAND2X0 U3150 ( .IN1(n1353), .IN2(n621), .QN(n3267) );
  NAND2X0 U3151 ( .IN1(n96), .IN2(n624), .QN(n3266) );
  OA22X1 U3152 ( .IN1(n3268), .IN2(n600), .IN3(n3269), .IN4(n615), .Q(n3264)
         );
  NOR2X0 U3153 ( .IN1(n1672), .IN2(n1489), .QN(n3269) );
  NOR2X0 U3154 ( .IN1(n1648), .IN2(n1490), .QN(n3268) );
  AND3X1 U3155 ( .IN1(n606), .IN2(n1047), .IN3(n1643), .Q(
        \fpu_div_ctl/i_d2stg_denorm_sng_in2/N3 ) );
  AND3X1 U3156 ( .IN1(n606), .IN2(n1047), .IN3(n1720), .Q(
        \fpu_div_ctl/i_d2stg_denorm_dbl_in2/N3 ) );
  NOR2X0 U3157 ( .IN1(n3270), .IN2(n1356), .QN(
        \fpu_div_ctl/i_d2stg_2zero_in/N3 ) );
  NAND3X0 U3158 ( .IN1(n627), .IN2(n604), .IN3(n88), .QN(n1356) );
  INVX0 U3159 ( .INP(\fpu_div_ctl/i_d2stg_zero_in2/N3 ), .ZN(n3270) );
  NOR2X0 U3160 ( .IN1(n253), .IN2(se), .QN(\fpu_div_ctl/i_d2stg_zero_in2/N3 )
         );
  NAND3X0 U3161 ( .IN1(n621), .IN2(n606), .IN3(n95), .QN(n253) );
  NOR2X0 U3162 ( .IN1(n3271), .IN2(n3228), .QN(
        \fpu_div_ctl/i_d2stg_2inf_in/N3 ) );
  AO21X1 U3163 ( .IN1(n3272), .IN2(n3273), .IN3(n1647), .Q(n3228) );
  NAND3X0 U3164 ( .IN1(n621), .IN2(n1401), .IN3(n1353), .QN(n3273) );
  NAND3X0 U3165 ( .IN1(n624), .IN2(n1547), .IN3(n96), .QN(n3272) );
  INVX0 U3166 ( .INP(\fpu_div_ctl/i_d2stg_inf_in1/N3 ), .ZN(n3271) );
  NOR2X0 U3167 ( .IN1(n3041), .IN2(se), .QN(\fpu_div_ctl/i_d2stg_inf_in1/N3 )
         );
  AO21X1 U3168 ( .IN1(n3274), .IN2(n3275), .IN3(n1543), .Q(n3041) );
  NAND3X0 U3169 ( .IN1(n627), .IN2(n1401), .IN3(n90), .QN(n3275) );
  NAND3X0 U3170 ( .IN1(n628), .IN2(n1547), .IN3(n89), .QN(n3274) );
  NOR2X0 U3171 ( .IN1(se), .IN2(n3234), .QN(\fpu_div_ctl/i_d234stg_fdiv/N7 )
         );
  NAND2X0 U3172 ( .IN1(n1781), .IN2(n3276), .QN(n3234) );
  NAND3X0 U3173 ( .IN1(n184), .IN2(n1549), .IN3(n2187), .QN(n3276) );
  NOR2X0 U3174 ( .IN1(n354), .IN2(n355), .QN(n2187) );
  NOR3X0 U3175 ( .IN1(n3277), .IN2(n148), .IN3(n1784), .QN(n355) );
  NOR3X0 U3176 ( .IN1(n3277), .IN2(n177), .IN3(n1785), .QN(n354) );
  NAND4X0 U3177 ( .IN1(n144), .IN2(n141), .IN3(n179), .IN4(n3278), .QN(n3277)
         );
  NOR3X0 U3178 ( .IN1(n142), .IN2(n146), .IN3(n145), .QN(n3278) );
  AND2X1 U3179 ( .IN1(inq_op[7]), .IN2(\fpu_div_ctl/i_d1stg_div/N7 ), .Q(
        \fpu_div_ctl/i_d1stg_op/N21 ) );
  AND2X1 U3180 ( .IN1(inq_op[6]), .IN2(\fpu_div_ctl/i_d1stg_div/N7 ), .Q(
        \fpu_div_ctl/i_d1stg_op/N20 ) );
  AND2X1 U3181 ( .IN1(inq_op[5]), .IN2(\fpu_div_ctl/i_d1stg_div/N7 ), .Q(
        \fpu_div_ctl/i_d1stg_op/N19 ) );
  AND2X1 U3182 ( .IN1(inq_op[4]), .IN2(\fpu_div_ctl/i_d1stg_div/N7 ), .Q(
        \fpu_div_ctl/i_d1stg_op/N18 ) );
  AND2X1 U3183 ( .IN1(inq_op[3]), .IN2(\fpu_div_ctl/i_d1stg_div/N7 ), .Q(
        \fpu_div_ctl/i_d1stg_op/N17 ) );
  AND2X1 U3184 ( .IN1(inq_op[2]), .IN2(\fpu_div_ctl/i_d1stg_div/N7 ), .Q(
        \fpu_div_ctl/i_d1stg_op/N16 ) );
  AND2X1 U3185 ( .IN1(inq_op[1]), .IN2(\fpu_div_ctl/i_d1stg_div/N7 ), .Q(
        \fpu_div_ctl/i_d1stg_op/N15 ) );
  AND2X1 U3186 ( .IN1(inq_op[0]), .IN2(\fpu_div_ctl/i_d1stg_div/N7 ), .Q(
        \fpu_div_ctl/i_d1stg_op/N14 ) );
  AND3X1 U3187 ( .IN1(n3236), .IN2(n1354), .IN3(inq_div), .Q(
        \fpu_div_ctl/i_d1stg_div/N7 ) );
  NOR2X0 U3188 ( .IN1(n152), .IN2(se), .QN(n1354) );
  INVX0 U3189 ( .INP(n3235), .ZN(n3236) );
  NAND4X0 U3190 ( .IN1(n150), .IN2(n149), .IN3(n126), .IN4(n117), .QN(n3235)
         );
  AND2X1 U3191 ( .IN1(grst_l), .IN2(n1047), .Q(\fpu_div_ctl/dffrl_div_ctl/N4 )
         );
  INVX0 U3192 ( .INP(se), .ZN(n1047) );
  AO22X1 U3193 ( .IN1(n2042), .IN2(\fpu_div_ctl/div_id_out[9] ), .IN3(n3279), 
        .IN4(n3280), .Q(div_id_out_in[9]) );
  AO22X1 U3194 ( .IN1(n2042), .IN2(\fpu_div_ctl/div_id_out[8] ), .IN3(n3279), 
        .IN4(n3281), .Q(div_id_out_in[8]) );
  NOR2X0 U3195 ( .IN1(n597), .IN2(n1351), .QN(n3279) );
  AO22X1 U3196 ( .IN1(n2042), .IN2(\fpu_div_ctl/div_id_out[7] ), .IN3(n3282), 
        .IN4(n1351), .Q(div_id_out_in[7]) );
  NOR2X0 U3197 ( .IN1(n597), .IN2(n3283), .QN(n3282) );
  AO22X1 U3198 ( .IN1(n2042), .IN2(\fpu_div_ctl/div_id_out[6] ), .IN3(n3284), 
        .IN4(n1351), .Q(div_id_out_in[6]) );
  NOR2X0 U3199 ( .IN1(n597), .IN2(n3285), .QN(n3284) );
  AO22X1 U3200 ( .IN1(n2042), .IN2(\fpu_div_ctl/div_id_out[5] ), .IN3(n3286), 
        .IN4(n597), .Q(div_id_out_in[5]) );
  NOR2X0 U3201 ( .IN1(n1351), .IN2(n3283), .QN(n3286) );
  AO22X1 U3202 ( .IN1(n2042), .IN2(\fpu_div_ctl/div_id_out[4] ), .IN3(n3287), 
        .IN4(n597), .Q(div_id_out_in[4]) );
  NOR2X0 U3203 ( .IN1(n1351), .IN2(n3285), .QN(n3287) );
  AO22X1 U3204 ( .IN1(n2042), .IN2(\fpu_div_ctl/div_id_out[3] ), .IN3(n3288), 
        .IN4(n597), .Q(div_id_out_in[3]) );
  NOR2X0 U3205 ( .IN1(n3283), .IN2(n1551), .QN(n3288) );
  INVX0 U3206 ( .INP(n3280), .ZN(n3283) );
  NOR2X0 U3207 ( .IN1(n2042), .IN2(n608), .QN(n3280) );
  AO22X1 U3208 ( .IN1(n2042), .IN2(\fpu_div_ctl/div_id_out[2] ), .IN3(n3289), 
        .IN4(n597), .Q(div_id_out_in[2]) );
  NOR2X0 U3209 ( .IN1(n3285), .IN2(n1551), .QN(n3289) );
  INVX0 U3210 ( .INP(n3281), .ZN(n3285) );
  NOR2X0 U3211 ( .IN1(n1715), .IN2(n2042), .QN(n3281) );
  MUX21X1 U3212 ( .IN1(n1722), .IN2(\fpu_div_ctl/div_id_out[1] ), .S(n2042), 
        .Q(div_id_out_in[1]) );
  MUX21X1 U3213 ( .IN1(n1723), .IN2(\fpu_div_ctl/div_id_out[0] ), .S(n2042), 
        .Q(div_id_out_in[0]) );
  NAND4X0 U3214 ( .IN1(n616), .IN2(n612), .IN3(n620), .IN4(n3290), .QN(n2042)
         );
  NOR4X0 U3215 ( .IN1(n2000), .IN2(n1395), .IN3(n1372), .IN4(n1541), .QN(n3290) );
  INVX0 U3216 ( .INP(n2854), .ZN(n2000) );
  NOR2X0 U3217 ( .IN1(n2033), .IN2(n191), .QN(n2854) );
  INVX0 U3218 ( .INP(n3291), .ZN(div_exc_out[3]) );
  NAND2X0 U3219 ( .IN1(n14), .IN2(n3291), .QN(div_exc_out[0]) );
  OA21X1 U3220 ( .IN1(n1783), .IN2(n2), .IN3(n19), .Q(n3291) );
  OA21X1 U3221 ( .IN1(n2033), .IN2(n1393), .IN3(n1781), .Q(d8stg_fdiv_in) );
  NOR2X0 U3222 ( .IN1(n196), .IN2(div_dest_rdy), .QN(n2033) );
endmodule

