
module fpu_rptr_groups ( inq_in1, inq_in2, inq_id, inq_op, inq_rnd_mode, 
        inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, inq_in1_53_32_neq_0, 
        inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0, 
        inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0, 
        inq_in2_exp_neq_ffs, ctu_tst_macrotest, ctu_tst_pre_grst_l, 
        ctu_tst_scan_disable, ctu_tst_scanmode, ctu_tst_short_chain, 
        global_shift_enable, grst_l, cluster_cken, se, arst_l, fpu_grst_l, 
        fmul_clken_l, fdiv_clken_l, scan_manual_6, si, so_unbuf, 
        pcx_fpio_data_px2, pcx_fpio_data_rdy_px2, fp_cpx_req_cq, 
        fp_cpx_data_ca, inq_sram_din_unbuf, inq_in1_add_buf1, inq_in1_mul_buf1, 
        inq_in1_div_buf1, inq_in2_add_buf1, inq_in2_mul_buf1, inq_in2_div_buf1, 
        inq_id_add_buf1, inq_id_mul_buf1, inq_id_div_buf1, inq_op_add_buf1, 
        inq_op_div_buf1, inq_op_mul_buf1, inq_rnd_mode_add_buf1, 
        inq_rnd_mode_div_buf1, inq_rnd_mode_mul_buf1, 
        inq_in1_50_0_neq_0_add_buf1, inq_in1_50_0_neq_0_mul_buf1, 
        inq_in1_50_0_neq_0_div_buf1, inq_in1_53_0_neq_0_add_buf1, 
        inq_in1_53_0_neq_0_mul_buf1, inq_in1_53_0_neq_0_div_buf1, 
        inq_in1_53_32_neq_0_add_buf1, inq_in1_53_32_neq_0_mul_buf1, 
        inq_in1_53_32_neq_0_div_buf1, inq_in1_exp_eq_0_add_buf1, 
        inq_in1_exp_eq_0_mul_buf1, inq_in1_exp_eq_0_div_buf1, 
        inq_in1_exp_neq_ffs_add_buf1, inq_in1_exp_neq_ffs_mul_buf1, 
        inq_in1_exp_neq_ffs_div_buf1, inq_in2_50_0_neq_0_add_buf1, 
        inq_in2_50_0_neq_0_mul_buf1, inq_in2_50_0_neq_0_div_buf1, 
        inq_in2_53_0_neq_0_add_buf1, inq_in2_53_0_neq_0_mul_buf1, 
        inq_in2_53_0_neq_0_div_buf1, inq_in2_53_32_neq_0_add_buf1, 
        inq_in2_53_32_neq_0_mul_buf1, inq_in2_53_32_neq_0_div_buf1, 
        inq_in2_exp_eq_0_add_buf1, inq_in2_exp_eq_0_mul_buf1, 
        inq_in2_exp_eq_0_div_buf1, inq_in2_exp_neq_ffs_add_buf1, 
        inq_in2_exp_neq_ffs_mul_buf1, inq_in2_exp_neq_ffs_div_buf1, 
        ctu_tst_macrotest_buf1, ctu_tst_pre_grst_l_buf1, 
        ctu_tst_scan_disable_buf1, ctu_tst_scanmode_buf1, 
        ctu_tst_short_chain_buf1, global_shift_enable_buf1, grst_l_buf1, 
        cluster_cken_buf1, se_add_exp_buf2, se_add_frac_buf2, se_out_buf2, 
        se_mul64_buf2, se_cluster_header_buf2, se_in_buf3, se_mul_buf4, 
        se_div_buf5, arst_l_div_buf2, arst_l_mul_buf2, 
        arst_l_cluster_header_buf2, arst_l_in_buf3, arst_l_out_buf3, 
        arst_l_add_buf4, fpu_grst_l_mul_buf1, fpu_grst_l_in_buf2, 
        fpu_grst_l_add_buf3, fmul_clken_l_buf1, fdiv_clken_l_div_exp_buf1, 
        fdiv_clken_l_div_frac_buf1, scan_manual_6_buf1, si_buf1, so, 
        pcx_fpio_data_px2_buf1, pcx_fpio_data_rdy_px2_buf1, fp_cpx_req_cq_buf1, 
        fp_cpx_data_ca_buf1, inq_sram_din_buf1 );
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  input [4:0] inq_id;
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [123:0] pcx_fpio_data_px2;
  input [7:0] fp_cpx_req_cq;
  input [144:0] fp_cpx_data_ca;
  input [155:0] inq_sram_din_unbuf;
  output [63:0] inq_in1_add_buf1;
  output [63:0] inq_in1_mul_buf1;
  output [63:0] inq_in1_div_buf1;
  output [63:0] inq_in2_add_buf1;
  output [63:0] inq_in2_mul_buf1;
  output [63:0] inq_in2_div_buf1;
  output [4:0] inq_id_add_buf1;
  output [4:0] inq_id_mul_buf1;
  output [4:0] inq_id_div_buf1;
  output [7:0] inq_op_add_buf1;
  output [7:0] inq_op_div_buf1;
  output [7:0] inq_op_mul_buf1;
  output [1:0] inq_rnd_mode_add_buf1;
  output [1:0] inq_rnd_mode_div_buf1;
  output [1:0] inq_rnd_mode_mul_buf1;
  output [123:0] pcx_fpio_data_px2_buf1;
  output [7:0] fp_cpx_req_cq_buf1;
  output [144:0] fp_cpx_data_ca_buf1;
  output [155:0] inq_sram_din_buf1;
  input inq_in1_50_0_neq_0, inq_in1_53_0_neq_0, inq_in1_53_32_neq_0,
         inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_50_0_neq_0,
         inq_in2_53_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0,
         inq_in2_exp_neq_ffs, ctu_tst_macrotest, ctu_tst_pre_grst_l,
         ctu_tst_scan_disable, ctu_tst_scanmode, ctu_tst_short_chain,
         global_shift_enable, grst_l, cluster_cken, se, arst_l, fpu_grst_l,
         fmul_clken_l, fdiv_clken_l, scan_manual_6, si, so_unbuf,
         pcx_fpio_data_rdy_px2;
  output inq_in1_50_0_neq_0_add_buf1, inq_in1_50_0_neq_0_mul_buf1,
         inq_in1_50_0_neq_0_div_buf1, inq_in1_53_0_neq_0_add_buf1,
         inq_in1_53_0_neq_0_mul_buf1, inq_in1_53_0_neq_0_div_buf1,
         inq_in1_53_32_neq_0_add_buf1, inq_in1_53_32_neq_0_mul_buf1,
         inq_in1_53_32_neq_0_div_buf1, inq_in1_exp_eq_0_add_buf1,
         inq_in1_exp_eq_0_mul_buf1, inq_in1_exp_eq_0_div_buf1,
         inq_in1_exp_neq_ffs_add_buf1, inq_in1_exp_neq_ffs_mul_buf1,
         inq_in1_exp_neq_ffs_div_buf1, inq_in2_50_0_neq_0_add_buf1,
         inq_in2_50_0_neq_0_mul_buf1, inq_in2_50_0_neq_0_div_buf1,
         inq_in2_53_0_neq_0_add_buf1, inq_in2_53_0_neq_0_mul_buf1,
         inq_in2_53_0_neq_0_div_buf1, inq_in2_53_32_neq_0_add_buf1,
         inq_in2_53_32_neq_0_mul_buf1, inq_in2_53_32_neq_0_div_buf1,
         inq_in2_exp_eq_0_add_buf1, inq_in2_exp_eq_0_mul_buf1,
         inq_in2_exp_eq_0_div_buf1, inq_in2_exp_neq_ffs_add_buf1,
         inq_in2_exp_neq_ffs_mul_buf1, inq_in2_exp_neq_ffs_div_buf1,
         ctu_tst_macrotest_buf1, ctu_tst_pre_grst_l_buf1,
         ctu_tst_scan_disable_buf1, ctu_tst_scanmode_buf1,
         ctu_tst_short_chain_buf1, global_shift_enable_buf1, grst_l_buf1,
         cluster_cken_buf1, se_add_exp_buf2, se_add_frac_buf2, se_out_buf2,
         se_mul64_buf2, se_cluster_header_buf2, se_in_buf3, se_mul_buf4,
         se_div_buf5, arst_l_div_buf2, arst_l_mul_buf2,
         arst_l_cluster_header_buf2, arst_l_in_buf3, arst_l_out_buf3,
         arst_l_add_buf4, fpu_grst_l_mul_buf1, fpu_grst_l_in_buf2,
         fpu_grst_l_add_buf3, fmul_clken_l_buf1, fdiv_clken_l_div_exp_buf1,
         fdiv_clken_l_div_frac_buf1, scan_manual_6_buf1, si_buf1, so,
         pcx_fpio_data_rdy_px2_buf1;
  wire   inq_in1_50_0_neq_0_div_buf1, inq_in1_53_0_neq_0_div_buf1,
         inq_in1_53_32_neq_0_div_buf1, inq_in1_exp_eq_0_div_buf1,
         inq_in1_exp_neq_ffs_div_buf1, inq_in2_50_0_neq_0_div_buf1,
         inq_in2_53_0_neq_0_div_buf1, inq_in2_53_32_neq_0_div_buf1,
         inq_in2_exp_eq_0_div_buf1, inq_in2_exp_neq_ffs_div_buf1,
         ctu_tst_macrotest_buf1, ctu_tst_pre_grst_l_buf1,
         ctu_tst_scan_disable_buf1, ctu_tst_scanmode_buf1,
         ctu_tst_short_chain_buf1, global_shift_enable_buf1, grst_l_buf1,
         cluster_cken_buf1, se_mul64_buf2, arst_l_in_buf3, fpu_grst_l_add_buf3,
         fmul_clken_l_buf1, fdiv_clken_l_div_exp_buf1, scan_manual_6_buf1,
         si_buf1, so, pcx_fpio_data_rdy_px2_buf1;
  assign inq_in1_mul_buf1[63] = inq_in1_div_buf1[63];
  assign inq_in1_add_buf1[63] = inq_in1_div_buf1[63];
  assign inq_in1_div_buf1[63] = inq_in1[63];
  assign inq_in1_mul_buf1[62] = inq_in1_div_buf1[62];
  assign inq_in1_add_buf1[62] = inq_in1_div_buf1[62];
  assign inq_in1_div_buf1[62] = inq_in1[62];
  assign inq_in1_mul_buf1[61] = inq_in1_div_buf1[61];
  assign inq_in1_add_buf1[61] = inq_in1_div_buf1[61];
  assign inq_in1_div_buf1[61] = inq_in1[61];
  assign inq_in1_mul_buf1[60] = inq_in1_div_buf1[60];
  assign inq_in1_add_buf1[60] = inq_in1_div_buf1[60];
  assign inq_in1_div_buf1[60] = inq_in1[60];
  assign inq_in1_mul_buf1[59] = inq_in1_div_buf1[59];
  assign inq_in1_add_buf1[59] = inq_in1_div_buf1[59];
  assign inq_in1_div_buf1[59] = inq_in1[59];
  assign inq_in1_mul_buf1[58] = inq_in1_div_buf1[58];
  assign inq_in1_add_buf1[58] = inq_in1_div_buf1[58];
  assign inq_in1_div_buf1[58] = inq_in1[58];
  assign inq_in1_mul_buf1[57] = inq_in1_div_buf1[57];
  assign inq_in1_add_buf1[57] = inq_in1_div_buf1[57];
  assign inq_in1_div_buf1[57] = inq_in1[57];
  assign inq_in1_mul_buf1[56] = inq_in1_div_buf1[56];
  assign inq_in1_add_buf1[56] = inq_in1_div_buf1[56];
  assign inq_in1_div_buf1[56] = inq_in1[56];
  assign inq_in1_mul_buf1[55] = inq_in1_div_buf1[55];
  assign inq_in1_add_buf1[55] = inq_in1_div_buf1[55];
  assign inq_in1_div_buf1[55] = inq_in1[55];
  assign inq_in1_mul_buf1[54] = inq_in1_div_buf1[54];
  assign inq_in1_add_buf1[54] = inq_in1_div_buf1[54];
  assign inq_in1_div_buf1[54] = inq_in1[54];
  assign inq_in1_mul_buf1[53] = inq_in1_div_buf1[53];
  assign inq_in1_add_buf1[53] = inq_in1_div_buf1[53];
  assign inq_in1_div_buf1[53] = inq_in1[53];
  assign inq_in1_mul_buf1[52] = inq_in1_div_buf1[52];
  assign inq_in1_add_buf1[52] = inq_in1_div_buf1[52];
  assign inq_in1_div_buf1[52] = inq_in1[52];
  assign inq_in1_mul_buf1[51] = inq_in1_div_buf1[51];
  assign inq_in1_add_buf1[51] = inq_in1_div_buf1[51];
  assign inq_in1_div_buf1[51] = inq_in1[51];
  assign inq_in1_mul_buf1[50] = inq_in1_div_buf1[50];
  assign inq_in1_add_buf1[50] = inq_in1_div_buf1[50];
  assign inq_in1_div_buf1[50] = inq_in1[50];
  assign inq_in1_mul_buf1[49] = inq_in1_div_buf1[49];
  assign inq_in1_add_buf1[49] = inq_in1_div_buf1[49];
  assign inq_in1_div_buf1[49] = inq_in1[49];
  assign inq_in1_mul_buf1[48] = inq_in1_div_buf1[48];
  assign inq_in1_add_buf1[48] = inq_in1_div_buf1[48];
  assign inq_in1_div_buf1[48] = inq_in1[48];
  assign inq_in1_mul_buf1[47] = inq_in1_div_buf1[47];
  assign inq_in1_add_buf1[47] = inq_in1_div_buf1[47];
  assign inq_in1_div_buf1[47] = inq_in1[47];
  assign inq_in1_mul_buf1[46] = inq_in1_div_buf1[46];
  assign inq_in1_add_buf1[46] = inq_in1_div_buf1[46];
  assign inq_in1_div_buf1[46] = inq_in1[46];
  assign inq_in1_mul_buf1[45] = inq_in1_div_buf1[45];
  assign inq_in1_add_buf1[45] = inq_in1_div_buf1[45];
  assign inq_in1_div_buf1[45] = inq_in1[45];
  assign inq_in1_mul_buf1[44] = inq_in1_div_buf1[44];
  assign inq_in1_add_buf1[44] = inq_in1_div_buf1[44];
  assign inq_in1_div_buf1[44] = inq_in1[44];
  assign inq_in1_mul_buf1[43] = inq_in1_div_buf1[43];
  assign inq_in1_add_buf1[43] = inq_in1_div_buf1[43];
  assign inq_in1_div_buf1[43] = inq_in1[43];
  assign inq_in1_mul_buf1[42] = inq_in1_div_buf1[42];
  assign inq_in1_add_buf1[42] = inq_in1_div_buf1[42];
  assign inq_in1_div_buf1[42] = inq_in1[42];
  assign inq_in1_mul_buf1[41] = inq_in1_div_buf1[41];
  assign inq_in1_add_buf1[41] = inq_in1_div_buf1[41];
  assign inq_in1_div_buf1[41] = inq_in1[41];
  assign inq_in1_mul_buf1[40] = inq_in1_div_buf1[40];
  assign inq_in1_add_buf1[40] = inq_in1_div_buf1[40];
  assign inq_in1_div_buf1[40] = inq_in1[40];
  assign inq_in1_mul_buf1[39] = inq_in1_div_buf1[39];
  assign inq_in1_add_buf1[39] = inq_in1_div_buf1[39];
  assign inq_in1_div_buf1[39] = inq_in1[39];
  assign inq_in1_mul_buf1[38] = inq_in1_div_buf1[38];
  assign inq_in1_add_buf1[38] = inq_in1_div_buf1[38];
  assign inq_in1_div_buf1[38] = inq_in1[38];
  assign inq_in1_mul_buf1[37] = inq_in1_div_buf1[37];
  assign inq_in1_add_buf1[37] = inq_in1_div_buf1[37];
  assign inq_in1_div_buf1[37] = inq_in1[37];
  assign inq_in1_mul_buf1[36] = inq_in1_div_buf1[36];
  assign inq_in1_add_buf1[36] = inq_in1_div_buf1[36];
  assign inq_in1_div_buf1[36] = inq_in1[36];
  assign inq_in1_mul_buf1[35] = inq_in1_div_buf1[35];
  assign inq_in1_add_buf1[35] = inq_in1_div_buf1[35];
  assign inq_in1_div_buf1[35] = inq_in1[35];
  assign inq_in1_mul_buf1[34] = inq_in1_div_buf1[34];
  assign inq_in1_add_buf1[34] = inq_in1_div_buf1[34];
  assign inq_in1_div_buf1[34] = inq_in1[34];
  assign inq_in1_mul_buf1[33] = inq_in1_div_buf1[33];
  assign inq_in1_add_buf1[33] = inq_in1_div_buf1[33];
  assign inq_in1_div_buf1[33] = inq_in1[33];
  assign inq_in1_mul_buf1[32] = inq_in1_div_buf1[32];
  assign inq_in1_add_buf1[32] = inq_in1_div_buf1[32];
  assign inq_in1_div_buf1[32] = inq_in1[32];
  assign inq_in1_mul_buf1[31] = inq_in1_div_buf1[31];
  assign inq_in1_add_buf1[31] = inq_in1_div_buf1[31];
  assign inq_in1_div_buf1[31] = inq_in1[31];
  assign inq_in1_mul_buf1[30] = inq_in1_div_buf1[30];
  assign inq_in1_add_buf1[30] = inq_in1_div_buf1[30];
  assign inq_in1_div_buf1[30] = inq_in1[30];
  assign inq_in1_mul_buf1[29] = inq_in1_div_buf1[29];
  assign inq_in1_add_buf1[29] = inq_in1_div_buf1[29];
  assign inq_in1_div_buf1[29] = inq_in1[29];
  assign inq_in1_mul_buf1[28] = inq_in1_div_buf1[28];
  assign inq_in1_add_buf1[28] = inq_in1_div_buf1[28];
  assign inq_in1_div_buf1[28] = inq_in1[28];
  assign inq_in1_mul_buf1[27] = inq_in1_div_buf1[27];
  assign inq_in1_add_buf1[27] = inq_in1_div_buf1[27];
  assign inq_in1_div_buf1[27] = inq_in1[27];
  assign inq_in1_mul_buf1[26] = inq_in1_div_buf1[26];
  assign inq_in1_add_buf1[26] = inq_in1_div_buf1[26];
  assign inq_in1_div_buf1[26] = inq_in1[26];
  assign inq_in1_mul_buf1[25] = inq_in1_div_buf1[25];
  assign inq_in1_add_buf1[25] = inq_in1_div_buf1[25];
  assign inq_in1_div_buf1[25] = inq_in1[25];
  assign inq_in1_mul_buf1[24] = inq_in1_div_buf1[24];
  assign inq_in1_add_buf1[24] = inq_in1_div_buf1[24];
  assign inq_in1_div_buf1[24] = inq_in1[24];
  assign inq_in1_mul_buf1[23] = inq_in1_div_buf1[23];
  assign inq_in1_add_buf1[23] = inq_in1_div_buf1[23];
  assign inq_in1_div_buf1[23] = inq_in1[23];
  assign inq_in1_mul_buf1[22] = inq_in1_div_buf1[22];
  assign inq_in1_add_buf1[22] = inq_in1_div_buf1[22];
  assign inq_in1_div_buf1[22] = inq_in1[22];
  assign inq_in1_mul_buf1[21] = inq_in1_div_buf1[21];
  assign inq_in1_add_buf1[21] = inq_in1_div_buf1[21];
  assign inq_in1_div_buf1[21] = inq_in1[21];
  assign inq_in1_mul_buf1[20] = inq_in1_div_buf1[20];
  assign inq_in1_add_buf1[20] = inq_in1_div_buf1[20];
  assign inq_in1_div_buf1[20] = inq_in1[20];
  assign inq_in1_mul_buf1[19] = inq_in1_div_buf1[19];
  assign inq_in1_add_buf1[19] = inq_in1_div_buf1[19];
  assign inq_in1_div_buf1[19] = inq_in1[19];
  assign inq_in1_mul_buf1[18] = inq_in1_div_buf1[18];
  assign inq_in1_add_buf1[18] = inq_in1_div_buf1[18];
  assign inq_in1_div_buf1[18] = inq_in1[18];
  assign inq_in1_mul_buf1[17] = inq_in1_div_buf1[17];
  assign inq_in1_add_buf1[17] = inq_in1_div_buf1[17];
  assign inq_in1_div_buf1[17] = inq_in1[17];
  assign inq_in1_mul_buf1[16] = inq_in1_div_buf1[16];
  assign inq_in1_add_buf1[16] = inq_in1_div_buf1[16];
  assign inq_in1_div_buf1[16] = inq_in1[16];
  assign inq_in1_mul_buf1[15] = inq_in1_div_buf1[15];
  assign inq_in1_add_buf1[15] = inq_in1_div_buf1[15];
  assign inq_in1_div_buf1[15] = inq_in1[15];
  assign inq_in1_mul_buf1[14] = inq_in1_div_buf1[14];
  assign inq_in1_add_buf1[14] = inq_in1_div_buf1[14];
  assign inq_in1_div_buf1[14] = inq_in1[14];
  assign inq_in1_mul_buf1[13] = inq_in1_div_buf1[13];
  assign inq_in1_add_buf1[13] = inq_in1_div_buf1[13];
  assign inq_in1_div_buf1[13] = inq_in1[13];
  assign inq_in1_mul_buf1[12] = inq_in1_div_buf1[12];
  assign inq_in1_add_buf1[12] = inq_in1_div_buf1[12];
  assign inq_in1_div_buf1[12] = inq_in1[12];
  assign inq_in1_mul_buf1[11] = inq_in1_div_buf1[11];
  assign inq_in1_add_buf1[11] = inq_in1_div_buf1[11];
  assign inq_in1_div_buf1[11] = inq_in1[11];
  assign inq_in1_mul_buf1[10] = inq_in1_div_buf1[10];
  assign inq_in1_add_buf1[10] = inq_in1_div_buf1[10];
  assign inq_in1_div_buf1[10] = inq_in1[10];
  assign inq_in1_mul_buf1[9] = inq_in1_div_buf1[9];
  assign inq_in1_add_buf1[9] = inq_in1_div_buf1[9];
  assign inq_in1_div_buf1[9] = inq_in1[9];
  assign inq_in1_mul_buf1[8] = inq_in1_div_buf1[8];
  assign inq_in1_add_buf1[8] = inq_in1_div_buf1[8];
  assign inq_in1_div_buf1[8] = inq_in1[8];
  assign inq_in1_mul_buf1[7] = inq_in1_div_buf1[7];
  assign inq_in1_add_buf1[7] = inq_in1_div_buf1[7];
  assign inq_in1_div_buf1[7] = inq_in1[7];
  assign inq_in1_mul_buf1[6] = inq_in1_div_buf1[6];
  assign inq_in1_add_buf1[6] = inq_in1_div_buf1[6];
  assign inq_in1_div_buf1[6] = inq_in1[6];
  assign inq_in1_mul_buf1[5] = inq_in1_div_buf1[5];
  assign inq_in1_add_buf1[5] = inq_in1_div_buf1[5];
  assign inq_in1_div_buf1[5] = inq_in1[5];
  assign inq_in1_mul_buf1[4] = inq_in1_div_buf1[4];
  assign inq_in1_add_buf1[4] = inq_in1_div_buf1[4];
  assign inq_in1_div_buf1[4] = inq_in1[4];
  assign inq_in1_mul_buf1[3] = inq_in1_div_buf1[3];
  assign inq_in1_add_buf1[3] = inq_in1_div_buf1[3];
  assign inq_in1_div_buf1[3] = inq_in1[3];
  assign inq_in1_mul_buf1[2] = inq_in1_div_buf1[2];
  assign inq_in1_add_buf1[2] = inq_in1_div_buf1[2];
  assign inq_in1_div_buf1[2] = inq_in1[2];
  assign inq_in1_mul_buf1[1] = inq_in1_div_buf1[1];
  assign inq_in1_add_buf1[1] = inq_in1_div_buf1[1];
  assign inq_in1_div_buf1[1] = inq_in1[1];
  assign inq_in1_mul_buf1[0] = inq_in1_div_buf1[0];
  assign inq_in1_add_buf1[0] = inq_in1_div_buf1[0];
  assign inq_in1_div_buf1[0] = inq_in1[0];
  assign inq_in2_mul_buf1[63] = inq_in2_div_buf1[63];
  assign inq_in2_add_buf1[63] = inq_in2_div_buf1[63];
  assign inq_in2_div_buf1[63] = inq_in2[63];
  assign inq_in2_mul_buf1[62] = inq_in2_div_buf1[62];
  assign inq_in2_add_buf1[62] = inq_in2_div_buf1[62];
  assign inq_in2_div_buf1[62] = inq_in2[62];
  assign inq_in2_mul_buf1[61] = inq_in2_div_buf1[61];
  assign inq_in2_add_buf1[61] = inq_in2_div_buf1[61];
  assign inq_in2_div_buf1[61] = inq_in2[61];
  assign inq_in2_mul_buf1[60] = inq_in2_div_buf1[60];
  assign inq_in2_add_buf1[60] = inq_in2_div_buf1[60];
  assign inq_in2_div_buf1[60] = inq_in2[60];
  assign inq_in2_mul_buf1[59] = inq_in2_div_buf1[59];
  assign inq_in2_add_buf1[59] = inq_in2_div_buf1[59];
  assign inq_in2_div_buf1[59] = inq_in2[59];
  assign inq_in2_mul_buf1[58] = inq_in2_div_buf1[58];
  assign inq_in2_add_buf1[58] = inq_in2_div_buf1[58];
  assign inq_in2_div_buf1[58] = inq_in2[58];
  assign inq_in2_mul_buf1[57] = inq_in2_div_buf1[57];
  assign inq_in2_add_buf1[57] = inq_in2_div_buf1[57];
  assign inq_in2_div_buf1[57] = inq_in2[57];
  assign inq_in2_mul_buf1[56] = inq_in2_div_buf1[56];
  assign inq_in2_add_buf1[56] = inq_in2_div_buf1[56];
  assign inq_in2_div_buf1[56] = inq_in2[56];
  assign inq_in2_mul_buf1[55] = inq_in2_div_buf1[55];
  assign inq_in2_add_buf1[55] = inq_in2_div_buf1[55];
  assign inq_in2_div_buf1[55] = inq_in2[55];
  assign inq_in2_mul_buf1[54] = inq_in2_div_buf1[54];
  assign inq_in2_add_buf1[54] = inq_in2_div_buf1[54];
  assign inq_in2_div_buf1[54] = inq_in2[54];
  assign inq_in2_mul_buf1[53] = inq_in2_div_buf1[53];
  assign inq_in2_add_buf1[53] = inq_in2_div_buf1[53];
  assign inq_in2_div_buf1[53] = inq_in2[53];
  assign inq_in2_mul_buf1[52] = inq_in2_div_buf1[52];
  assign inq_in2_add_buf1[52] = inq_in2_div_buf1[52];
  assign inq_in2_div_buf1[52] = inq_in2[52];
  assign inq_in2_mul_buf1[51] = inq_in2_div_buf1[51];
  assign inq_in2_add_buf1[51] = inq_in2_div_buf1[51];
  assign inq_in2_div_buf1[51] = inq_in2[51];
  assign inq_in2_mul_buf1[50] = inq_in2_div_buf1[50];
  assign inq_in2_add_buf1[50] = inq_in2_div_buf1[50];
  assign inq_in2_div_buf1[50] = inq_in2[50];
  assign inq_in2_mul_buf1[49] = inq_in2_div_buf1[49];
  assign inq_in2_add_buf1[49] = inq_in2_div_buf1[49];
  assign inq_in2_div_buf1[49] = inq_in2[49];
  assign inq_in2_mul_buf1[48] = inq_in2_div_buf1[48];
  assign inq_in2_add_buf1[48] = inq_in2_div_buf1[48];
  assign inq_in2_div_buf1[48] = inq_in2[48];
  assign inq_in2_mul_buf1[47] = inq_in2_div_buf1[47];
  assign inq_in2_add_buf1[47] = inq_in2_div_buf1[47];
  assign inq_in2_div_buf1[47] = inq_in2[47];
  assign inq_in2_mul_buf1[46] = inq_in2_div_buf1[46];
  assign inq_in2_add_buf1[46] = inq_in2_div_buf1[46];
  assign inq_in2_div_buf1[46] = inq_in2[46];
  assign inq_in2_mul_buf1[45] = inq_in2_div_buf1[45];
  assign inq_in2_add_buf1[45] = inq_in2_div_buf1[45];
  assign inq_in2_div_buf1[45] = inq_in2[45];
  assign inq_in2_mul_buf1[44] = inq_in2_div_buf1[44];
  assign inq_in2_add_buf1[44] = inq_in2_div_buf1[44];
  assign inq_in2_div_buf1[44] = inq_in2[44];
  assign inq_in2_mul_buf1[43] = inq_in2_div_buf1[43];
  assign inq_in2_add_buf1[43] = inq_in2_div_buf1[43];
  assign inq_in2_div_buf1[43] = inq_in2[43];
  assign inq_in2_mul_buf1[42] = inq_in2_div_buf1[42];
  assign inq_in2_add_buf1[42] = inq_in2_div_buf1[42];
  assign inq_in2_div_buf1[42] = inq_in2[42];
  assign inq_in2_mul_buf1[41] = inq_in2_div_buf1[41];
  assign inq_in2_add_buf1[41] = inq_in2_div_buf1[41];
  assign inq_in2_div_buf1[41] = inq_in2[41];
  assign inq_in2_mul_buf1[40] = inq_in2_div_buf1[40];
  assign inq_in2_add_buf1[40] = inq_in2_div_buf1[40];
  assign inq_in2_div_buf1[40] = inq_in2[40];
  assign inq_in2_mul_buf1[39] = inq_in2_div_buf1[39];
  assign inq_in2_add_buf1[39] = inq_in2_div_buf1[39];
  assign inq_in2_div_buf1[39] = inq_in2[39];
  assign inq_in2_mul_buf1[38] = inq_in2_div_buf1[38];
  assign inq_in2_add_buf1[38] = inq_in2_div_buf1[38];
  assign inq_in2_div_buf1[38] = inq_in2[38];
  assign inq_in2_mul_buf1[37] = inq_in2_div_buf1[37];
  assign inq_in2_add_buf1[37] = inq_in2_div_buf1[37];
  assign inq_in2_div_buf1[37] = inq_in2[37];
  assign inq_in2_mul_buf1[36] = inq_in2_div_buf1[36];
  assign inq_in2_add_buf1[36] = inq_in2_div_buf1[36];
  assign inq_in2_div_buf1[36] = inq_in2[36];
  assign inq_in2_mul_buf1[35] = inq_in2_div_buf1[35];
  assign inq_in2_add_buf1[35] = inq_in2_div_buf1[35];
  assign inq_in2_div_buf1[35] = inq_in2[35];
  assign inq_in2_mul_buf1[34] = inq_in2_div_buf1[34];
  assign inq_in2_add_buf1[34] = inq_in2_div_buf1[34];
  assign inq_in2_div_buf1[34] = inq_in2[34];
  assign inq_in2_mul_buf1[33] = inq_in2_div_buf1[33];
  assign inq_in2_add_buf1[33] = inq_in2_div_buf1[33];
  assign inq_in2_div_buf1[33] = inq_in2[33];
  assign inq_in2_mul_buf1[32] = inq_in2_div_buf1[32];
  assign inq_in2_add_buf1[32] = inq_in2_div_buf1[32];
  assign inq_in2_div_buf1[32] = inq_in2[32];
  assign inq_in2_mul_buf1[31] = inq_in2_div_buf1[31];
  assign inq_in2_add_buf1[31] = inq_in2_div_buf1[31];
  assign inq_in2_div_buf1[31] = inq_in2[31];
  assign inq_in2_mul_buf1[30] = inq_in2_div_buf1[30];
  assign inq_in2_add_buf1[30] = inq_in2_div_buf1[30];
  assign inq_in2_div_buf1[30] = inq_in2[30];
  assign inq_in2_mul_buf1[29] = inq_in2_div_buf1[29];
  assign inq_in2_add_buf1[29] = inq_in2_div_buf1[29];
  assign inq_in2_div_buf1[29] = inq_in2[29];
  assign inq_in2_mul_buf1[28] = inq_in2_div_buf1[28];
  assign inq_in2_add_buf1[28] = inq_in2_div_buf1[28];
  assign inq_in2_div_buf1[28] = inq_in2[28];
  assign inq_in2_mul_buf1[27] = inq_in2_div_buf1[27];
  assign inq_in2_add_buf1[27] = inq_in2_div_buf1[27];
  assign inq_in2_div_buf1[27] = inq_in2[27];
  assign inq_in2_mul_buf1[26] = inq_in2_div_buf1[26];
  assign inq_in2_add_buf1[26] = inq_in2_div_buf1[26];
  assign inq_in2_div_buf1[26] = inq_in2[26];
  assign inq_in2_mul_buf1[25] = inq_in2_div_buf1[25];
  assign inq_in2_add_buf1[25] = inq_in2_div_buf1[25];
  assign inq_in2_div_buf1[25] = inq_in2[25];
  assign inq_in2_mul_buf1[24] = inq_in2_div_buf1[24];
  assign inq_in2_add_buf1[24] = inq_in2_div_buf1[24];
  assign inq_in2_div_buf1[24] = inq_in2[24];
  assign inq_in2_mul_buf1[23] = inq_in2_div_buf1[23];
  assign inq_in2_add_buf1[23] = inq_in2_div_buf1[23];
  assign inq_in2_div_buf1[23] = inq_in2[23];
  assign inq_in2_mul_buf1[22] = inq_in2_div_buf1[22];
  assign inq_in2_add_buf1[22] = inq_in2_div_buf1[22];
  assign inq_in2_div_buf1[22] = inq_in2[22];
  assign inq_in2_mul_buf1[21] = inq_in2_div_buf1[21];
  assign inq_in2_add_buf1[21] = inq_in2_div_buf1[21];
  assign inq_in2_div_buf1[21] = inq_in2[21];
  assign inq_in2_mul_buf1[20] = inq_in2_div_buf1[20];
  assign inq_in2_add_buf1[20] = inq_in2_div_buf1[20];
  assign inq_in2_div_buf1[20] = inq_in2[20];
  assign inq_in2_mul_buf1[19] = inq_in2_div_buf1[19];
  assign inq_in2_add_buf1[19] = inq_in2_div_buf1[19];
  assign inq_in2_div_buf1[19] = inq_in2[19];
  assign inq_in2_mul_buf1[18] = inq_in2_div_buf1[18];
  assign inq_in2_add_buf1[18] = inq_in2_div_buf1[18];
  assign inq_in2_div_buf1[18] = inq_in2[18];
  assign inq_in2_mul_buf1[17] = inq_in2_div_buf1[17];
  assign inq_in2_add_buf1[17] = inq_in2_div_buf1[17];
  assign inq_in2_div_buf1[17] = inq_in2[17];
  assign inq_in2_mul_buf1[16] = inq_in2_div_buf1[16];
  assign inq_in2_add_buf1[16] = inq_in2_div_buf1[16];
  assign inq_in2_div_buf1[16] = inq_in2[16];
  assign inq_in2_mul_buf1[15] = inq_in2_div_buf1[15];
  assign inq_in2_add_buf1[15] = inq_in2_div_buf1[15];
  assign inq_in2_div_buf1[15] = inq_in2[15];
  assign inq_in2_mul_buf1[14] = inq_in2_div_buf1[14];
  assign inq_in2_add_buf1[14] = inq_in2_div_buf1[14];
  assign inq_in2_div_buf1[14] = inq_in2[14];
  assign inq_in2_mul_buf1[13] = inq_in2_div_buf1[13];
  assign inq_in2_add_buf1[13] = inq_in2_div_buf1[13];
  assign inq_in2_div_buf1[13] = inq_in2[13];
  assign inq_in2_mul_buf1[12] = inq_in2_div_buf1[12];
  assign inq_in2_add_buf1[12] = inq_in2_div_buf1[12];
  assign inq_in2_div_buf1[12] = inq_in2[12];
  assign inq_in2_mul_buf1[11] = inq_in2_div_buf1[11];
  assign inq_in2_add_buf1[11] = inq_in2_div_buf1[11];
  assign inq_in2_div_buf1[11] = inq_in2[11];
  assign inq_in2_mul_buf1[10] = inq_in2_div_buf1[10];
  assign inq_in2_add_buf1[10] = inq_in2_div_buf1[10];
  assign inq_in2_div_buf1[10] = inq_in2[10];
  assign inq_in2_mul_buf1[9] = inq_in2_div_buf1[9];
  assign inq_in2_add_buf1[9] = inq_in2_div_buf1[9];
  assign inq_in2_div_buf1[9] = inq_in2[9];
  assign inq_in2_mul_buf1[8] = inq_in2_div_buf1[8];
  assign inq_in2_add_buf1[8] = inq_in2_div_buf1[8];
  assign inq_in2_div_buf1[8] = inq_in2[8];
  assign inq_in2_mul_buf1[7] = inq_in2_div_buf1[7];
  assign inq_in2_add_buf1[7] = inq_in2_div_buf1[7];
  assign inq_in2_div_buf1[7] = inq_in2[7];
  assign inq_in2_mul_buf1[6] = inq_in2_div_buf1[6];
  assign inq_in2_add_buf1[6] = inq_in2_div_buf1[6];
  assign inq_in2_div_buf1[6] = inq_in2[6];
  assign inq_in2_mul_buf1[5] = inq_in2_div_buf1[5];
  assign inq_in2_add_buf1[5] = inq_in2_div_buf1[5];
  assign inq_in2_div_buf1[5] = inq_in2[5];
  assign inq_in2_mul_buf1[4] = inq_in2_div_buf1[4];
  assign inq_in2_add_buf1[4] = inq_in2_div_buf1[4];
  assign inq_in2_div_buf1[4] = inq_in2[4];
  assign inq_in2_mul_buf1[3] = inq_in2_div_buf1[3];
  assign inq_in2_add_buf1[3] = inq_in2_div_buf1[3];
  assign inq_in2_div_buf1[3] = inq_in2[3];
  assign inq_in2_mul_buf1[2] = inq_in2_div_buf1[2];
  assign inq_in2_add_buf1[2] = inq_in2_div_buf1[2];
  assign inq_in2_div_buf1[2] = inq_in2[2];
  assign inq_in2_mul_buf1[1] = inq_in2_div_buf1[1];
  assign inq_in2_add_buf1[1] = inq_in2_div_buf1[1];
  assign inq_in2_div_buf1[1] = inq_in2[1];
  assign inq_in2_mul_buf1[0] = inq_in2_div_buf1[0];
  assign inq_in2_add_buf1[0] = inq_in2_div_buf1[0];
  assign inq_in2_div_buf1[0] = inq_in2[0];
  assign inq_id_mul_buf1[4] = inq_id_div_buf1[4];
  assign inq_id_add_buf1[4] = inq_id_div_buf1[4];
  assign inq_id_div_buf1[4] = inq_id[4];
  assign inq_id_mul_buf1[3] = inq_id_div_buf1[3];
  assign inq_id_add_buf1[3] = inq_id_div_buf1[3];
  assign inq_id_div_buf1[3] = inq_id[3];
  assign inq_id_mul_buf1[2] = inq_id_div_buf1[2];
  assign inq_id_add_buf1[2] = inq_id_div_buf1[2];
  assign inq_id_div_buf1[2] = inq_id[2];
  assign inq_id_mul_buf1[1] = inq_id_div_buf1[1];
  assign inq_id_add_buf1[1] = inq_id_div_buf1[1];
  assign inq_id_div_buf1[1] = inq_id[1];
  assign inq_id_mul_buf1[0] = inq_id_div_buf1[0];
  assign inq_id_add_buf1[0] = inq_id_div_buf1[0];
  assign inq_id_div_buf1[0] = inq_id[0];
  assign inq_op_mul_buf1[7] = inq_op_div_buf1[7];
  assign inq_op_add_buf1[7] = inq_op_div_buf1[7];
  assign inq_op_div_buf1[7] = inq_op[7];
  assign inq_op_mul_buf1[6] = inq_op_div_buf1[6];
  assign inq_op_add_buf1[6] = inq_op_div_buf1[6];
  assign inq_op_div_buf1[6] = inq_op[6];
  assign inq_op_mul_buf1[5] = inq_op_div_buf1[5];
  assign inq_op_add_buf1[5] = inq_op_div_buf1[5];
  assign inq_op_div_buf1[5] = inq_op[5];
  assign inq_op_mul_buf1[4] = inq_op_div_buf1[4];
  assign inq_op_add_buf1[4] = inq_op_div_buf1[4];
  assign inq_op_div_buf1[4] = inq_op[4];
  assign inq_op_mul_buf1[3] = inq_op_div_buf1[3];
  assign inq_op_add_buf1[3] = inq_op_div_buf1[3];
  assign inq_op_div_buf1[3] = inq_op[3];
  assign inq_op_mul_buf1[2] = inq_op_div_buf1[2];
  assign inq_op_add_buf1[2] = inq_op_div_buf1[2];
  assign inq_op_div_buf1[2] = inq_op[2];
  assign inq_op_mul_buf1[1] = inq_op_div_buf1[1];
  assign inq_op_add_buf1[1] = inq_op_div_buf1[1];
  assign inq_op_div_buf1[1] = inq_op[1];
  assign inq_op_mul_buf1[0] = inq_op_div_buf1[0];
  assign inq_op_add_buf1[0] = inq_op_div_buf1[0];
  assign inq_op_div_buf1[0] = inq_op[0];
  assign inq_rnd_mode_mul_buf1[1] = inq_rnd_mode_div_buf1[1];
  assign inq_rnd_mode_add_buf1[1] = inq_rnd_mode_div_buf1[1];
  assign inq_rnd_mode_div_buf1[1] = inq_rnd_mode[1];
  assign inq_rnd_mode_mul_buf1[0] = inq_rnd_mode_div_buf1[0];
  assign inq_rnd_mode_add_buf1[0] = inq_rnd_mode_div_buf1[0];
  assign inq_rnd_mode_div_buf1[0] = inq_rnd_mode[0];
  assign inq_in1_50_0_neq_0_mul_buf1 = inq_in1_50_0_neq_0_div_buf1;
  assign inq_in1_50_0_neq_0_add_buf1 = inq_in1_50_0_neq_0_div_buf1;
  assign inq_in1_50_0_neq_0_div_buf1 = inq_in1_50_0_neq_0;
  assign inq_in1_53_0_neq_0_mul_buf1 = inq_in1_53_0_neq_0_div_buf1;
  assign inq_in1_53_0_neq_0_add_buf1 = inq_in1_53_0_neq_0_div_buf1;
  assign inq_in1_53_0_neq_0_div_buf1 = inq_in1_53_0_neq_0;
  assign inq_in1_53_32_neq_0_mul_buf1 = inq_in1_53_32_neq_0_div_buf1;
  assign inq_in1_53_32_neq_0_add_buf1 = inq_in1_53_32_neq_0_div_buf1;
  assign inq_in1_53_32_neq_0_div_buf1 = inq_in1_53_32_neq_0;
  assign inq_in1_exp_eq_0_mul_buf1 = inq_in1_exp_eq_0_div_buf1;
  assign inq_in1_exp_eq_0_add_buf1 = inq_in1_exp_eq_0_div_buf1;
  assign inq_in1_exp_eq_0_div_buf1 = inq_in1_exp_eq_0;
  assign inq_in1_exp_neq_ffs_mul_buf1 = inq_in1_exp_neq_ffs_div_buf1;
  assign inq_in1_exp_neq_ffs_add_buf1 = inq_in1_exp_neq_ffs_div_buf1;
  assign inq_in1_exp_neq_ffs_div_buf1 = inq_in1_exp_neq_ffs;
  assign inq_in2_50_0_neq_0_mul_buf1 = inq_in2_50_0_neq_0_div_buf1;
  assign inq_in2_50_0_neq_0_add_buf1 = inq_in2_50_0_neq_0_div_buf1;
  assign inq_in2_50_0_neq_0_div_buf1 = inq_in2_50_0_neq_0;
  assign inq_in2_53_0_neq_0_mul_buf1 = inq_in2_53_0_neq_0_div_buf1;
  assign inq_in2_53_0_neq_0_add_buf1 = inq_in2_53_0_neq_0_div_buf1;
  assign inq_in2_53_0_neq_0_div_buf1 = inq_in2_53_0_neq_0;
  assign inq_in2_53_32_neq_0_mul_buf1 = inq_in2_53_32_neq_0_div_buf1;
  assign inq_in2_53_32_neq_0_add_buf1 = inq_in2_53_32_neq_0_div_buf1;
  assign inq_in2_53_32_neq_0_div_buf1 = inq_in2_53_32_neq_0;
  assign inq_in2_exp_eq_0_mul_buf1 = inq_in2_exp_eq_0_div_buf1;
  assign inq_in2_exp_eq_0_add_buf1 = inq_in2_exp_eq_0_div_buf1;
  assign inq_in2_exp_eq_0_div_buf1 = inq_in2_exp_eq_0;
  assign inq_in2_exp_neq_ffs_mul_buf1 = inq_in2_exp_neq_ffs_div_buf1;
  assign inq_in2_exp_neq_ffs_add_buf1 = inq_in2_exp_neq_ffs_div_buf1;
  assign inq_in2_exp_neq_ffs_div_buf1 = inq_in2_exp_neq_ffs;
  assign ctu_tst_macrotest_buf1 = ctu_tst_macrotest;
  assign ctu_tst_pre_grst_l_buf1 = ctu_tst_pre_grst_l;
  assign ctu_tst_scan_disable_buf1 = ctu_tst_scan_disable;
  assign ctu_tst_scanmode_buf1 = ctu_tst_scanmode;
  assign ctu_tst_short_chain_buf1 = ctu_tst_short_chain;
  assign global_shift_enable_buf1 = global_shift_enable;
  assign grst_l_buf1 = grst_l;
  assign cluster_cken_buf1 = cluster_cken;
  assign se_div_buf5 = se_mul64_buf2;
  assign se_mul_buf4 = se_mul64_buf2;
  assign se_in_buf3 = se_mul64_buf2;
  assign se_cluster_header_buf2 = se_mul64_buf2;
  assign se_out_buf2 = se_mul64_buf2;
  assign se_add_frac_buf2 = se_mul64_buf2;
  assign se_add_exp_buf2 = se_mul64_buf2;
  assign se_mul64_buf2 = se;
  assign arst_l_add_buf4 = arst_l_in_buf3;
  assign arst_l_out_buf3 = arst_l_in_buf3;
  assign arst_l_cluster_header_buf2 = arst_l_in_buf3;
  assign arst_l_mul_buf2 = arst_l_in_buf3;
  assign arst_l_div_buf2 = arst_l_in_buf3;
  assign arst_l_in_buf3 = arst_l;
  assign fpu_grst_l_in_buf2 = fpu_grst_l_add_buf3;
  assign fpu_grst_l_mul_buf1 = fpu_grst_l_add_buf3;
  assign fpu_grst_l_add_buf3 = fpu_grst_l;
  assign fmul_clken_l_buf1 = fmul_clken_l;
  assign fdiv_clken_l_div_frac_buf1 = fdiv_clken_l_div_exp_buf1;
  assign fdiv_clken_l_div_exp_buf1 = fdiv_clken_l;
  assign scan_manual_6_buf1 = scan_manual_6;
  assign si_buf1 = si;
  assign so = so_unbuf;
  assign pcx_fpio_data_px2_buf1[123] = pcx_fpio_data_px2[123];
  assign pcx_fpio_data_px2_buf1[122] = pcx_fpio_data_px2[122];
  assign pcx_fpio_data_px2_buf1[121] = pcx_fpio_data_px2[121];
  assign pcx_fpio_data_px2_buf1[120] = pcx_fpio_data_px2[120];
  assign pcx_fpio_data_px2_buf1[119] = pcx_fpio_data_px2[119];
  assign pcx_fpio_data_px2_buf1[118] = pcx_fpio_data_px2[118];
  assign pcx_fpio_data_px2_buf1[117] = pcx_fpio_data_px2[117];
  assign pcx_fpio_data_px2_buf1[116] = pcx_fpio_data_px2[116];
  assign pcx_fpio_data_px2_buf1[115] = pcx_fpio_data_px2[115];
  assign pcx_fpio_data_px2_buf1[114] = pcx_fpio_data_px2[114];
  assign pcx_fpio_data_px2_buf1[113] = pcx_fpio_data_px2[113];
  assign pcx_fpio_data_px2_buf1[112] = pcx_fpio_data_px2[112];
  assign pcx_fpio_data_px2_buf1[111] = pcx_fpio_data_px2[111];
  assign pcx_fpio_data_px2_buf1[110] = pcx_fpio_data_px2[110];
  assign pcx_fpio_data_px2_buf1[109] = pcx_fpio_data_px2[109];
  assign pcx_fpio_data_px2_buf1[108] = pcx_fpio_data_px2[108];
  assign pcx_fpio_data_px2_buf1[107] = pcx_fpio_data_px2[107];
  assign pcx_fpio_data_px2_buf1[106] = pcx_fpio_data_px2[106];
  assign pcx_fpio_data_px2_buf1[105] = pcx_fpio_data_px2[105];
  assign pcx_fpio_data_px2_buf1[104] = pcx_fpio_data_px2[104];
  assign pcx_fpio_data_px2_buf1[103] = pcx_fpio_data_px2[103];
  assign pcx_fpio_data_px2_buf1[102] = pcx_fpio_data_px2[102];
  assign pcx_fpio_data_px2_buf1[101] = pcx_fpio_data_px2[101];
  assign pcx_fpio_data_px2_buf1[100] = pcx_fpio_data_px2[100];
  assign pcx_fpio_data_px2_buf1[99] = pcx_fpio_data_px2[99];
  assign pcx_fpio_data_px2_buf1[98] = pcx_fpio_data_px2[98];
  assign pcx_fpio_data_px2_buf1[97] = pcx_fpio_data_px2[97];
  assign pcx_fpio_data_px2_buf1[96] = pcx_fpio_data_px2[96];
  assign pcx_fpio_data_px2_buf1[95] = pcx_fpio_data_px2[95];
  assign pcx_fpio_data_px2_buf1[94] = pcx_fpio_data_px2[94];
  assign pcx_fpio_data_px2_buf1[93] = pcx_fpio_data_px2[93];
  assign pcx_fpio_data_px2_buf1[92] = pcx_fpio_data_px2[92];
  assign pcx_fpio_data_px2_buf1[91] = pcx_fpio_data_px2[91];
  assign pcx_fpio_data_px2_buf1[90] = pcx_fpio_data_px2[90];
  assign pcx_fpio_data_px2_buf1[89] = pcx_fpio_data_px2[89];
  assign pcx_fpio_data_px2_buf1[88] = pcx_fpio_data_px2[88];
  assign pcx_fpio_data_px2_buf1[87] = pcx_fpio_data_px2[87];
  assign pcx_fpio_data_px2_buf1[86] = pcx_fpio_data_px2[86];
  assign pcx_fpio_data_px2_buf1[85] = pcx_fpio_data_px2[85];
  assign pcx_fpio_data_px2_buf1[84] = pcx_fpio_data_px2[84];
  assign pcx_fpio_data_px2_buf1[83] = pcx_fpio_data_px2[83];
  assign pcx_fpio_data_px2_buf1[82] = pcx_fpio_data_px2[82];
  assign pcx_fpio_data_px2_buf1[81] = pcx_fpio_data_px2[81];
  assign pcx_fpio_data_px2_buf1[80] = pcx_fpio_data_px2[80];
  assign pcx_fpio_data_px2_buf1[79] = pcx_fpio_data_px2[79];
  assign pcx_fpio_data_px2_buf1[78] = pcx_fpio_data_px2[78];
  assign pcx_fpio_data_px2_buf1[77] = pcx_fpio_data_px2[77];
  assign pcx_fpio_data_px2_buf1[76] = pcx_fpio_data_px2[76];
  assign pcx_fpio_data_px2_buf1[75] = pcx_fpio_data_px2[75];
  assign pcx_fpio_data_px2_buf1[74] = pcx_fpio_data_px2[74];
  assign pcx_fpio_data_px2_buf1[73] = pcx_fpio_data_px2[73];
  assign pcx_fpio_data_px2_buf1[72] = pcx_fpio_data_px2[72];
  assign pcx_fpio_data_px2_buf1[71] = pcx_fpio_data_px2[71];
  assign pcx_fpio_data_px2_buf1[70] = pcx_fpio_data_px2[70];
  assign pcx_fpio_data_px2_buf1[69] = pcx_fpio_data_px2[69];
  assign pcx_fpio_data_px2_buf1[68] = pcx_fpio_data_px2[68];
  assign pcx_fpio_data_px2_buf1[67] = pcx_fpio_data_px2[67];
  assign pcx_fpio_data_px2_buf1[66] = pcx_fpio_data_px2[66];
  assign pcx_fpio_data_px2_buf1[65] = pcx_fpio_data_px2[65];
  assign pcx_fpio_data_px2_buf1[64] = pcx_fpio_data_px2[64];
  assign pcx_fpio_data_px2_buf1[63] = pcx_fpio_data_px2[63];
  assign pcx_fpio_data_px2_buf1[62] = pcx_fpio_data_px2[62];
  assign pcx_fpio_data_px2_buf1[61] = pcx_fpio_data_px2[61];
  assign pcx_fpio_data_px2_buf1[60] = pcx_fpio_data_px2[60];
  assign pcx_fpio_data_px2_buf1[59] = pcx_fpio_data_px2[59];
  assign pcx_fpio_data_px2_buf1[58] = pcx_fpio_data_px2[58];
  assign pcx_fpio_data_px2_buf1[57] = pcx_fpio_data_px2[57];
  assign pcx_fpio_data_px2_buf1[56] = pcx_fpio_data_px2[56];
  assign pcx_fpio_data_px2_buf1[55] = pcx_fpio_data_px2[55];
  assign pcx_fpio_data_px2_buf1[54] = pcx_fpio_data_px2[54];
  assign pcx_fpio_data_px2_buf1[53] = pcx_fpio_data_px2[53];
  assign pcx_fpio_data_px2_buf1[52] = pcx_fpio_data_px2[52];
  assign pcx_fpio_data_px2_buf1[51] = pcx_fpio_data_px2[51];
  assign pcx_fpio_data_px2_buf1[50] = pcx_fpio_data_px2[50];
  assign pcx_fpio_data_px2_buf1[49] = pcx_fpio_data_px2[49];
  assign pcx_fpio_data_px2_buf1[48] = pcx_fpio_data_px2[48];
  assign pcx_fpio_data_px2_buf1[47] = pcx_fpio_data_px2[47];
  assign pcx_fpio_data_px2_buf1[46] = pcx_fpio_data_px2[46];
  assign pcx_fpio_data_px2_buf1[45] = pcx_fpio_data_px2[45];
  assign pcx_fpio_data_px2_buf1[44] = pcx_fpio_data_px2[44];
  assign pcx_fpio_data_px2_buf1[43] = pcx_fpio_data_px2[43];
  assign pcx_fpio_data_px2_buf1[42] = pcx_fpio_data_px2[42];
  assign pcx_fpio_data_px2_buf1[41] = pcx_fpio_data_px2[41];
  assign pcx_fpio_data_px2_buf1[40] = pcx_fpio_data_px2[40];
  assign pcx_fpio_data_px2_buf1[39] = pcx_fpio_data_px2[39];
  assign pcx_fpio_data_px2_buf1[38] = pcx_fpio_data_px2[38];
  assign pcx_fpio_data_px2_buf1[37] = pcx_fpio_data_px2[37];
  assign pcx_fpio_data_px2_buf1[36] = pcx_fpio_data_px2[36];
  assign pcx_fpio_data_px2_buf1[35] = pcx_fpio_data_px2[35];
  assign pcx_fpio_data_px2_buf1[34] = pcx_fpio_data_px2[34];
  assign pcx_fpio_data_px2_buf1[33] = pcx_fpio_data_px2[33];
  assign pcx_fpio_data_px2_buf1[32] = pcx_fpio_data_px2[32];
  assign pcx_fpio_data_px2_buf1[31] = pcx_fpio_data_px2[31];
  assign pcx_fpio_data_px2_buf1[30] = pcx_fpio_data_px2[30];
  assign pcx_fpio_data_px2_buf1[29] = pcx_fpio_data_px2[29];
  assign pcx_fpio_data_px2_buf1[28] = pcx_fpio_data_px2[28];
  assign pcx_fpio_data_px2_buf1[27] = pcx_fpio_data_px2[27];
  assign pcx_fpio_data_px2_buf1[26] = pcx_fpio_data_px2[26];
  assign pcx_fpio_data_px2_buf1[25] = pcx_fpio_data_px2[25];
  assign pcx_fpio_data_px2_buf1[24] = pcx_fpio_data_px2[24];
  assign pcx_fpio_data_px2_buf1[23] = pcx_fpio_data_px2[23];
  assign pcx_fpio_data_px2_buf1[22] = pcx_fpio_data_px2[22];
  assign pcx_fpio_data_px2_buf1[21] = pcx_fpio_data_px2[21];
  assign pcx_fpio_data_px2_buf1[20] = pcx_fpio_data_px2[20];
  assign pcx_fpio_data_px2_buf1[19] = pcx_fpio_data_px2[19];
  assign pcx_fpio_data_px2_buf1[18] = pcx_fpio_data_px2[18];
  assign pcx_fpio_data_px2_buf1[17] = pcx_fpio_data_px2[17];
  assign pcx_fpio_data_px2_buf1[16] = pcx_fpio_data_px2[16];
  assign pcx_fpio_data_px2_buf1[15] = pcx_fpio_data_px2[15];
  assign pcx_fpio_data_px2_buf1[14] = pcx_fpio_data_px2[14];
  assign pcx_fpio_data_px2_buf1[13] = pcx_fpio_data_px2[13];
  assign pcx_fpio_data_px2_buf1[12] = pcx_fpio_data_px2[12];
  assign pcx_fpio_data_px2_buf1[11] = pcx_fpio_data_px2[11];
  assign pcx_fpio_data_px2_buf1[10] = pcx_fpio_data_px2[10];
  assign pcx_fpio_data_px2_buf1[9] = pcx_fpio_data_px2[9];
  assign pcx_fpio_data_px2_buf1[8] = pcx_fpio_data_px2[8];
  assign pcx_fpio_data_px2_buf1[7] = pcx_fpio_data_px2[7];
  assign pcx_fpio_data_px2_buf1[6] = pcx_fpio_data_px2[6];
  assign pcx_fpio_data_px2_buf1[5] = pcx_fpio_data_px2[5];
  assign pcx_fpio_data_px2_buf1[4] = pcx_fpio_data_px2[4];
  assign pcx_fpio_data_px2_buf1[3] = pcx_fpio_data_px2[3];
  assign pcx_fpio_data_px2_buf1[2] = pcx_fpio_data_px2[2];
  assign pcx_fpio_data_px2_buf1[1] = pcx_fpio_data_px2[1];
  assign pcx_fpio_data_px2_buf1[0] = pcx_fpio_data_px2[0];
  assign pcx_fpio_data_rdy_px2_buf1 = pcx_fpio_data_rdy_px2;
  assign fp_cpx_req_cq_buf1[7] = fp_cpx_req_cq[7];
  assign fp_cpx_req_cq_buf1[6] = fp_cpx_req_cq[6];
  assign fp_cpx_req_cq_buf1[5] = fp_cpx_req_cq[5];
  assign fp_cpx_req_cq_buf1[4] = fp_cpx_req_cq[4];
  assign fp_cpx_req_cq_buf1[3] = fp_cpx_req_cq[3];
  assign fp_cpx_req_cq_buf1[2] = fp_cpx_req_cq[2];
  assign fp_cpx_req_cq_buf1[1] = fp_cpx_req_cq[1];
  assign fp_cpx_req_cq_buf1[0] = fp_cpx_req_cq[0];
  assign fp_cpx_data_ca_buf1[144] = fp_cpx_data_ca[144];
  assign fp_cpx_data_ca_buf1[143] = fp_cpx_data_ca[143];
  assign fp_cpx_data_ca_buf1[142] = fp_cpx_data_ca[142];
  assign fp_cpx_data_ca_buf1[141] = fp_cpx_data_ca[141];
  assign fp_cpx_data_ca_buf1[140] = fp_cpx_data_ca[140];
  assign fp_cpx_data_ca_buf1[139] = fp_cpx_data_ca[139];
  assign fp_cpx_data_ca_buf1[138] = fp_cpx_data_ca[138];
  assign fp_cpx_data_ca_buf1[137] = fp_cpx_data_ca[137];
  assign fp_cpx_data_ca_buf1[136] = fp_cpx_data_ca[136];
  assign fp_cpx_data_ca_buf1[135] = fp_cpx_data_ca[135];
  assign fp_cpx_data_ca_buf1[134] = fp_cpx_data_ca[134];
  assign fp_cpx_data_ca_buf1[133] = fp_cpx_data_ca[133];
  assign fp_cpx_data_ca_buf1[132] = fp_cpx_data_ca[132];
  assign fp_cpx_data_ca_buf1[131] = fp_cpx_data_ca[131];
  assign fp_cpx_data_ca_buf1[130] = fp_cpx_data_ca[130];
  assign fp_cpx_data_ca_buf1[129] = fp_cpx_data_ca[129];
  assign fp_cpx_data_ca_buf1[128] = fp_cpx_data_ca[128];
  assign fp_cpx_data_ca_buf1[127] = fp_cpx_data_ca[127];
  assign fp_cpx_data_ca_buf1[126] = fp_cpx_data_ca[126];
  assign fp_cpx_data_ca_buf1[125] = fp_cpx_data_ca[125];
  assign fp_cpx_data_ca_buf1[124] = fp_cpx_data_ca[124];
  assign fp_cpx_data_ca_buf1[123] = fp_cpx_data_ca[123];
  assign fp_cpx_data_ca_buf1[122] = fp_cpx_data_ca[122];
  assign fp_cpx_data_ca_buf1[121] = fp_cpx_data_ca[121];
  assign fp_cpx_data_ca_buf1[120] = fp_cpx_data_ca[120];
  assign fp_cpx_data_ca_buf1[119] = fp_cpx_data_ca[119];
  assign fp_cpx_data_ca_buf1[118] = fp_cpx_data_ca[118];
  assign fp_cpx_data_ca_buf1[117] = fp_cpx_data_ca[117];
  assign fp_cpx_data_ca_buf1[116] = fp_cpx_data_ca[116];
  assign fp_cpx_data_ca_buf1[115] = fp_cpx_data_ca[115];
  assign fp_cpx_data_ca_buf1[114] = fp_cpx_data_ca[114];
  assign fp_cpx_data_ca_buf1[113] = fp_cpx_data_ca[113];
  assign fp_cpx_data_ca_buf1[112] = fp_cpx_data_ca[112];
  assign fp_cpx_data_ca_buf1[111] = fp_cpx_data_ca[111];
  assign fp_cpx_data_ca_buf1[110] = fp_cpx_data_ca[110];
  assign fp_cpx_data_ca_buf1[109] = fp_cpx_data_ca[109];
  assign fp_cpx_data_ca_buf1[108] = fp_cpx_data_ca[108];
  assign fp_cpx_data_ca_buf1[107] = fp_cpx_data_ca[107];
  assign fp_cpx_data_ca_buf1[106] = fp_cpx_data_ca[106];
  assign fp_cpx_data_ca_buf1[105] = fp_cpx_data_ca[105];
  assign fp_cpx_data_ca_buf1[104] = fp_cpx_data_ca[104];
  assign fp_cpx_data_ca_buf1[103] = fp_cpx_data_ca[103];
  assign fp_cpx_data_ca_buf1[102] = fp_cpx_data_ca[102];
  assign fp_cpx_data_ca_buf1[101] = fp_cpx_data_ca[101];
  assign fp_cpx_data_ca_buf1[100] = fp_cpx_data_ca[100];
  assign fp_cpx_data_ca_buf1[99] = fp_cpx_data_ca[99];
  assign fp_cpx_data_ca_buf1[98] = fp_cpx_data_ca[98];
  assign fp_cpx_data_ca_buf1[97] = fp_cpx_data_ca[97];
  assign fp_cpx_data_ca_buf1[96] = fp_cpx_data_ca[96];
  assign fp_cpx_data_ca_buf1[95] = fp_cpx_data_ca[95];
  assign fp_cpx_data_ca_buf1[94] = fp_cpx_data_ca[94];
  assign fp_cpx_data_ca_buf1[93] = fp_cpx_data_ca[93];
  assign fp_cpx_data_ca_buf1[92] = fp_cpx_data_ca[92];
  assign fp_cpx_data_ca_buf1[91] = fp_cpx_data_ca[91];
  assign fp_cpx_data_ca_buf1[90] = fp_cpx_data_ca[90];
  assign fp_cpx_data_ca_buf1[89] = fp_cpx_data_ca[89];
  assign fp_cpx_data_ca_buf1[88] = fp_cpx_data_ca[88];
  assign fp_cpx_data_ca_buf1[87] = fp_cpx_data_ca[87];
  assign fp_cpx_data_ca_buf1[86] = fp_cpx_data_ca[86];
  assign fp_cpx_data_ca_buf1[85] = fp_cpx_data_ca[85];
  assign fp_cpx_data_ca_buf1[84] = fp_cpx_data_ca[84];
  assign fp_cpx_data_ca_buf1[83] = fp_cpx_data_ca[83];
  assign fp_cpx_data_ca_buf1[82] = fp_cpx_data_ca[82];
  assign fp_cpx_data_ca_buf1[81] = fp_cpx_data_ca[81];
  assign fp_cpx_data_ca_buf1[80] = fp_cpx_data_ca[80];
  assign fp_cpx_data_ca_buf1[79] = fp_cpx_data_ca[79];
  assign fp_cpx_data_ca_buf1[78] = fp_cpx_data_ca[78];
  assign fp_cpx_data_ca_buf1[77] = fp_cpx_data_ca[77];
  assign fp_cpx_data_ca_buf1[76] = fp_cpx_data_ca[76];
  assign fp_cpx_data_ca_buf1[75] = fp_cpx_data_ca[75];
  assign fp_cpx_data_ca_buf1[74] = fp_cpx_data_ca[74];
  assign fp_cpx_data_ca_buf1[73] = fp_cpx_data_ca[73];
  assign fp_cpx_data_ca_buf1[72] = fp_cpx_data_ca[72];
  assign fp_cpx_data_ca_buf1[71] = fp_cpx_data_ca[71];
  assign fp_cpx_data_ca_buf1[70] = fp_cpx_data_ca[70];
  assign fp_cpx_data_ca_buf1[69] = fp_cpx_data_ca[69];
  assign fp_cpx_data_ca_buf1[68] = fp_cpx_data_ca[68];
  assign fp_cpx_data_ca_buf1[67] = fp_cpx_data_ca[67];
  assign fp_cpx_data_ca_buf1[66] = fp_cpx_data_ca[66];
  assign fp_cpx_data_ca_buf1[65] = fp_cpx_data_ca[65];
  assign fp_cpx_data_ca_buf1[64] = fp_cpx_data_ca[64];
  assign fp_cpx_data_ca_buf1[63] = fp_cpx_data_ca[63];
  assign fp_cpx_data_ca_buf1[62] = fp_cpx_data_ca[62];
  assign fp_cpx_data_ca_buf1[61] = fp_cpx_data_ca[61];
  assign fp_cpx_data_ca_buf1[60] = fp_cpx_data_ca[60];
  assign fp_cpx_data_ca_buf1[59] = fp_cpx_data_ca[59];
  assign fp_cpx_data_ca_buf1[58] = fp_cpx_data_ca[58];
  assign fp_cpx_data_ca_buf1[57] = fp_cpx_data_ca[57];
  assign fp_cpx_data_ca_buf1[56] = fp_cpx_data_ca[56];
  assign fp_cpx_data_ca_buf1[55] = fp_cpx_data_ca[55];
  assign fp_cpx_data_ca_buf1[54] = fp_cpx_data_ca[54];
  assign fp_cpx_data_ca_buf1[53] = fp_cpx_data_ca[53];
  assign fp_cpx_data_ca_buf1[52] = fp_cpx_data_ca[52];
  assign fp_cpx_data_ca_buf1[51] = fp_cpx_data_ca[51];
  assign fp_cpx_data_ca_buf1[50] = fp_cpx_data_ca[50];
  assign fp_cpx_data_ca_buf1[49] = fp_cpx_data_ca[49];
  assign fp_cpx_data_ca_buf1[48] = fp_cpx_data_ca[48];
  assign fp_cpx_data_ca_buf1[47] = fp_cpx_data_ca[47];
  assign fp_cpx_data_ca_buf1[46] = fp_cpx_data_ca[46];
  assign fp_cpx_data_ca_buf1[45] = fp_cpx_data_ca[45];
  assign fp_cpx_data_ca_buf1[44] = fp_cpx_data_ca[44];
  assign fp_cpx_data_ca_buf1[43] = fp_cpx_data_ca[43];
  assign fp_cpx_data_ca_buf1[42] = fp_cpx_data_ca[42];
  assign fp_cpx_data_ca_buf1[41] = fp_cpx_data_ca[41];
  assign fp_cpx_data_ca_buf1[40] = fp_cpx_data_ca[40];
  assign fp_cpx_data_ca_buf1[39] = fp_cpx_data_ca[39];
  assign fp_cpx_data_ca_buf1[38] = fp_cpx_data_ca[38];
  assign fp_cpx_data_ca_buf1[37] = fp_cpx_data_ca[37];
  assign fp_cpx_data_ca_buf1[36] = fp_cpx_data_ca[36];
  assign fp_cpx_data_ca_buf1[35] = fp_cpx_data_ca[35];
  assign fp_cpx_data_ca_buf1[34] = fp_cpx_data_ca[34];
  assign fp_cpx_data_ca_buf1[33] = fp_cpx_data_ca[33];
  assign fp_cpx_data_ca_buf1[32] = fp_cpx_data_ca[32];
  assign fp_cpx_data_ca_buf1[31] = fp_cpx_data_ca[31];
  assign fp_cpx_data_ca_buf1[30] = fp_cpx_data_ca[30];
  assign fp_cpx_data_ca_buf1[29] = fp_cpx_data_ca[29];
  assign fp_cpx_data_ca_buf1[28] = fp_cpx_data_ca[28];
  assign fp_cpx_data_ca_buf1[27] = fp_cpx_data_ca[27];
  assign fp_cpx_data_ca_buf1[26] = fp_cpx_data_ca[26];
  assign fp_cpx_data_ca_buf1[25] = fp_cpx_data_ca[25];
  assign fp_cpx_data_ca_buf1[24] = fp_cpx_data_ca[24];
  assign fp_cpx_data_ca_buf1[23] = fp_cpx_data_ca[23];
  assign fp_cpx_data_ca_buf1[22] = fp_cpx_data_ca[22];
  assign fp_cpx_data_ca_buf1[21] = fp_cpx_data_ca[21];
  assign fp_cpx_data_ca_buf1[20] = fp_cpx_data_ca[20];
  assign fp_cpx_data_ca_buf1[19] = fp_cpx_data_ca[19];
  assign fp_cpx_data_ca_buf1[18] = fp_cpx_data_ca[18];
  assign fp_cpx_data_ca_buf1[17] = fp_cpx_data_ca[17];
  assign fp_cpx_data_ca_buf1[16] = fp_cpx_data_ca[16];
  assign fp_cpx_data_ca_buf1[15] = fp_cpx_data_ca[15];
  assign fp_cpx_data_ca_buf1[14] = fp_cpx_data_ca[14];
  assign fp_cpx_data_ca_buf1[13] = fp_cpx_data_ca[13];
  assign fp_cpx_data_ca_buf1[12] = fp_cpx_data_ca[12];
  assign fp_cpx_data_ca_buf1[11] = fp_cpx_data_ca[11];
  assign fp_cpx_data_ca_buf1[10] = fp_cpx_data_ca[10];
  assign fp_cpx_data_ca_buf1[9] = fp_cpx_data_ca[9];
  assign fp_cpx_data_ca_buf1[8] = fp_cpx_data_ca[8];
  assign fp_cpx_data_ca_buf1[7] = fp_cpx_data_ca[7];
  assign fp_cpx_data_ca_buf1[6] = fp_cpx_data_ca[6];
  assign fp_cpx_data_ca_buf1[5] = fp_cpx_data_ca[5];
  assign fp_cpx_data_ca_buf1[4] = fp_cpx_data_ca[4];
  assign fp_cpx_data_ca_buf1[3] = fp_cpx_data_ca[3];
  assign fp_cpx_data_ca_buf1[2] = fp_cpx_data_ca[2];
  assign fp_cpx_data_ca_buf1[1] = fp_cpx_data_ca[1];
  assign fp_cpx_data_ca_buf1[0] = fp_cpx_data_ca[0];
  assign inq_sram_din_buf1[155] = inq_sram_din_unbuf[155];
  assign inq_sram_din_buf1[154] = inq_sram_din_unbuf[154];
  assign inq_sram_din_buf1[153] = inq_sram_din_unbuf[153];
  assign inq_sram_din_buf1[152] = inq_sram_din_unbuf[152];
  assign inq_sram_din_buf1[151] = inq_sram_din_unbuf[151];
  assign inq_sram_din_buf1[150] = inq_sram_din_unbuf[150];
  assign inq_sram_din_buf1[149] = inq_sram_din_unbuf[149];
  assign inq_sram_din_buf1[148] = inq_sram_din_unbuf[148];
  assign inq_sram_din_buf1[147] = inq_sram_din_unbuf[147];
  assign inq_sram_din_buf1[146] = inq_sram_din_unbuf[146];
  assign inq_sram_din_buf1[145] = inq_sram_din_unbuf[145];
  assign inq_sram_din_buf1[144] = inq_sram_din_unbuf[144];
  assign inq_sram_din_buf1[143] = inq_sram_din_unbuf[143];
  assign inq_sram_din_buf1[142] = inq_sram_din_unbuf[142];
  assign inq_sram_din_buf1[141] = inq_sram_din_unbuf[141];
  assign inq_sram_din_buf1[140] = inq_sram_din_unbuf[140];
  assign inq_sram_din_buf1[139] = inq_sram_din_unbuf[139];
  assign inq_sram_din_buf1[138] = inq_sram_din_unbuf[138];
  assign inq_sram_din_buf1[137] = inq_sram_din_unbuf[137];
  assign inq_sram_din_buf1[136] = inq_sram_din_unbuf[136];
  assign inq_sram_din_buf1[135] = inq_sram_din_unbuf[135];
  assign inq_sram_din_buf1[134] = inq_sram_din_unbuf[134];
  assign inq_sram_din_buf1[133] = inq_sram_din_unbuf[133];
  assign inq_sram_din_buf1[132] = inq_sram_din_unbuf[132];
  assign inq_sram_din_buf1[131] = inq_sram_din_unbuf[131];
  assign inq_sram_din_buf1[130] = inq_sram_din_unbuf[130];
  assign inq_sram_din_buf1[129] = inq_sram_din_unbuf[129];
  assign inq_sram_din_buf1[128] = inq_sram_din_unbuf[128];
  assign inq_sram_din_buf1[127] = inq_sram_din_unbuf[127];
  assign inq_sram_din_buf1[126] = inq_sram_din_unbuf[126];
  assign inq_sram_din_buf1[125] = inq_sram_din_unbuf[125];
  assign inq_sram_din_buf1[124] = inq_sram_din_unbuf[124];
  assign inq_sram_din_buf1[123] = inq_sram_din_unbuf[123];
  assign inq_sram_din_buf1[122] = inq_sram_din_unbuf[122];
  assign inq_sram_din_buf1[121] = inq_sram_din_unbuf[121];
  assign inq_sram_din_buf1[120] = inq_sram_din_unbuf[120];
  assign inq_sram_din_buf1[119] = inq_sram_din_unbuf[119];
  assign inq_sram_din_buf1[118] = inq_sram_din_unbuf[118];
  assign inq_sram_din_buf1[117] = inq_sram_din_unbuf[117];
  assign inq_sram_din_buf1[116] = inq_sram_din_unbuf[116];
  assign inq_sram_din_buf1[115] = inq_sram_din_unbuf[115];
  assign inq_sram_din_buf1[114] = inq_sram_din_unbuf[114];
  assign inq_sram_din_buf1[113] = inq_sram_din_unbuf[113];
  assign inq_sram_din_buf1[112] = inq_sram_din_unbuf[112];
  assign inq_sram_din_buf1[111] = inq_sram_din_unbuf[111];
  assign inq_sram_din_buf1[110] = inq_sram_din_unbuf[110];
  assign inq_sram_din_buf1[109] = inq_sram_din_unbuf[109];
  assign inq_sram_din_buf1[108] = inq_sram_din_unbuf[108];
  assign inq_sram_din_buf1[107] = inq_sram_din_unbuf[107];
  assign inq_sram_din_buf1[106] = inq_sram_din_unbuf[106];
  assign inq_sram_din_buf1[105] = inq_sram_din_unbuf[105];
  assign inq_sram_din_buf1[104] = inq_sram_din_unbuf[104];
  assign inq_sram_din_buf1[103] = inq_sram_din_unbuf[103];
  assign inq_sram_din_buf1[102] = inq_sram_din_unbuf[102];
  assign inq_sram_din_buf1[101] = inq_sram_din_unbuf[101];
  assign inq_sram_din_buf1[100] = inq_sram_din_unbuf[100];
  assign inq_sram_din_buf1[99] = inq_sram_din_unbuf[99];
  assign inq_sram_din_buf1[98] = inq_sram_din_unbuf[98];
  assign inq_sram_din_buf1[97] = inq_sram_din_unbuf[97];
  assign inq_sram_din_buf1[96] = inq_sram_din_unbuf[96];
  assign inq_sram_din_buf1[95] = inq_sram_din_unbuf[95];
  assign inq_sram_din_buf1[94] = inq_sram_din_unbuf[94];
  assign inq_sram_din_buf1[93] = inq_sram_din_unbuf[93];
  assign inq_sram_din_buf1[92] = inq_sram_din_unbuf[92];
  assign inq_sram_din_buf1[91] = inq_sram_din_unbuf[91];
  assign inq_sram_din_buf1[90] = inq_sram_din_unbuf[90];
  assign inq_sram_din_buf1[89] = inq_sram_din_unbuf[89];
  assign inq_sram_din_buf1[88] = inq_sram_din_unbuf[88];
  assign inq_sram_din_buf1[87] = inq_sram_din_unbuf[87];
  assign inq_sram_din_buf1[86] = inq_sram_din_unbuf[86];
  assign inq_sram_din_buf1[85] = inq_sram_din_unbuf[85];
  assign inq_sram_din_buf1[84] = inq_sram_din_unbuf[84];
  assign inq_sram_din_buf1[83] = inq_sram_din_unbuf[83];
  assign inq_sram_din_buf1[82] = inq_sram_din_unbuf[82];
  assign inq_sram_din_buf1[81] = inq_sram_din_unbuf[81];
  assign inq_sram_din_buf1[80] = inq_sram_din_unbuf[80];
  assign inq_sram_din_buf1[79] = inq_sram_din_unbuf[79];
  assign inq_sram_din_buf1[78] = inq_sram_din_unbuf[78];
  assign inq_sram_din_buf1[77] = inq_sram_din_unbuf[77];
  assign inq_sram_din_buf1[76] = inq_sram_din_unbuf[76];
  assign inq_sram_din_buf1[75] = inq_sram_din_unbuf[75];
  assign inq_sram_din_buf1[74] = inq_sram_din_unbuf[74];
  assign inq_sram_din_buf1[73] = inq_sram_din_unbuf[73];
  assign inq_sram_din_buf1[72] = inq_sram_din_unbuf[72];
  assign inq_sram_din_buf1[71] = inq_sram_din_unbuf[71];
  assign inq_sram_din_buf1[70] = inq_sram_din_unbuf[70];
  assign inq_sram_din_buf1[69] = inq_sram_din_unbuf[69];
  assign inq_sram_din_buf1[68] = inq_sram_din_unbuf[68];
  assign inq_sram_din_buf1[67] = inq_sram_din_unbuf[67];
  assign inq_sram_din_buf1[66] = inq_sram_din_unbuf[66];
  assign inq_sram_din_buf1[65] = inq_sram_din_unbuf[65];
  assign inq_sram_din_buf1[64] = inq_sram_din_unbuf[64];
  assign inq_sram_din_buf1[63] = inq_sram_din_unbuf[63];
  assign inq_sram_din_buf1[62] = inq_sram_din_unbuf[62];
  assign inq_sram_din_buf1[61] = inq_sram_din_unbuf[61];
  assign inq_sram_din_buf1[60] = inq_sram_din_unbuf[60];
  assign inq_sram_din_buf1[59] = inq_sram_din_unbuf[59];
  assign inq_sram_din_buf1[58] = inq_sram_din_unbuf[58];
  assign inq_sram_din_buf1[57] = inq_sram_din_unbuf[57];
  assign inq_sram_din_buf1[56] = inq_sram_din_unbuf[56];
  assign inq_sram_din_buf1[55] = inq_sram_din_unbuf[55];
  assign inq_sram_din_buf1[54] = inq_sram_din_unbuf[54];
  assign inq_sram_din_buf1[53] = inq_sram_din_unbuf[53];
  assign inq_sram_din_buf1[52] = inq_sram_din_unbuf[52];
  assign inq_sram_din_buf1[51] = inq_sram_din_unbuf[51];
  assign inq_sram_din_buf1[50] = inq_sram_din_unbuf[50];
  assign inq_sram_din_buf1[49] = inq_sram_din_unbuf[49];
  assign inq_sram_din_buf1[48] = inq_sram_din_unbuf[48];
  assign inq_sram_din_buf1[47] = inq_sram_din_unbuf[47];
  assign inq_sram_din_buf1[46] = inq_sram_din_unbuf[46];
  assign inq_sram_din_buf1[45] = inq_sram_din_unbuf[45];
  assign inq_sram_din_buf1[44] = inq_sram_din_unbuf[44];
  assign inq_sram_din_buf1[43] = inq_sram_din_unbuf[43];
  assign inq_sram_din_buf1[42] = inq_sram_din_unbuf[42];
  assign inq_sram_din_buf1[41] = inq_sram_din_unbuf[41];
  assign inq_sram_din_buf1[40] = inq_sram_din_unbuf[40];
  assign inq_sram_din_buf1[39] = inq_sram_din_unbuf[39];
  assign inq_sram_din_buf1[38] = inq_sram_din_unbuf[38];
  assign inq_sram_din_buf1[37] = inq_sram_din_unbuf[37];
  assign inq_sram_din_buf1[36] = inq_sram_din_unbuf[36];
  assign inq_sram_din_buf1[35] = inq_sram_din_unbuf[35];
  assign inq_sram_din_buf1[34] = inq_sram_din_unbuf[34];
  assign inq_sram_din_buf1[33] = inq_sram_din_unbuf[33];
  assign inq_sram_din_buf1[32] = inq_sram_din_unbuf[32];
  assign inq_sram_din_buf1[31] = inq_sram_din_unbuf[31];
  assign inq_sram_din_buf1[30] = inq_sram_din_unbuf[30];
  assign inq_sram_din_buf1[29] = inq_sram_din_unbuf[29];
  assign inq_sram_din_buf1[28] = inq_sram_din_unbuf[28];
  assign inq_sram_din_buf1[27] = inq_sram_din_unbuf[27];
  assign inq_sram_din_buf1[26] = inq_sram_din_unbuf[26];
  assign inq_sram_din_buf1[25] = inq_sram_din_unbuf[25];
  assign inq_sram_din_buf1[24] = inq_sram_din_unbuf[24];
  assign inq_sram_din_buf1[23] = inq_sram_din_unbuf[23];
  assign inq_sram_din_buf1[22] = inq_sram_din_unbuf[22];
  assign inq_sram_din_buf1[21] = inq_sram_din_unbuf[21];
  assign inq_sram_din_buf1[20] = inq_sram_din_unbuf[20];
  assign inq_sram_din_buf1[19] = inq_sram_din_unbuf[19];
  assign inq_sram_din_buf1[18] = inq_sram_din_unbuf[18];
  assign inq_sram_din_buf1[17] = inq_sram_din_unbuf[17];
  assign inq_sram_din_buf1[16] = inq_sram_din_unbuf[16];
  assign inq_sram_din_buf1[15] = inq_sram_din_unbuf[15];
  assign inq_sram_din_buf1[14] = inq_sram_din_unbuf[14];
  assign inq_sram_din_buf1[13] = inq_sram_din_unbuf[13];
  assign inq_sram_din_buf1[12] = inq_sram_din_unbuf[12];
  assign inq_sram_din_buf1[11] = inq_sram_din_unbuf[11];
  assign inq_sram_din_buf1[10] = inq_sram_din_unbuf[10];
  assign inq_sram_din_buf1[9] = inq_sram_din_unbuf[9];
  assign inq_sram_din_buf1[8] = inq_sram_din_unbuf[8];
  assign inq_sram_din_buf1[7] = inq_sram_din_unbuf[7];
  assign inq_sram_din_buf1[6] = inq_sram_din_unbuf[6];
  assign inq_sram_din_buf1[5] = inq_sram_din_unbuf[5];
  assign inq_sram_din_buf1[4] = inq_sram_din_unbuf[4];
  assign inq_sram_din_buf1[3] = inq_sram_din_unbuf[3];
  assign inq_sram_din_buf1[2] = inq_sram_din_unbuf[2];
  assign inq_sram_din_buf1[1] = inq_sram_din_unbuf[1];
  assign inq_sram_din_buf1[0] = inq_sram_din_unbuf[0];

endmodule

