
module fpu_mul ( inq_op, inq_rnd_mode, inq_id, inq_in1, inq_in1_53_0_neq_0, 
        inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1_exp_eq_0, 
        inq_in1_exp_neq_ffs, inq_in2, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0, 
        inq_in2_53_32_neq_0, inq_in2_exp_eq_0, inq_in2_exp_neq_ffs, inq_mul, 
        mul_dest_rdy, mul_dest_rdya, fmul_clken_l, fmul_clken_l_buf1, arst_l, 
        grst_l, rclk, mul_pipe_active, m1stg_step, m6stg_fmul_in, m6stg_id_in, 
        mul_exc_out, m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out, 
        mul_exp_out, mul_frac_out, se_mul, se_mul64, si, so );
  input [7:0] inq_op;
  input [1:0] inq_rnd_mode;
  input [4:0] inq_id;
  input [63:0] inq_in1;
  input [63:0] inq_in2;
  output [9:0] m6stg_id_in;
  output [4:0] mul_exc_out;
  output [10:0] mul_exp_out;
  output [51:0] mul_frac_out;
  input inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0,
         inq_in1_exp_eq_0, inq_in1_exp_neq_ffs, inq_in2_53_0_neq_0,
         inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2_exp_eq_0,
         inq_in2_exp_neq_ffs, inq_mul, mul_dest_rdy, mul_dest_rdya,
         fmul_clken_l, fmul_clken_l_buf1, arst_l, grst_l, rclk, se_mul,
         se_mul64, si;
  output mul_pipe_active, m1stg_step, m6stg_fmul_in, m6stg_fmul_dbl_dst,
         m6stg_fmuls, mul_sign_out, so;
  wire   m1stg_sngop, m1stg_dblop, m1stg_dblop_inv, m2stg_fmuls, m2stg_fmuld,
         m2stg_fsmuld, m5stg_fmuls, m5stg_fmuld, m5stg_fmulda, m2stg_exp_017f,
         m4stg_inc_exp_54, m4stg_inc_exp_55, m4stg_inc_exp_105, mul_rst_l,
         m4stg_frac_105, m4stg_shl_54, m4stg_shl_55,
         \fpu_mul_exp_dp/m5stg_inc_exp_105 , \fpu_mul_exp_dp/m5stg_inc_exp_55 ,
         \fpu_mul_exp_dp/m5stg_inc_exp_54 , \fpu_mul_exp_dp/m5stg_shl_54 ,
         \fpu_mul_exp_dp/m5stg_shl_55 , \fpu_mul_exp_dp/m5stg_exp_pre2[11] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[10] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[9] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[8] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[7] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[6] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[5] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[4] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[3] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[2] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[1] ,
         \fpu_mul_exp_dp/m5stg_exp_pre2[0] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[12] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[11] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[10] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[9] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[8] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[7] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[6] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[5] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[4] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[3] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[2] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[1] ,
         \fpu_mul_exp_dp/m5stg_exp_pre1[0] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[11] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[10] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[9] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[8] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[7] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[6] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[5] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[4] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[3] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[2] ,
         \fpu_mul_exp_dp/m4stg_exp_plus1[1] , \fpu_mul_exp_dp/m3stg_expa[12] ,
         \fpu_mul_exp_dp/m3stg_expa[11] , \fpu_mul_exp_dp/m3stg_expa[9] ,
         \fpu_mul_exp_dp/m3stg_expa[8] , \fpu_mul_exp_dp/m3stg_expa[1] ,
         \fpu_mul_exp_dp/m3bstg_exp[9] , \fpu_mul_exp_dp/m3bstg_exp[11] ,
         \fpu_mul_exp_dp/m2stg_exp[12] , \fpu_mul_exp_dp/m2stg_exp[8] ,
         \fpu_mul_exp_dp/ckbuf_mul_exp_dp/clken ,
         \fpu_mul_exp_dp/ckbuf_mul_exp_dp/N1 , n4, n5, n6, n7, n8, n9, n10,
         n12, n17, n18, n20, n22, n24, n26, n28, n29, n30, n32, n34, n36, n37,
         n38, n40, n43, n44, n45, n47, n49, n51, n52, n53, n55, n57, n59, n60,
         n61, n63, n94, n98, n103, n104, n106, n107, n110, n111, n112, n114,
         n115, n118, n119, n120, n122, n130, n132, n134, n135, n136, n137,
         n138, n140, n142, n143, n144, n145, n146, n147, n148, n156, n158,
         n160, n162, n164, n166, n168, n172, n174, n176, n178, n180, n189,
         n190, n191, n192, n193, n194, n195, n196, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n269, n270, n271,
         n272, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n438, n439, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n452, n453, n454, n455, n456, n594, n603, n604, n709, n876, n877,
         n878, \fpu_mul_ctl/n735 , \fpu_mul_ctl/n733 , \fpu_mul_ctl/n732 ,
         \fpu_mul_ctl/n731 , \fpu_mul_ctl/n730 , \fpu_mul_ctl/n105 ,
         \fpu_mul_ctl/n273 , \fpu_mul_ctl/n272 , \fpu_mul_ctl/n271 ,
         \fpu_mul_ctl/n270 , \fpu_mul_ctl/n269 , \fpu_mul_ctl/n268 ,
         \fpu_mul_ctl/n267 , \fpu_mul_ctl/n266 , \fpu_mul_ctl/n265 ,
         \fpu_mul_ctl/n264 , \fpu_mul_ctl/n263 , \fpu_mul_ctl/n262 ,
         \fpu_mul_ctl/n261 , \fpu_mul_ctl/n260 , \fpu_mul_ctl/n259 ,
         \fpu_mul_ctl/n257 , \fpu_mul_ctl/n256 , \fpu_mul_ctl/n253 ,
         \fpu_mul_ctl/n561 , \fpu_mul_ctl/n560 , \fpu_mul_ctl/n559 ,
         \fpu_mul_ctl/n558 , \fpu_mul_ctl/n557 , \fpu_mul_ctl/n556 ,
         \fpu_mul_ctl/n555 , \fpu_mul_ctl/n554 , \fpu_mul_ctl/n553 ,
         \fpu_mul_ctl/n552 , \fpu_mul_ctl/n551 , \fpu_mul_ctl/n550 ,
         \fpu_mul_ctl/n549 , \fpu_mul_ctl/n548 , \fpu_mul_ctl/n547 ,
         \fpu_mul_ctl/n546 , \fpu_mul_ctl/n545 , \fpu_mul_ctl/n544 ,
         \fpu_mul_ctl/n543 , \fpu_mul_ctl/n542 , \fpu_mul_ctl/n541 ,
         \fpu_mul_ctl/n540 , \fpu_mul_ctl/n539 , \fpu_mul_ctl/n538 ,
         \fpu_mul_ctl/n537 , \fpu_mul_ctl/n536 , \fpu_mul_ctl/n535 ,
         \fpu_mul_ctl/n534 , \fpu_mul_ctl/n533 , \fpu_mul_ctl/n532 ,
         \fpu_mul_ctl/n531 , \fpu_mul_ctl/n530 , \fpu_mul_ctl/n529 ,
         \fpu_mul_ctl/n528 , \fpu_mul_ctl/n527 , \fpu_mul_ctl/n526 ,
         \fpu_mul_ctl/n525 , \fpu_mul_ctl/n524 , \fpu_mul_ctl/n523 ,
         \fpu_mul_ctl/n522 , \fpu_mul_ctl/n521 , \fpu_mul_ctl/n520 ,
         \fpu_mul_ctl/n519 , \fpu_mul_ctl/n518 , \fpu_mul_ctl/n517 ,
         \fpu_mul_ctl/n516 , \fpu_mul_ctl/n515 , \fpu_mul_ctl/n514 ,
         \fpu_mul_ctl/n513 , \fpu_mul_ctl/n512 , \fpu_mul_ctl/n511 ,
         \fpu_mul_ctl/n510 , \fpu_mul_ctl/n509 , \fpu_mul_ctl/n508 ,
         \fpu_mul_ctl/n507 , \fpu_mul_ctl/n506 , \fpu_mul_ctl/n505 ,
         \fpu_mul_ctl/n504 , \fpu_mul_ctl/n503 , \fpu_mul_ctl/n502 ,
         \fpu_mul_ctl/n501 , \fpu_mul_ctl/n500 , \fpu_mul_ctl/n499 ,
         \fpu_mul_ctl/n498 , \fpu_mul_ctl/n497 , \fpu_mul_ctl/n496 ,
         \fpu_mul_ctl/n495 , \fpu_mul_ctl/n494 , \fpu_mul_ctl/n493 ,
         \fpu_mul_ctl/n492 , \fpu_mul_ctl/n491 , \fpu_mul_ctl/n490 ,
         \fpu_mul_ctl/n489 , \fpu_mul_ctl/n488 , \fpu_mul_ctl/n487 ,
         \fpu_mul_ctl/n486 , \fpu_mul_ctl/n485 , \fpu_mul_ctl/n484 ,
         \fpu_mul_ctl/n483 , \fpu_mul_ctl/n482 , \fpu_mul_ctl/n481 ,
         \fpu_mul_ctl/n480 , \fpu_mul_ctl/n479 , \fpu_mul_ctl/n478 ,
         \fpu_mul_ctl/n477 , \fpu_mul_ctl/n476 , \fpu_mul_ctl/n475 ,
         \fpu_mul_ctl/n474 , \fpu_mul_ctl/n473 , \fpu_mul_ctl/n472 ,
         \fpu_mul_ctl/n471 , \fpu_mul_ctl/n470 , \fpu_mul_ctl/n469 ,
         \fpu_mul_ctl/n468 , \fpu_mul_ctl/n467 , \fpu_mul_ctl/n466 ,
         \fpu_mul_ctl/n465 , \fpu_mul_ctl/n464 , \fpu_mul_ctl/n463 ,
         \fpu_mul_ctl/n462 , \fpu_mul_ctl/n461 , \fpu_mul_ctl/n460 ,
         \fpu_mul_ctl/n459 , \fpu_mul_ctl/n458 , \fpu_mul_ctl/n457 ,
         \fpu_mul_ctl/n456 , \fpu_mul_ctl/n455 , \fpu_mul_ctl/n454 ,
         \fpu_mul_ctl/n453 , \fpu_mul_ctl/n452 , \fpu_mul_ctl/n451 ,
         \fpu_mul_ctl/n450 , \fpu_mul_ctl/n449 , \fpu_mul_ctl/n448 ,
         \fpu_mul_ctl/n447 , \fpu_mul_ctl/n446 , \fpu_mul_ctl/n445 ,
         \fpu_mul_ctl/n444 , \fpu_mul_ctl/n443 , \fpu_mul_ctl/n442 ,
         \fpu_mul_ctl/n441 , \fpu_mul_ctl/n440 , \fpu_mul_ctl/n439 ,
         \fpu_mul_ctl/n438 , \fpu_mul_ctl/n437 , \fpu_mul_ctl/n436 ,
         \fpu_mul_ctl/n435 , \fpu_mul_ctl/n434 , \fpu_mul_ctl/n433 ,
         \fpu_mul_ctl/n432 , \fpu_mul_ctl/n431 , \fpu_mul_ctl/n430 ,
         \fpu_mul_ctl/n429 , \fpu_mul_ctl/n428 , \fpu_mul_ctl/n427 ,
         \fpu_mul_ctl/n426 , \fpu_mul_ctl/n425 , \fpu_mul_ctl/n424 ,
         \fpu_mul_ctl/n423 , \fpu_mul_ctl/n422 , \fpu_mul_ctl/n421 ,
         \fpu_mul_ctl/n420 , \fpu_mul_ctl/n419 , \fpu_mul_ctl/n418 ,
         \fpu_mul_ctl/n417 , \fpu_mul_ctl/n416 , \fpu_mul_ctl/n415 ,
         \fpu_mul_ctl/n414 , \fpu_mul_ctl/n413 , \fpu_mul_ctl/n412 ,
         \fpu_mul_ctl/n411 , \fpu_mul_ctl/n410 , \fpu_mul_ctl/n409 ,
         \fpu_mul_ctl/n408 , \fpu_mul_ctl/n407 , \fpu_mul_ctl/n406 ,
         \fpu_mul_ctl/n405 , \fpu_mul_ctl/n404 , \fpu_mul_ctl/n403 ,
         \fpu_mul_ctl/n402 , \fpu_mul_ctl/n401 , \fpu_mul_ctl/n400 ,
         \fpu_mul_ctl/n399 , \fpu_mul_ctl/n398 , \fpu_mul_ctl/n397 ,
         \fpu_mul_ctl/n396 , \fpu_mul_ctl/n395 , \fpu_mul_ctl/n394 ,
         \fpu_mul_ctl/n393 , \fpu_mul_ctl/n392 , \fpu_mul_ctl/n391 ,
         \fpu_mul_ctl/n390 , \fpu_mul_ctl/n389 , \fpu_mul_ctl/n388 ,
         \fpu_mul_ctl/n387 , \fpu_mul_ctl/n386 , \fpu_mul_ctl/n385 ,
         \fpu_mul_ctl/n384 , \fpu_mul_ctl/n380 , \fpu_mul_ctl/n379 ,
         \fpu_mul_ctl/n163 , \fpu_mul_ctl/n156 , \fpu_mul_ctl/n143 ,
         \fpu_mul_ctl/n142 , \fpu_mul_ctl/n141 , \fpu_mul_ctl/n140 ,
         \fpu_mul_ctl/n139 , \fpu_mul_ctl/n138 , \fpu_mul_ctl/n137 ,
         \fpu_mul_ctl/n136 , \fpu_mul_ctl/n135 , \fpu_mul_ctl/n134 ,
         \fpu_mul_ctl/n133 , \fpu_mul_ctl/n132 , \fpu_mul_ctl/n131 ,
         \fpu_mul_ctl/n130 , \fpu_mul_ctl/n123 , \fpu_mul_ctl/n120 ,
         \fpu_mul_ctl/n117 , \fpu_mul_ctl/n116 , \fpu_mul_ctl/n112 ,
         \fpu_mul_ctl/n111 , \fpu_mul_ctl/n110 , \fpu_mul_ctl/n107 ,
         \fpu_mul_ctl/n106 , \fpu_mul_ctl/n104 , \fpu_mul_ctl/n103 ,
         \fpu_mul_ctl/n102 , \fpu_mul_ctl/n100 , \fpu_mul_ctl/n98 ,
         \fpu_mul_ctl/n97 , \fpu_mul_ctl/n96 , \fpu_mul_ctl/n95 ,
         \fpu_mul_ctl/n94 , \fpu_mul_ctl/n93 , \fpu_mul_ctl/n52 ,
         \fpu_mul_ctl/n51 , \fpu_mul_ctl/n50 , \fpu_mul_ctl/n32 ,
         \fpu_mul_ctl/n31 , \fpu_mul_ctl/n30 , \fpu_mul_ctl/n28 ,
         \fpu_mul_ctl/n26 , \fpu_mul_ctl/n25 , \fpu_mul_ctl/n24 ,
         \fpu_mul_ctl/n23 , \fpu_mul_ctl/n22 , \fpu_mul_ctl/n20 ,
         \fpu_mul_ctl/n19 , \fpu_mul_ctl/n18 , \fpu_mul_ctl/n17 ,
         \fpu_mul_ctl/n16 , \fpu_mul_ctl/n1 , \fpu_mul_ctl/i_m1stg_mul/N3 ,
         \fpu_mul_ctl/i_m1stg_op/N3 , \fpu_mul_ctl/i_m1stg_op/N4 ,
         \fpu_mul_ctl/i_m1stg_op/N5 , \fpu_mul_ctl/i_m1stg_op/N6 ,
         \fpu_mul_ctl/i_m1stg_op/N7 , \fpu_mul_ctl/i_m1stg_op/N8 ,
         \fpu_mul_ctl/i_m1stg_op/N9 , \fpu_mul_ctl/i_m1stg_op/N10 ,
         \fpu_mul_ctl/dffrl_mul_ctl/N4 , \fpu_mul_ctl/m4stg_right_shift ,
         \fpu_mul_ctl/m4stg_expadd_eq_0 , \fpu_mul_ctl/m2stg_ld0_2[3] ,
         \fpu_mul_ctl/m2stg_ld0_2[1] , \fpu_mul_ctl/m2stg_ld0_1[5] ,
         \fpu_mul_ctl/m2stg_ld0_1[4] , \fpu_mul_ctl/m2stg_ld0_1[3] ,
         \fpu_mul_ctl/m2stg_ld0_1[2] , \fpu_mul_ctl/m2stg_ld0_1[1] ,
         \fpu_mul_ctl/mul_of_out_cout , \fpu_mul_ctl/mul_of_out_tmp2 ,
         \fpu_mul_ctl/m2stg_sign2 , \fpu_mul_ctl/m5stg_id[4] ,
         \fpu_mul_ctl/m5stg_rnd_mode[0] , \fpu_mul_ctl/m5stg_opdec[4] ,
         \fpu_mul_ctl/m4stg_id[4] , \fpu_mul_ctl/m4stg_rnd_mode[0] ,
         \fpu_mul_ctl/m3stg_id[4] , \fpu_mul_ctl/m3stg_rnd_mode[0] ,
         \fpu_mul_ctl/m3bstg_id[4] , \fpu_mul_ctl/m3bstg_rnd_mode[0] ,
         \fpu_mul_ctl/m3astg_id[4] , \fpu_mul_ctl/m3astg_rnd_mode[0] ,
         \fpu_mul_ctl/m2stg_id[4] , \fpu_mul_ctl/m2stg_rnd_mode[0] ,
         \fpu_mul_ctl/m2stg_zero_in , \fpu_mul_frac_dp/n838 ,
         \fpu_mul_frac_dp/n837 , \fpu_mul_frac_dp/n836 ,
         \fpu_mul_frac_dp/n834 , \fpu_mul_frac_dp/n833 ,
         \fpu_mul_frac_dp/n832 , \fpu_mul_frac_dp/n831 ,
         \fpu_mul_frac_dp/n829 , \fpu_mul_frac_dp/n828 ,
         \fpu_mul_frac_dp/n827 , \fpu_mul_frac_dp/n826 ,
         \fpu_mul_frac_dp/n825 , \fpu_mul_frac_dp/n824 ,
         \fpu_mul_frac_dp/n823 , \fpu_mul_frac_dp/n822 ,
         \fpu_mul_frac_dp/n821 , \fpu_mul_frac_dp/n820 ,
         \fpu_mul_frac_dp/n819 , \fpu_mul_frac_dp/n818 ,
         \fpu_mul_frac_dp/n817 , \fpu_mul_frac_dp/n816 ,
         \fpu_mul_frac_dp/n815 , \fpu_mul_frac_dp/n814 ,
         \fpu_mul_frac_dp/n813 , \fpu_mul_frac_dp/n812 ,
         \fpu_mul_frac_dp/n811 , \fpu_mul_frac_dp/n810 ,
         \fpu_mul_frac_dp/n809 , \fpu_mul_frac_dp/n808 ,
         \fpu_mul_frac_dp/n807 , \fpu_mul_frac_dp/n806 ,
         \fpu_mul_frac_dp/n805 , \fpu_mul_frac_dp/n804 ,
         \fpu_mul_frac_dp/n803 , \fpu_mul_frac_dp/n802 ,
         \fpu_mul_frac_dp/n801 , \fpu_mul_frac_dp/n800 ,
         \fpu_mul_frac_dp/n797 , \fpu_mul_frac_dp/n796 ,
         \fpu_mul_frac_dp/n795 , \fpu_mul_frac_dp/n794 ,
         \fpu_mul_frac_dp/n793 , \fpu_mul_frac_dp/n792 ,
         \fpu_mul_frac_dp/n791 , \fpu_mul_frac_dp/n790 ,
         \fpu_mul_frac_dp/n789 , \fpu_mul_frac_dp/n788 ,
         \fpu_mul_frac_dp/n787 , \fpu_mul_frac_dp/n786 ,
         \fpu_mul_frac_dp/n785 , \fpu_mul_frac_dp/n784 ,
         \fpu_mul_frac_dp/n783 , \fpu_mul_frac_dp/n782 ,
         \fpu_mul_frac_dp/n781 , \fpu_mul_frac_dp/n780 ,
         \fpu_mul_frac_dp/n779 , \fpu_mul_frac_dp/n778 ,
         \fpu_mul_frac_dp/n777 , \fpu_mul_frac_dp/n776 ,
         \fpu_mul_frac_dp/n775 , \fpu_mul_frac_dp/n767 ,
         \fpu_mul_frac_dp/n766 , \fpu_mul_frac_dp/n765 ,
         \fpu_mul_frac_dp/n764 , \fpu_mul_frac_dp/n763 ,
         \fpu_mul_frac_dp/n762 , \fpu_mul_frac_dp/n761 ,
         \fpu_mul_frac_dp/n760 , \fpu_mul_frac_dp/n759 ,
         \fpu_mul_frac_dp/n758 , \fpu_mul_frac_dp/n757 ,
         \fpu_mul_frac_dp/n756 , \fpu_mul_frac_dp/n754 ,
         \fpu_mul_frac_dp/n753 , \fpu_mul_frac_dp/n752 ,
         \fpu_mul_frac_dp/n751 , \fpu_mul_frac_dp/n750 ,
         \fpu_mul_frac_dp/n749 , \fpu_mul_frac_dp/n1097 ,
         \fpu_mul_frac_dp/n1096 , \fpu_mul_frac_dp/n1095 ,
         \fpu_mul_frac_dp/n1094 , \fpu_mul_frac_dp/n1093 ,
         \fpu_mul_frac_dp/n1092 , \fpu_mul_frac_dp/n1091 ,
         \fpu_mul_frac_dp/n1090 , \fpu_mul_frac_dp/n1089 ,
         \fpu_mul_frac_dp/n1088 , \fpu_mul_frac_dp/n1087 ,
         \fpu_mul_frac_dp/n1086 , \fpu_mul_frac_dp/n1085 ,
         \fpu_mul_frac_dp/n1084 , \fpu_mul_frac_dp/n1083 ,
         \fpu_mul_frac_dp/n1082 , \fpu_mul_frac_dp/n1081 ,
         \fpu_mul_frac_dp/n1080 , \fpu_mul_frac_dp/n1079 ,
         \fpu_mul_frac_dp/n1078 , \fpu_mul_frac_dp/n1077 ,
         \fpu_mul_frac_dp/n1076 , \fpu_mul_frac_dp/n1075 ,
         \fpu_mul_frac_dp/n1074 , \fpu_mul_frac_dp/n1073 ,
         \fpu_mul_frac_dp/n1072 , \fpu_mul_frac_dp/n1071 ,
         \fpu_mul_frac_dp/n1070 , \fpu_mul_frac_dp/n1069 ,
         \fpu_mul_frac_dp/n1068 , \fpu_mul_frac_dp/n1067 ,
         \fpu_mul_frac_dp/n1066 , \fpu_mul_frac_dp/n1065 ,
         \fpu_mul_frac_dp/n1064 , \fpu_mul_frac_dp/n1063 ,
         \fpu_mul_frac_dp/n1062 , \fpu_mul_frac_dp/n1061 ,
         \fpu_mul_frac_dp/n1060 , \fpu_mul_frac_dp/n1059 ,
         \fpu_mul_frac_dp/n1058 , \fpu_mul_frac_dp/n1057 ,
         \fpu_mul_frac_dp/n1056 , \fpu_mul_frac_dp/n1055 ,
         \fpu_mul_frac_dp/n1054 , \fpu_mul_frac_dp/n1053 ,
         \fpu_mul_frac_dp/n1052 , \fpu_mul_frac_dp/n1051 ,
         \fpu_mul_frac_dp/n1050 , \fpu_mul_frac_dp/n1049 ,
         \fpu_mul_frac_dp/n1048 , \fpu_mul_frac_dp/n1047 ,
         \fpu_mul_frac_dp/n1046 , \fpu_mul_frac_dp/n1045 ,
         \fpu_mul_frac_dp/n1044 , \fpu_mul_frac_dp/n1043 ,
         \fpu_mul_frac_dp/n1042 , \fpu_mul_frac_dp/n1041 ,
         \fpu_mul_frac_dp/n1040 , \fpu_mul_frac_dp/n1039 ,
         \fpu_mul_frac_dp/n1038 , \fpu_mul_frac_dp/n1037 ,
         \fpu_mul_frac_dp/n1036 , \fpu_mul_frac_dp/n1035 ,
         \fpu_mul_frac_dp/n1034 , \fpu_mul_frac_dp/n1033 ,
         \fpu_mul_frac_dp/n1032 , \fpu_mul_frac_dp/n1031 ,
         \fpu_mul_frac_dp/n1030 , \fpu_mul_frac_dp/n1029 ,
         \fpu_mul_frac_dp/n1028 , \fpu_mul_frac_dp/n1027 ,
         \fpu_mul_frac_dp/n1026 , \fpu_mul_frac_dp/n1025 ,
         \fpu_mul_frac_dp/n1024 , \fpu_mul_frac_dp/n1023 ,
         \fpu_mul_frac_dp/n1022 , \fpu_mul_frac_dp/n1021 ,
         \fpu_mul_frac_dp/n1020 , \fpu_mul_frac_dp/n1019 ,
         \fpu_mul_frac_dp/n1018 , \fpu_mul_frac_dp/n1017 ,
         \fpu_mul_frac_dp/n1016 , \fpu_mul_frac_dp/n1015 ,
         \fpu_mul_frac_dp/n1014 , \fpu_mul_frac_dp/n1013 ,
         \fpu_mul_frac_dp/n1012 , \fpu_mul_frac_dp/n1011 ,
         \fpu_mul_frac_dp/n1010 , \fpu_mul_frac_dp/n1009 ,
         \fpu_mul_frac_dp/n1008 , \fpu_mul_frac_dp/n1007 ,
         \fpu_mul_frac_dp/n1006 , \fpu_mul_frac_dp/n1005 ,
         \fpu_mul_frac_dp/n1004 , \fpu_mul_frac_dp/n1003 ,
         \fpu_mul_frac_dp/n1002 , \fpu_mul_frac_dp/n1001 ,
         \fpu_mul_frac_dp/n1000 , \fpu_mul_frac_dp/n999 ,
         \fpu_mul_frac_dp/n998 , \fpu_mul_frac_dp/n997 ,
         \fpu_mul_frac_dp/n996 , \fpu_mul_frac_dp/n995 ,
         \fpu_mul_frac_dp/n994 , \fpu_mul_frac_dp/n993 ,
         \fpu_mul_frac_dp/n992 , \fpu_mul_frac_dp/n991 ,
         \fpu_mul_frac_dp/n990 , \fpu_mul_frac_dp/n989 ,
         \fpu_mul_frac_dp/n988 , \fpu_mul_frac_dp/n987 ,
         \fpu_mul_frac_dp/n986 , \fpu_mul_frac_dp/n985 ,
         \fpu_mul_frac_dp/n984 , \fpu_mul_frac_dp/n983 ,
         \fpu_mul_frac_dp/n982 , \fpu_mul_frac_dp/n981 ,
         \fpu_mul_frac_dp/n980 , \fpu_mul_frac_dp/n979 ,
         \fpu_mul_frac_dp/n978 , \fpu_mul_frac_dp/n977 ,
         \fpu_mul_frac_dp/n976 , \fpu_mul_frac_dp/n975 ,
         \fpu_mul_frac_dp/n974 , \fpu_mul_frac_dp/n973 ,
         \fpu_mul_frac_dp/n972 , \fpu_mul_frac_dp/n971 ,
         \fpu_mul_frac_dp/n970 , \fpu_mul_frac_dp/n969 ,
         \fpu_mul_frac_dp/n968 , \fpu_mul_frac_dp/n967 ,
         \fpu_mul_frac_dp/n966 , \fpu_mul_frac_dp/n965 ,
         \fpu_mul_frac_dp/n964 , \fpu_mul_frac_dp/n963 ,
         \fpu_mul_frac_dp/n962 , \fpu_mul_frac_dp/n961 ,
         \fpu_mul_frac_dp/n960 , \fpu_mul_frac_dp/n959 ,
         \fpu_mul_frac_dp/n958 , \fpu_mul_frac_dp/n957 ,
         \fpu_mul_frac_dp/n956 , \fpu_mul_frac_dp/n955 ,
         \fpu_mul_frac_dp/n954 , \fpu_mul_frac_dp/n953 ,
         \fpu_mul_frac_dp/n952 , \fpu_mul_frac_dp/n951 ,
         \fpu_mul_frac_dp/n950 , \fpu_mul_frac_dp/n949 ,
         \fpu_mul_frac_dp/n948 , \fpu_mul_frac_dp/n947 ,
         \fpu_mul_frac_dp/n946 , \fpu_mul_frac_dp/n945 ,
         \fpu_mul_frac_dp/n944 , \fpu_mul_frac_dp/n943 ,
         \fpu_mul_frac_dp/n942 , \fpu_mul_frac_dp/n941 ,
         \fpu_mul_frac_dp/n940 , \fpu_mul_frac_dp/n939 ,
         \fpu_mul_frac_dp/n938 , \fpu_mul_frac_dp/n937 ,
         \fpu_mul_frac_dp/n936 , \fpu_mul_frac_dp/n935 ,
         \fpu_mul_frac_dp/n934 , \fpu_mul_frac_dp/n933 ,
         \fpu_mul_frac_dp/n932 , \fpu_mul_frac_dp/n931 ,
         \fpu_mul_frac_dp/n930 , \fpu_mul_frac_dp/n929 ,
         \fpu_mul_frac_dp/n928 , \fpu_mul_frac_dp/n927 ,
         \fpu_mul_frac_dp/n926 , \fpu_mul_frac_dp/n925 ,
         \fpu_mul_frac_dp/n924 , \fpu_mul_frac_dp/n923 ,
         \fpu_mul_frac_dp/n922 , \fpu_mul_frac_dp/n425 ,
         \fpu_mul_frac_dp/n383 , \fpu_mul_frac_dp/n382 ,
         \fpu_mul_frac_dp/n360 , \fpu_mul_frac_dp/n359 ,
         \fpu_mul_frac_dp/n358 , \fpu_mul_frac_dp/n357 ,
         \fpu_mul_frac_dp/n356 , \fpu_mul_frac_dp/n355 ,
         \fpu_mul_frac_dp/n354 , \fpu_mul_frac_dp/n353 ,
         \fpu_mul_frac_dp/n352 , \fpu_mul_frac_dp/n351 ,
         \fpu_mul_frac_dp/n350 , \fpu_mul_frac_dp/n349 ,
         \fpu_mul_frac_dp/n348 , \fpu_mul_frac_dp/n347 ,
         \fpu_mul_frac_dp/n346 , \fpu_mul_frac_dp/n345 ,
         \fpu_mul_frac_dp/n344 , \fpu_mul_frac_dp/n343 ,
         \fpu_mul_frac_dp/n342 , \fpu_mul_frac_dp/n341 ,
         \fpu_mul_frac_dp/n340 , \fpu_mul_frac_dp/n339 ,
         \fpu_mul_frac_dp/n338 , \fpu_mul_frac_dp/n337 ,
         \fpu_mul_frac_dp/n336 , \fpu_mul_frac_dp/n335 ,
         \fpu_mul_frac_dp/n334 , \fpu_mul_frac_dp/n311 ,
         \fpu_mul_frac_dp/n310 , \fpu_mul_frac_dp/n309 ,
         \fpu_mul_frac_dp/n307 , \fpu_mul_frac_dp/n306 ,
         \fpu_mul_frac_dp/n305 , \fpu_mul_frac_dp/n303 ,
         \fpu_mul_frac_dp/n300 , \fpu_mul_frac_dp/n289 ,
         \fpu_mul_frac_dp/n287 , \fpu_mul_frac_dp/n286 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N4 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N5 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N6 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N7 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N8 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N9 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N10 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N11 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N12 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N13 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N14 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N15 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N16 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N17 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N18 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N19 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N20 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N21 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N22 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N23 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N24 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N25 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N26 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N27 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N28 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N29 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N30 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N31 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N32 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N33 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N34 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N35 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N36 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N37 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N38 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N39 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N40 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N41 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N42 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N43 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N44 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N45 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N46 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N47 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N48 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N49 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N50 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N51 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N52 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N53 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N54 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N55 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N56 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre4/N57 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N3 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N4 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N5 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N6 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N7 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N8 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N9 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N10 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N11 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N12 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N13 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N14 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N15 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N16 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N17 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N18 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N19 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N20 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N21 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N22 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N23 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N24 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N25 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N26 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N27 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N28 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N29 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N30 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N31 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N32 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N33 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N34 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N35 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N36 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N37 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N38 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N39 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N40 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N41 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N42 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N43 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N44 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N45 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N46 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N47 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N48 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N49 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N50 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N51 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N52 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N53 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N54 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N55 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N56 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre3/N57 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N4 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N5 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N6 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N7 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N8 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N9 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N10 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N11 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N12 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N13 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N14 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N15 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N16 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N17 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N18 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N19 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N20 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N21 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N22 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N23 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N24 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N25 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N26 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N27 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N28 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N29 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N30 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N31 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N32 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N33 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N34 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N35 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N36 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N37 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N38 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N39 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N40 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N41 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N42 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N43 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N44 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N45 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N46 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N47 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N48 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N49 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N50 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N51 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N52 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N53 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N54 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N55 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N56 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre2/N57 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N3 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N4 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N5 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N6 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N7 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N8 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N9 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N10 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N11 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N12 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N13 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N14 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N15 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N16 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N17 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N18 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N19 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N20 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N21 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N22 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N23 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N24 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N25 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N26 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N27 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N28 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N29 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N30 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N31 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N32 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N33 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N34 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N35 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N36 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N37 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N38 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N39 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N40 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N41 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N42 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N43 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N44 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N45 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N46 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N47 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N48 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N49 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N50 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N51 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N52 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N53 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N54 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N55 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N56 ,
         \fpu_mul_frac_dp/i_m5stg_frac_pre1/N57 ,
         \fpu_mul_frac_dp/ckbuf_mul_frac_dp/N1 ,
         \fpu_mul_frac_dp/ckbuf_mul_frac_dp/clken ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[54] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[53] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[52] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[51] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[50] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[49] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[48] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[47] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[46] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[45] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[44] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[43] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[42] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[41] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[40] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[39] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[38] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[37] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[36] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[35] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[34] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[33] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[32] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[31] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[30] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[29] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[28] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[27] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[26] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[25] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[24] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[23] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[22] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[21] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[20] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[19] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[18] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[17] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[16] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[15] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[14] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[13] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[12] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[11] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[10] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[9] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[8] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[7] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[6] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[5] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[4] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[3] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[2] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[1] ,
         \fpu_mul_frac_dp/m5stg_frac_pre4[0] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[54] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[53] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[52] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[51] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[50] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[49] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[48] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[47] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[46] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[45] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[44] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[43] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[42] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[41] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[40] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[39] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[38] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[37] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[36] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[35] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[34] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[33] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[32] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[31] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[30] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[29] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[28] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[27] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[26] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[25] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[24] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[23] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[22] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[21] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[20] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[19] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[18] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[17] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[16] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[15] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[14] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[13] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[12] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[11] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[10] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[9] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[8] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[7] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[6] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[5] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[4] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[3] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[2] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[1] ,
         \fpu_mul_frac_dp/m5stg_frac_pre3[0] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[54] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[53] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[52] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[51] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[50] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[49] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[48] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[47] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[46] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[45] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[44] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[43] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[42] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[41] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[40] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[39] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[38] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[37] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[36] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[35] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[34] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[33] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[32] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[31] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[30] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[29] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[28] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[27] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[26] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[25] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[24] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[23] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[22] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[21] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[20] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[19] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[18] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[17] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[16] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[15] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[14] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[13] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[12] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[11] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[10] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[9] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[8] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[7] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[6] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[5] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[4] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[3] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[2] ,
         \fpu_mul_frac_dp/m5stg_frac_pre2[1] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[54] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[53] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[52] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[51] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[50] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[49] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[48] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[47] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[46] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[45] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[44] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[43] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[42] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[41] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[40] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[39] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[38] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[37] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[36] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[35] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[34] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[33] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[32] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[31] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[30] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[29] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[28] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[27] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[26] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[25] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[24] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[23] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[22] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[21] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[20] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[19] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[18] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[17] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[16] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[15] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[14] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[13] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[12] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[11] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[10] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[9] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[8] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[7] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[6] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[5] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[4] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[3] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[2] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[1] ,
         \fpu_mul_frac_dp/m5stg_frac_pre1[0] , \i_m4stg_frac/n1285 ,
         \i_m4stg_frac/n1283 , \i_m4stg_frac/n1281 , \i_m4stg_frac/n1277 ,
         \i_m4stg_frac/n854 , \i_m4stg_frac/n850 , \i_m4stg_frac/n637 ,
         \i_m4stg_frac/n635 , \i_m4stg_frac/n633 , \i_m4stg_frac/n631 ,
         \i_m4stg_frac/n629 , \i_m4stg_frac/n627 , \i_m4stg_frac/n625 ,
         \i_m4stg_frac/n623 , \i_m4stg_frac/n621 , \i_m4stg_frac/n619 ,
         \i_m4stg_frac/n617 , \i_m4stg_frac/n615 , \i_m4stg_frac/n613 ,
         \i_m4stg_frac/n611 , \i_m4stg_frac/n609 , \i_m4stg_frac/n607 ,
         \i_m4stg_frac/n605 , \i_m4stg_frac/n603 , \i_m4stg_frac/n601 ,
         \i_m4stg_frac/n599 , \i_m4stg_frac/n597 , \i_m4stg_frac/n595 ,
         \i_m4stg_frac/n593 , \i_m4stg_frac/n591 , \i_m4stg_frac/n589 ,
         \i_m4stg_frac/n587 , \i_m4stg_frac/n585 , \i_m4stg_frac/n583 ,
         \i_m4stg_frac/n581 , \i_m4stg_frac/n579 , \i_m4stg_frac/n577 ,
         \i_m4stg_frac/n575 , \i_m4stg_frac/n573 , \i_m4stg_frac/n571 ,
         \i_m4stg_frac/n569 , \i_m4stg_frac/n567 , \i_m4stg_frac/n565 ,
         \i_m4stg_frac/n563 , \i_m4stg_frac/n561 , \i_m4stg_frac/n559 ,
         \i_m4stg_frac/n557 , \i_m4stg_frac/n555 , \i_m4stg_frac/n553 ,
         \i_m4stg_frac/n551 , \i_m4stg_frac/n549 , \i_m4stg_frac/n547 ,
         \i_m4stg_frac/n545 , \i_m4stg_frac/n543 , \i_m4stg_frac/n541 ,
         \i_m4stg_frac/n539 , \i_m4stg_frac/n537 , \i_m4stg_frac/n535 ,
         \i_m4stg_frac/n533 , \i_m4stg_frac/n531 , \i_m4stg_frac/n529 ,
         \i_m4stg_frac/n527 , \i_m4stg_frac/n525 , \i_m4stg_frac/n523 ,
         \i_m4stg_frac/n521 , \i_m4stg_frac/n519 , \i_m4stg_frac/n517 ,
         \i_m4stg_frac/n515 , \i_m4stg_frac/n513 , \i_m4stg_frac/n511 ,
         \i_m4stg_frac/n509 , \i_m4stg_frac/n507 , \i_m4stg_frac/n505 ,
         \i_m4stg_frac/n503 , \i_m4stg_frac/n501 , \i_m4stg_frac/n499 ,
         \i_m4stg_frac/n497 , \i_m4stg_frac/n495 , \i_m4stg_frac/n493 ,
         \i_m4stg_frac/n492 , \i_m4stg_frac/n491 , \i_m4stg_frac/n489 ,
         \i_m4stg_frac/n487 , \i_m4stg_frac/n485 , \i_m4stg_frac/n483 ,
         \i_m4stg_frac/n481 , \i_m4stg_frac/n479 , \i_m4stg_frac/n477 ,
         \i_m4stg_frac/n475 , \i_m4stg_frac/n473 , \i_m4stg_frac/n471 ,
         \i_m4stg_frac/n469 , \i_m4stg_frac/n467 , \i_m4stg_frac/n465 ,
         \i_m4stg_frac/n463 , \i_m4stg_frac/n461 , \i_m4stg_frac/n459 ,
         \i_m4stg_frac/n457 , \i_m4stg_frac/n455 , \i_m4stg_frac/n453 ,
         \i_m4stg_frac/n451 , \i_m4stg_frac/n449 , \i_m4stg_frac/n447 ,
         \i_m4stg_frac/n445 , \i_m4stg_frac/n443 , \i_m4stg_frac/n441 ,
         \i_m4stg_frac/n439 , \i_m4stg_frac/n437 , \i_m4stg_frac/n435 ,
         \i_m4stg_frac/n433 , \i_m4stg_frac/n431 , \i_m4stg_frac/n429 ,
         \i_m4stg_frac/n427 , \i_m4stg_frac/n425 , \i_m4stg_frac/n423 ,
         \i_m4stg_frac/n421 , \i_m4stg_frac/n419 , \i_m4stg_frac/n417 ,
         \i_m4stg_frac/n415 , \i_m4stg_frac/n413 , \i_m4stg_frac/n411 ,
         \i_m4stg_frac/n409 , \i_m4stg_frac/n407 , \i_m4stg_frac/n405 ,
         \i_m4stg_frac/n403 , \i_m4stg_frac/n401 , \i_m4stg_frac/n399 ,
         \i_m4stg_frac/n397 , \i_m4stg_frac/n395 , \i_m4stg_frac/n393 ,
         \i_m4stg_frac/n391 , \i_m4stg_frac/n389 , \i_m4stg_frac/n387 ,
         \i_m4stg_frac/n385 , \i_m4stg_frac/n383 , \i_m4stg_frac/n381 ,
         \i_m4stg_frac/n379 , \i_m4stg_frac/n377 , \i_m4stg_frac/n375 ,
         \i_m4stg_frac/n373 , \i_m4stg_frac/n371 , \i_m4stg_frac/n369 ,
         \i_m4stg_frac/n367 , \i_m4stg_frac/n365 , \i_m4stg_frac/n363 ,
         \i_m4stg_frac/n361 , \i_m4stg_frac/n359 , \i_m4stg_frac/n357 ,
         \i_m4stg_frac/n355 , \i_m4stg_frac/n345 , \i_m4stg_frac/n343 ,
         \i_m4stg_frac/n341 , \i_m4stg_frac/n339 , \i_m4stg_frac/n337 ,
         \i_m4stg_frac/n336 , \i_m4stg_frac/n335 , \i_m4stg_frac/n334 ,
         \i_m4stg_frac/n333 , \i_m4stg_frac/n300 , \i_m4stg_frac/n215 ,
         \i_m4stg_frac/n213 , \i_m4stg_frac/n211 , \i_m4stg_frac/n209 ,
         \i_m4stg_frac/n207 , \i_m4stg_frac/n205 , \i_m4stg_frac/n203 ,
         \i_m4stg_frac/n201 , \i_m4stg_frac/n199 , \i_m4stg_frac/n1693 ,
         \i_m4stg_frac/n1692 , \i_m4stg_frac/n1684 , \i_m4stg_frac/n1532 ,
         \i_m4stg_frac/n1530 , \i_m4stg_frac/n1519 , \i_m4stg_frac/n1518 ,
         \i_m4stg_frac/n1517 , \i_m4stg_frac/n1516 , \i_m4stg_frac/n1515 ,
         \i_m4stg_frac/n1514 , \i_m4stg_frac/n1513 , \i_m4stg_frac/n1512 ,
         \i_m4stg_frac/n1511 , \i_m4stg_frac/n1510 , \i_m4stg_frac/n1509 ,
         \i_m4stg_frac/n1508 , \i_m4stg_frac/n1507 , \i_m4stg_frac/n1506 ,
         \i_m4stg_frac/n1505 , \i_m4stg_frac/n1504 , \i_m4stg_frac/n1503 ,
         \i_m4stg_frac/n1502 , \i_m4stg_frac/n1501 , \i_m4stg_frac/n1500 ,
         \i_m4stg_frac/n1499 , \i_m4stg_frac/n1498 , \i_m4stg_frac/n1497 ,
         \i_m4stg_frac/n1496 , \i_m4stg_frac/n1495 , \i_m4stg_frac/n1494 ,
         \i_m4stg_frac/n1493 , \i_m4stg_frac/n1492 , \i_m4stg_frac/n1491 ,
         \i_m4stg_frac/n1490 , \i_m4stg_frac/n1489 , \i_m4stg_frac/n1488 ,
         \i_m4stg_frac/n1487 , \i_m4stg_frac/n1486 , \i_m4stg_frac/n1485 ,
         \i_m4stg_frac/n1484 , \i_m4stg_frac/n1483 , \i_m4stg_frac/n1482 ,
         \i_m4stg_frac/n1481 , \i_m4stg_frac/n1480 , \i_m4stg_frac/n1479 ,
         \i_m4stg_frac/n1478 , \i_m4stg_frac/n1477 , \i_m4stg_frac/n1476 ,
         \i_m4stg_frac/n1475 , \i_m4stg_frac/n1474 , \i_m4stg_frac/n1473 ,
         \i_m4stg_frac/n1472 , \i_m4stg_frac/n1471 , \i_m4stg_frac/n1470 ,
         \i_m4stg_frac/n1469 , \i_m4stg_frac/n1468 , \i_m4stg_frac/n1467 ,
         \i_m4stg_frac/n1464 , \i_m4stg_frac/n1462 , \i_m4stg_frac/n1329 ,
         \i_m4stg_frac/n1056 , \i_m4stg_frac/n1055 , \i_m4stg_frac/n1021 ,
         \i_m4stg_frac/n1020 , \i_m4stg_frac/n1019 , \i_m4stg_frac/n1018 ,
         \i_m4stg_frac/n1017 , \i_m4stg_frac/n1016 , \i_m4stg_frac/n1015 ,
         \i_m4stg_frac/n1013 , \i_m4stg_frac/n1012 , \i_m4stg_frac/n1011 ,
         \i_m4stg_frac/n1010 , \i_m4stg_frac/n1009 , \i_m4stg_frac/n1008 ,
         \i_m4stg_frac/n1007 , \i_m4stg_frac/n1006 , \i_m4stg_frac/n1004 ,
         \i_m4stg_frac/n1003 , \i_m4stg_frac/n1002 , \i_m4stg_frac/n1001 ,
         \i_m4stg_frac/n1000 , \i_m4stg_frac/n999 , \i_m4stg_frac/n998 ,
         \i_m4stg_frac/n997 , \i_m4stg_frac/n989 , \i_m4stg_frac/n985 ,
         \i_m4stg_frac/n969 , \i_m4stg_frac/n965 , \i_m4stg_frac/n963 ,
         \i_m4stg_frac/n961 , \i_m4stg_frac/n959 , \i_m4stg_frac/n957 ,
         \i_m4stg_frac/n955 , \i_m4stg_frac/n953 , \i_m4stg_frac/n951 ,
         \i_m4stg_frac/n949 , \i_m4stg_frac/n947 , \i_m4stg_frac/n945 ,
         \i_m4stg_frac/n943 , \i_m4stg_frac/n941 , \i_m4stg_frac/n939 ,
         \i_m4stg_frac/n937 , \i_m4stg_frac/n935 , \i_m4stg_frac/n933 ,
         \i_m4stg_frac/n931 , \i_m4stg_frac/n929 , \i_m4stg_frac/n927 ,
         \i_m4stg_frac/n925 , \i_m4stg_frac/n923 , \i_m4stg_frac/n921 ,
         \i_m4stg_frac/n919 , \i_m4stg_frac/n917 , \i_m4stg_frac/n915 ,
         \i_m4stg_frac/n913 , \i_m4stg_frac/n911 , \i_m4stg_frac/n909 ,
         \i_m4stg_frac/n907 , \i_m4stg_frac/n905 , \i_m4stg_frac/n903 ,
         \i_m4stg_frac/n901 , \i_m4stg_frac/n899 , \i_m4stg_frac/n897 ,
         \i_m4stg_frac/n895 , \i_m4stg_frac/n893 , \i_m4stg_frac/n891 ,
         \i_m4stg_frac/n889 , \i_m4stg_frac/n887 , \i_m4stg_frac/n885 ,
         \i_m4stg_frac/n883 , \i_m4stg_frac/n881 , \i_m4stg_frac/n879 ,
         \i_m4stg_frac/n877 , \i_m4stg_frac/n875 , \i_m4stg_frac/n873 ,
         \i_m4stg_frac/n871 , \i_m4stg_frac/n869 , \i_m4stg_frac/n867 ,
         \i_m4stg_frac/n865 , \i_m4stg_frac/n863 , \i_m4stg_frac/n861 ,
         \i_m4stg_frac/n859 , \i_m4stg_frac/n857 , \i_m4stg_frac/n855 ,
         \i_m4stg_frac/n853 , \i_m4stg_frac/n851 , \i_m4stg_frac/n849 ,
         \i_m4stg_frac/n847 , \i_m4stg_frac/n845 , \i_m4stg_frac/n843 ,
         \i_m4stg_frac/n841 , \i_m4stg_frac/n839 , \i_m4stg_frac/n837 ,
         \i_m4stg_frac/n833 , \i_m4stg_frac/n831 , \i_m4stg_frac/n827 ,
         \i_m4stg_frac/n825 , \i_m4stg_frac/n823 , \i_m4stg_frac/n821 ,
         \i_m4stg_frac/n819 , \i_m4stg_frac/n817 , \i_m4stg_frac/n815 ,
         \i_m4stg_frac/n811 , \i_m4stg_frac/n809 , \i_m4stg_frac/n807 ,
         \i_m4stg_frac/n805 , \i_m4stg_frac/n803 , \i_m4stg_frac/n801 ,
         \i_m4stg_frac/n799 , \i_m4stg_frac/n797 , \i_m4stg_frac/n795 ,
         \i_m4stg_frac/n793 , \i_m4stg_frac/n791 , \i_m4stg_frac/n789 ,
         \i_m4stg_frac/n787 , \i_m4stg_frac/n785 , \i_m4stg_frac/n783 ,
         \i_m4stg_frac/n781 , \i_m4stg_frac/n779 , \i_m4stg_frac/n777 ,
         \i_m4stg_frac/n775 , \i_m4stg_frac/n773 , \i_m4stg_frac/n771 ,
         \i_m4stg_frac/n769 , \i_m4stg_frac/n767 , \i_m4stg_frac/n765 ,
         \i_m4stg_frac/n763 , \i_m4stg_frac/n761 , \i_m4stg_frac/n759 ,
         \i_m4stg_frac/n757 , \i_m4stg_frac/n755 , \i_m4stg_frac/n753 ,
         \i_m4stg_frac/n751 , \i_m4stg_frac/n749 , \i_m4stg_frac/n747 ,
         \i_m4stg_frac/n745 , \i_m4stg_frac/n743 , \i_m4stg_frac/n741 ,
         \i_m4stg_frac/n739 , \i_m4stg_frac/n737 , \i_m4stg_frac/n735 ,
         \i_m4stg_frac/n733 , \i_m4stg_frac/n731 , \i_m4stg_frac/n729 ,
         \i_m4stg_frac/n727 , \i_m4stg_frac/n725 , \i_m4stg_frac/n723 ,
         \i_m4stg_frac/n721 , \i_m4stg_frac/n719 , \i_m4stg_frac/n717 ,
         \i_m4stg_frac/n715 , \i_m4stg_frac/n713 , \i_m4stg_frac/n711 ,
         \i_m4stg_frac/n707 , \i_m4stg_frac/n705 , \i_m4stg_frac/n703 ,
         \i_m4stg_frac/n701 , \i_m4stg_frac/n699 , \i_m4stg_frac/n697 ,
         \i_m4stg_frac/n695 , \i_m4stg_frac/n693 , \i_m4stg_frac/n691 ,
         \i_m4stg_frac/n689 , \i_m4stg_frac/n687 , \i_m4stg_frac/n685 ,
         \i_m4stg_frac/n683 , \i_m4stg_frac/n677 , \i_m4stg_frac/n676 ,
         \i_m4stg_frac/n675 , \i_m4stg_frac/n674 , \i_m4stg_frac/n673 ,
         \i_m4stg_frac/n672 , \i_m4stg_frac/n671 , \i_m4stg_frac/n669 ,
         \i_m4stg_frac/n668 , \i_m4stg_frac/n667 , \i_m4stg_frac/n666 ,
         \i_m4stg_frac/n665 , \i_m4stg_frac/n664 , \i_m4stg_frac/n663 ,
         \i_m4stg_frac/n662 , \i_m4stg_frac/n660 , \i_m4stg_frac/n659 ,
         \i_m4stg_frac/n658 , \i_m4stg_frac/n657 , \i_m4stg_frac/n656 ,
         \i_m4stg_frac/n655 , \i_m4stg_frac/n654 , \i_m4stg_frac/n652 ,
         \i_m4stg_frac/n642 , \i_m4stg_frac/n550 , \i_m4stg_frac/n548 ,
         \i_m4stg_frac/n546 , \i_m4stg_frac/n544 , \i_m4stg_frac/n542 ,
         \i_m4stg_frac/n540 , \i_m4stg_frac/n538 , \i_m4stg_frac/n536 ,
         \i_m4stg_frac/n534 , \i_m4stg_frac/n532 , \i_m4stg_frac/n530 ,
         \i_m4stg_frac/n528 , \i_m4stg_frac/n526 , \i_m4stg_frac/n524 ,
         \i_m4stg_frac/n522 , \i_m4stg_frac/n520 , \i_m4stg_frac/n518 ,
         \i_m4stg_frac/n516 , \i_m4stg_frac/n514 , \i_m4stg_frac/n512 ,
         \i_m4stg_frac/n510 , \i_m4stg_frac/n508 , \i_m4stg_frac/n506 ,
         \i_m4stg_frac/n504 , \i_m4stg_frac/n502 , \i_m4stg_frac/n500 ,
         \i_m4stg_frac/n498 , \i_m4stg_frac/n496 , \i_m4stg_frac/n494 ,
         \i_m4stg_frac/n490 , \i_m4stg_frac/n488 , \i_m4stg_frac/n486 ,
         \i_m4stg_frac/n484 , \i_m4stg_frac/n482 , \i_m4stg_frac/n480 ,
         \i_m4stg_frac/n478 , \i_m4stg_frac/n476 , \i_m4stg_frac/n474 ,
         \i_m4stg_frac/n472 , \i_m4stg_frac/n470 , \i_m4stg_frac/n468 ,
         \i_m4stg_frac/n466 , \i_m4stg_frac/n464 , \i_m4stg_frac/n462 ,
         \i_m4stg_frac/n460 , \i_m4stg_frac/n458 , \i_m4stg_frac/n456 ,
         \i_m4stg_frac/n454 , \i_m4stg_frac/n452 , \i_m4stg_frac/n450 ,
         \i_m4stg_frac/n448 , \i_m4stg_frac/n446 , \i_m4stg_frac/n444 ,
         \i_m4stg_frac/n442 , \i_m4stg_frac/n440 , \i_m4stg_frac/n438 ,
         \i_m4stg_frac/n436 , \i_m4stg_frac/n434 , \i_m4stg_frac/n432 ,
         \i_m4stg_frac/n430 , \i_m4stg_frac/n428 , \i_m4stg_frac/n426 ,
         \i_m4stg_frac/n424 , \i_m4stg_frac/n422 , \i_m4stg_frac/n420 ,
         \i_m4stg_frac/n418 , \i_m4stg_frac/n416 , \i_m4stg_frac/n414 ,
         \i_m4stg_frac/n412 , \i_m4stg_frac/n410 , \i_m4stg_frac/n408 ,
         \i_m4stg_frac/n406 , \i_m4stg_frac/n404 , \i_m4stg_frac/n402 ,
         \i_m4stg_frac/n400 , \i_m4stg_frac/n398 , \i_m4stg_frac/n396 ,
         \i_m4stg_frac/n394 , \i_m4stg_frac/n392 , \i_m4stg_frac/n390 ,
         \i_m4stg_frac/n388 , \i_m4stg_frac/n386 , \i_m4stg_frac/n384 ,
         \i_m4stg_frac/n382 , \i_m4stg_frac/n380 , \i_m4stg_frac/n378 ,
         \i_m4stg_frac/n376 , \i_m4stg_frac/n374 , \i_m4stg_frac/n372 ,
         \i_m4stg_frac/n370 , \i_m4stg_frac/n368 , \i_m4stg_frac/n366 ,
         \i_m4stg_frac/n364 , \i_m4stg_frac/n362 , \i_m4stg_frac/n360 ,
         \i_m4stg_frac/n358 , \i_m4stg_frac/n356 , \i_m4stg_frac/n354 ,
         \i_m4stg_frac/n352 , \i_m4stg_frac/n350 , \i_m4stg_frac/n348 ,
         \i_m4stg_frac/n346 , \i_m4stg_frac/n344 , \i_m4stg_frac/n342 ,
         \i_m4stg_frac/n340 , \i_m4stg_frac/n338 , \i_m4stg_frac/n332 ,
         \i_m4stg_frac/n331 , \i_m4stg_frac/n329 , \i_m4stg_frac/n328 ,
         \i_m4stg_frac/n327 , \i_m4stg_frac/n326 , \i_m4stg_frac/n325 ,
         \i_m4stg_frac/n324 , \i_m4stg_frac/n323 , \i_m4stg_frac/n322 ,
         \i_m4stg_frac/n321 , \i_m4stg_frac/n320 , \i_m4stg_frac/n319 ,
         \i_m4stg_frac/n318 , \i_m4stg_frac/n317 , \i_m4stg_frac/n316 ,
         \i_m4stg_frac/n315 , \i_m4stg_frac/n314 , \i_m4stg_frac/n313 ,
         \i_m4stg_frac/n312 , \i_m4stg_frac/n311 , \i_m4stg_frac/n310 ,
         \i_m4stg_frac/n309 , \i_m4stg_frac/n308 , \i_m4stg_frac/n307 ,
         \i_m4stg_frac/n306 , \i_m4stg_frac/n305 , \i_m4stg_frac/n304 ,
         \i_m4stg_frac/n303 , \i_m4stg_frac/n302 , \i_m4stg_frac/n301 ,
         \i_m4stg_frac/n299 , \i_m4stg_frac/n297 , \i_m4stg_frac/n295 ,
         \i_m4stg_frac/n293 , \i_m4stg_frac/n291 , \i_m4stg_frac/n289 ,
         \i_m4stg_frac/n287 , \i_m4stg_frac/n285 , \i_m4stg_frac/n283 ,
         \i_m4stg_frac/n281 , \i_m4stg_frac/n279 , \i_m4stg_frac/n277 ,
         \i_m4stg_frac/n275 , \i_m4stg_frac/n273 , \i_m4stg_frac/n271 ,
         \i_m4stg_frac/n269 , \i_m4stg_frac/n267 , \i_m4stg_frac/n265 ,
         \i_m4stg_frac/n263 , \i_m4stg_frac/n261 , \i_m4stg_frac/n259 ,
         \i_m4stg_frac/n257 , \i_m4stg_frac/n255 , \i_m4stg_frac/n253 ,
         \i_m4stg_frac/n251 , \i_m4stg_frac/n249 , \i_m4stg_frac/n247 ,
         \i_m4stg_frac/n245 , \i_m4stg_frac/n243 , \i_m4stg_frac/n241 ,
         \i_m4stg_frac/n239 , \i_m4stg_frac/n237 , \i_m4stg_frac/n235 ,
         \i_m4stg_frac/n233 , \i_m4stg_frac/n231 , \i_m4stg_frac/n229 ,
         \i_m4stg_frac/n227 , \i_m4stg_frac/n225 , \i_m4stg_frac/n223 ,
         \i_m4stg_frac/n221 , \i_m4stg_frac/n219 , \i_m4stg_frac/n217 ,
         \i_m4stg_frac/n164 , \i_m4stg_frac/n163 , \i_m4stg_frac/n162 ,
         \i_m4stg_frac/n161 , \i_m4stg_frac/n160 , \i_m4stg_frac/n159 ,
         \i_m4stg_frac/n158 , \i_m4stg_frac/n157 , \i_m4stg_frac/n156 ,
         \i_m4stg_frac/n155 , \i_m4stg_frac/n154 , \i_m4stg_frac/n153 ,
         \i_m4stg_frac/n152 , \i_m4stg_frac/n150 , \i_m4stg_frac/n149 ,
         \i_m4stg_frac/n148 , \i_m4stg_frac/n147 , \i_m4stg_frac/n146 ,
         \i_m4stg_frac/n145 , \i_m4stg_frac/n144 , \i_m4stg_frac/n143 ,
         \i_m4stg_frac/n142 , \i_m4stg_frac/n141 , \i_m4stg_frac/n140 ,
         \i_m4stg_frac/n139 , \i_m4stg_frac/n138 , \i_m4stg_frac/n137 ,
         \i_m4stg_frac/n136 , \i_m4stg_frac/n134 , \i_m4stg_frac/n132 ,
         \i_m4stg_frac/n130 , \i_m4stg_frac/n128 , \i_m4stg_frac/n126 ,
         \i_m4stg_frac/n124 , \i_m4stg_frac/n122 , \i_m4stg_frac/n120 ,
         \i_m4stg_frac/n118 , \i_m4stg_frac/n116 , \i_m4stg_frac/n114 ,
         \i_m4stg_frac/n112 , \i_m4stg_frac/n110 , \i_m4stg_frac/n108 ,
         \i_m4stg_frac/n106 , \i_m4stg_frac/n104 , \i_m4stg_frac/n102 ,
         \i_m4stg_frac/n100 , \i_m4stg_frac/n98 , \i_m4stg_frac/n96 ,
         \i_m4stg_frac/n94 , \i_m4stg_frac/n92 , \i_m4stg_frac/n90 ,
         \i_m4stg_frac/n88 , \i_m4stg_frac/n86 , \i_m4stg_frac/n84 ,
         \i_m4stg_frac/n82 , \i_m4stg_frac/n80 , \i_m4stg_frac/n78 ,
         \i_m4stg_frac/n76 , \i_m4stg_frac/n74 , \i_m4stg_frac/n72 ,
         \i_m4stg_frac/n70 , \i_m4stg_frac/n68 , \i_m4stg_frac/n66 ,
         \i_m4stg_frac/n64 , \i_m4stg_frac/n62 , \i_m4stg_frac/n60 ,
         \i_m4stg_frac/n58 , \i_m4stg_frac/n56 , \i_m4stg_frac/n54 ,
         \i_m4stg_frac/n52 , \i_m4stg_frac/booth/out_dff15/N3 ,
         \i_m4stg_frac/booth/out_dff15/N4 , \i_m4stg_frac/booth/out_dff15/N5 ,
         \i_m4stg_frac/booth/out_dff14/N3 , \i_m4stg_frac/booth/out_dff14/N4 ,
         \i_m4stg_frac/booth/out_dff14/N5 , \i_m4stg_frac/booth/out_dff13/N3 ,
         \i_m4stg_frac/booth/out_dff13/N4 , \i_m4stg_frac/booth/out_dff13/N5 ,
         \i_m4stg_frac/booth/out_dff12/N3 , \i_m4stg_frac/booth/out_dff12/N4 ,
         \i_m4stg_frac/booth/out_dff12/N5 , \i_m4stg_frac/booth/out_dff11/N3 ,
         \i_m4stg_frac/booth/out_dff11/N4 , \i_m4stg_frac/booth/out_dff11/N5 ,
         \i_m4stg_frac/booth/out_dff10/N3 , \i_m4stg_frac/booth/out_dff10/N4 ,
         \i_m4stg_frac/booth/out_dff9/N3 , \i_m4stg_frac/booth/out_dff9/N4 ,
         \i_m4stg_frac/booth/out_dff9/N5 , \i_m4stg_frac/booth/out_dff8/N3 ,
         \i_m4stg_frac/booth/out_dff8/N4 , \i_m4stg_frac/booth/out_dff8/N5 ,
         \i_m4stg_frac/booth/out_dff7/N3 , \i_m4stg_frac/booth/out_dff7/N4 ,
         \i_m4stg_frac/booth/out_dff7/N5 , \i_m4stg_frac/booth/out_dff6/N3 ,
         \i_m4stg_frac/booth/out_dff6/N4 , \i_m4stg_frac/booth/out_dff6/N5 ,
         \i_m4stg_frac/booth/out_dff5/N3 , \i_m4stg_frac/booth/out_dff5/N4 ,
         \i_m4stg_frac/booth/out_dff5/N5 , \i_m4stg_frac/booth/out_dff4/N3 ,
         \i_m4stg_frac/booth/out_dff4/N4 , \i_m4stg_frac/booth/out_dff4/N5 ,
         \i_m4stg_frac/booth/out_dff3/N3 , \i_m4stg_frac/booth/out_dff3/N4 ,
         \i_m4stg_frac/booth/out_dff3/N5 , \i_m4stg_frac/booth/out_dff2/N3 ,
         \i_m4stg_frac/booth/out_dff2/N4 , \i_m4stg_frac/booth/out_dff2/N5 ,
         \i_m4stg_frac/booth/out_dff1/N3 , \i_m4stg_frac/booth/out_dff1/N4 ,
         \i_m4stg_frac/booth/out_dff0/N3 , \i_m4stg_frac/booth/ckbuf_1/clken ,
         \i_m4stg_frac/booth/ckbuf_0/clken , \i_m4stg_frac/co31_dff/N3 ,
         \i_m4stg_frac/pcout_dff/N4 , \i_m4stg_frac/pcout_dff/N5 ,
         \i_m4stg_frac/pcout_dff/N6 , \i_m4stg_frac/pcout_dff/N7 ,
         \i_m4stg_frac/pcout_dff/N8 , \i_m4stg_frac/pcout_dff/N9 ,
         \i_m4stg_frac/pcout_dff/N10 , \i_m4stg_frac/pcout_dff/N11 ,
         \i_m4stg_frac/pcout_dff/N12 , \i_m4stg_frac/pcout_dff/N13 ,
         \i_m4stg_frac/pcout_dff/N14 , \i_m4stg_frac/pcout_dff/N15 ,
         \i_m4stg_frac/pcout_dff/N16 , \i_m4stg_frac/pcout_dff/N17 ,
         \i_m4stg_frac/pcout_dff/N18 , \i_m4stg_frac/pcout_dff/N19 ,
         \i_m4stg_frac/pcout_dff/N20 , \i_m4stg_frac/pcout_dff/N21 ,
         \i_m4stg_frac/pcout_dff/N22 , \i_m4stg_frac/pcout_dff/N23 ,
         \i_m4stg_frac/pcout_dff/N24 , \i_m4stg_frac/pcout_dff/N25 ,
         \i_m4stg_frac/pcout_dff/N26 , \i_m4stg_frac/pcout_dff/N27 ,
         \i_m4stg_frac/pcout_dff/N28 , \i_m4stg_frac/pcout_dff/N29 ,
         \i_m4stg_frac/pcout_dff/N30 , \i_m4stg_frac/pcout_dff/N31 ,
         \i_m4stg_frac/pcout_dff/N32 , \i_m4stg_frac/pcout_dff/N33 ,
         \i_m4stg_frac/pcout_dff/N34 , \i_m4stg_frac/pcout_dff/N35 ,
         \i_m4stg_frac/pcout_dff/N36 , \i_m4stg_frac/pcout_dff/N37 ,
         \i_m4stg_frac/pcout_dff/N38 , \i_m4stg_frac/pcout_dff/N39 ,
         \i_m4stg_frac/pcout_dff/N40 , \i_m4stg_frac/pcout_dff/N41 ,
         \i_m4stg_frac/pcout_dff/N42 , \i_m4stg_frac/pcout_dff/N43 ,
         \i_m4stg_frac/pcout_dff/N44 , \i_m4stg_frac/pcout_dff/N45 ,
         \i_m4stg_frac/pcout_dff/N46 , \i_m4stg_frac/pcout_dff/N47 ,
         \i_m4stg_frac/pcout_dff/N48 , \i_m4stg_frac/pcout_dff/N49 ,
         \i_m4stg_frac/pcout_dff/N50 , \i_m4stg_frac/pcout_dff/N51 ,
         \i_m4stg_frac/pcout_dff/N52 , \i_m4stg_frac/pcout_dff/N53 ,
         \i_m4stg_frac/pcout_dff/N54 , \i_m4stg_frac/pcout_dff/N55 ,
         \i_m4stg_frac/pcout_dff/N56 , \i_m4stg_frac/pcout_dff/N57 ,
         \i_m4stg_frac/pcout_dff/N58 , \i_m4stg_frac/pcout_dff/N59 ,
         \i_m4stg_frac/pcout_dff/N60 , \i_m4stg_frac/pcout_dff/N61 ,
         \i_m4stg_frac/pcout_dff/N62 , \i_m4stg_frac/pcout_dff/N63 ,
         \i_m4stg_frac/pcout_dff/N64 , \i_m4stg_frac/pcout_dff/N65 ,
         \i_m4stg_frac/pcout_dff/N66 , \i_m4stg_frac/pcout_dff/N67 ,
         \i_m4stg_frac/pcout_dff/N68 , \i_m4stg_frac/pcout_dff/N69 ,
         \i_m4stg_frac/pcout_dff/N70 , \i_m4stg_frac/psum_dff/N4 ,
         \i_m4stg_frac/psum_dff/N5 , \i_m4stg_frac/psum_dff/N6 ,
         \i_m4stg_frac/psum_dff/N7 , \i_m4stg_frac/psum_dff/N8 ,
         \i_m4stg_frac/psum_dff/N9 , \i_m4stg_frac/psum_dff/N10 ,
         \i_m4stg_frac/psum_dff/N11 , \i_m4stg_frac/psum_dff/N12 ,
         \i_m4stg_frac/psum_dff/N13 , \i_m4stg_frac/psum_dff/N14 ,
         \i_m4stg_frac/psum_dff/N15 , \i_m4stg_frac/psum_dff/N16 ,
         \i_m4stg_frac/psum_dff/N17 , \i_m4stg_frac/psum_dff/N18 ,
         \i_m4stg_frac/psum_dff/N19 , \i_m4stg_frac/psum_dff/N20 ,
         \i_m4stg_frac/psum_dff/N21 , \i_m4stg_frac/psum_dff/N22 ,
         \i_m4stg_frac/psum_dff/N23 , \i_m4stg_frac/psum_dff/N24 ,
         \i_m4stg_frac/psum_dff/N25 , \i_m4stg_frac/psum_dff/N26 ,
         \i_m4stg_frac/psum_dff/N27 , \i_m4stg_frac/psum_dff/N28 ,
         \i_m4stg_frac/psum_dff/N29 , \i_m4stg_frac/psum_dff/N30 ,
         \i_m4stg_frac/psum_dff/N31 , \i_m4stg_frac/psum_dff/N32 ,
         \i_m4stg_frac/psum_dff/N33 , \i_m4stg_frac/psum_dff/N34 ,
         \i_m4stg_frac/psum_dff/N35 , \i_m4stg_frac/psum_dff/N36 ,
         \i_m4stg_frac/psum_dff/N37 , \i_m4stg_frac/psum_dff/N38 ,
         \i_m4stg_frac/psum_dff/N39 , \i_m4stg_frac/psum_dff/N40 ,
         \i_m4stg_frac/psum_dff/N41 , \i_m4stg_frac/psum_dff/N42 ,
         \i_m4stg_frac/psum_dff/N43 , \i_m4stg_frac/psum_dff/N44 ,
         \i_m4stg_frac/psum_dff/N45 , \i_m4stg_frac/psum_dff/N46 ,
         \i_m4stg_frac/psum_dff/N47 , \i_m4stg_frac/psum_dff/N48 ,
         \i_m4stg_frac/psum_dff/N49 , \i_m4stg_frac/psum_dff/N50 ,
         \i_m4stg_frac/psum_dff/N51 , \i_m4stg_frac/psum_dff/N52 ,
         \i_m4stg_frac/psum_dff/N53 , \i_m4stg_frac/psum_dff/N54 ,
         \i_m4stg_frac/psum_dff/N55 , \i_m4stg_frac/psum_dff/N56 ,
         \i_m4stg_frac/psum_dff/N57 , \i_m4stg_frac/psum_dff/N58 ,
         \i_m4stg_frac/psum_dff/N59 , \i_m4stg_frac/psum_dff/N60 ,
         \i_m4stg_frac/psum_dff/N61 , \i_m4stg_frac/psum_dff/N62 ,
         \i_m4stg_frac/psum_dff/N63 , \i_m4stg_frac/psum_dff/N64 ,
         \i_m4stg_frac/psum_dff/N65 , \i_m4stg_frac/psum_dff/N66 ,
         \i_m4stg_frac/psum_dff/N67 , \i_m4stg_frac/psum_dff/N68 ,
         \i_m4stg_frac/psum_dff/N69 , \i_m4stg_frac/psum_dff/N70 ,
         \i_m4stg_frac/a2cot_dff/N19 , \i_m4stg_frac/booth/b[50] ,
         \i_m4stg_frac/booth/b[48] , \i_m4stg_frac/booth/b[44] ,
         \i_m4stg_frac/booth/b[38] , \i_m4stg_frac/booth/b[36] ,
         \i_m4stg_frac/booth/b[34] , \i_m4stg_frac/booth/b[31] ,
         \i_m4stg_frac/booth/b0_in1[2] , \i_m4stg_frac/ckbuf_1/N1 ,
         \i_m4stg_frac/cyc3_dff/N7 , \i_m4stg_frac/cyc2_dff/N7 ,
         \i_m4stg_frac/cyc1_dff/N7 , \i_m4stg_frac/ckbuf_0/N1 ,
         \i_m4stg_frac/addout[73] , \i_m4stg_frac/addout[72] ,
         \i_m4stg_frac/addout[71] , \i_m4stg_frac/addout[70] ,
         \i_m4stg_frac/addout[69] , \i_m4stg_frac/addout[68] ,
         \i_m4stg_frac/addout[67] , \i_m4stg_frac/addout[66] ,
         \i_m4stg_frac/addout[65] , \i_m4stg_frac/addout[64] ,
         \i_m4stg_frac/addout[63] , \i_m4stg_frac/addout[62] ,
         \i_m4stg_frac/addout[61] , \i_m4stg_frac/addout[60] ,
         \i_m4stg_frac/addout[59] , \i_m4stg_frac/addout[58] ,
         \i_m4stg_frac/addout[57] , \i_m4stg_frac/addout[56] ,
         \i_m4stg_frac/addout[55] , \i_m4stg_frac/addout[54] ,
         \i_m4stg_frac/addout[53] , \i_m4stg_frac/addout[52] ,
         \i_m4stg_frac/addout[51] , \i_m4stg_frac/addout[50] ,
         \i_m4stg_frac/addout[49] , \i_m4stg_frac/addout[48] ,
         \i_m4stg_frac/addout[47] , \i_m4stg_frac/addout[46] ,
         \i_m4stg_frac/addout[45] , \i_m4stg_frac/addout[44] ,
         \i_m4stg_frac/addout[43] , \i_m4stg_frac/addout[42] ,
         \i_m4stg_frac/addout[41] , \i_m4stg_frac/addout[40] ,
         \i_m4stg_frac/addout[39] , \i_m4stg_frac/addout[38] ,
         \i_m4stg_frac/addout[37] , \i_m4stg_frac/addout[36] ,
         \i_m4stg_frac/addout[35] , \i_m4stg_frac/addout[34] ,
         \i_m4stg_frac/addout[33] , \i_m4stg_frac/addout[32] ,
         \i_m4stg_frac/addout[31] , \i_m4stg_frac/addout[30] ,
         \i_m4stg_frac/addout[29] , \i_m4stg_frac/addout[28] ,
         \i_m4stg_frac/addout[27] , \i_m4stg_frac/addout[26] ,
         \i_m4stg_frac/addout[25] , \i_m4stg_frac/addout[24] ,
         \i_m4stg_frac/addout[23] , \i_m4stg_frac/addout[22] ,
         \i_m4stg_frac/addout[21] , \i_m4stg_frac/addout[20] ,
         \i_m4stg_frac/addout[19] , \i_m4stg_frac/addout[18] ,
         \i_m4stg_frac/addout[17] , \i_m4stg_frac/addout[16] ,
         \i_m4stg_frac/addout[15] , \i_m4stg_frac/addout[14] ,
         \i_m4stg_frac/addout[13] , \i_m4stg_frac/addout[12] ,
         \i_m4stg_frac/addout[11] , \i_m4stg_frac/addout[10] ,
         \i_m4stg_frac/addout[9] , \i_m4stg_frac/addout[8] ,
         \i_m4stg_frac/addout[7] , \i_m4stg_frac/addout[6] ,
         \i_m4stg_frac/addout[5] , \i_m4stg_frac/addout[4] ,
         \i_m4stg_frac/addout[3] , \i_m4stg_frac/addout[2] ,
         \i_m4stg_frac/addout[1] , \i_m4stg_frac/addout[0] ,
         \i_m4stg_frac/addin_cin , \i_m4stg_frac/addin_sum[73] ,
         \i_m4stg_frac/addin_sum[72] , \i_m4stg_frac/addin_sum[71] ,
         \i_m4stg_frac/addin_sum[70] , \i_m4stg_frac/addin_sum[69] ,
         \i_m4stg_frac/addin_sum[68] , \i_m4stg_frac/addin_sum[67] ,
         \i_m4stg_frac/addin_sum[66] , \i_m4stg_frac/addin_sum[65] ,
         \i_m4stg_frac/addin_sum[64] , \i_m4stg_frac/addin_sum[63] ,
         \i_m4stg_frac/addin_sum[62] , \i_m4stg_frac/addin_sum[61] ,
         \i_m4stg_frac/addin_sum[60] , \i_m4stg_frac/addin_sum[59] ,
         \i_m4stg_frac/addin_sum[58] , \i_m4stg_frac/addin_sum[57] ,
         \i_m4stg_frac/addin_sum[56] , \i_m4stg_frac/addin_sum[55] ,
         \i_m4stg_frac/addin_sum[54] , \i_m4stg_frac/addin_sum[53] ,
         \i_m4stg_frac/addin_sum[52] , \i_m4stg_frac/addin_sum[51] ,
         \i_m4stg_frac/addin_sum[50] , \i_m4stg_frac/addin_sum[49] ,
         \i_m4stg_frac/addin_sum[48] , \i_m4stg_frac/addin_sum[47] ,
         \i_m4stg_frac/addin_sum[46] , \i_m4stg_frac/addin_sum[45] ,
         \i_m4stg_frac/addin_sum[44] , \i_m4stg_frac/addin_sum[43] ,
         \i_m4stg_frac/addin_sum[42] , \i_m4stg_frac/addin_sum[41] ,
         \i_m4stg_frac/addin_sum[40] , \i_m4stg_frac/addin_sum[39] ,
         \i_m4stg_frac/addin_sum[38] , \i_m4stg_frac/addin_sum[37] ,
         \i_m4stg_frac/addin_sum[36] , \i_m4stg_frac/addin_sum[35] ,
         \i_m4stg_frac/addin_sum[34] , \i_m4stg_frac/addin_sum[33] ,
         \i_m4stg_frac/addin_sum[32] , \i_m4stg_frac/addin_sum[31] ,
         \i_m4stg_frac/addin_sum[30] , \i_m4stg_frac/addin_sum[29] ,
         \i_m4stg_frac/addin_sum[28] , \i_m4stg_frac/addin_sum[27] ,
         \i_m4stg_frac/addin_sum[26] , \i_m4stg_frac/addin_sum[25] ,
         \i_m4stg_frac/addin_sum[24] , \i_m4stg_frac/addin_sum[23] ,
         \i_m4stg_frac/addin_sum[22] , \i_m4stg_frac/addin_sum[21] ,
         \i_m4stg_frac/addin_sum[20] , \i_m4stg_frac/addin_sum[19] ,
         \i_m4stg_frac/addin_sum[18] , \i_m4stg_frac/addin_sum[17] ,
         \i_m4stg_frac/addin_sum[16] , \i_m4stg_frac/addin_sum[15] ,
         \i_m4stg_frac/addin_sum[14] , \i_m4stg_frac/addin_sum[13] ,
         \i_m4stg_frac/addin_sum[12] , \i_m4stg_frac/addin_sum[11] ,
         \i_m4stg_frac/addin_sum[10] , \i_m4stg_frac/addin_sum[9] ,
         \i_m4stg_frac/addin_sum[8] , \i_m4stg_frac/addin_sum[7] ,
         \i_m4stg_frac/addin_sum[6] , \i_m4stg_frac/addin_sum[5] ,
         \i_m4stg_frac/addin_sum[4] , \i_m4stg_frac/addin_sum[3] ,
         \i_m4stg_frac/addin_sum[1] , \i_m4stg_frac/addin_sum[0] ,
         \i_m4stg_frac/addin_cout[72] , \i_m4stg_frac/addin_cout[71] ,
         \i_m4stg_frac/addin_cout[70] , \i_m4stg_frac/addin_cout[69] ,
         \i_m4stg_frac/addin_cout[68] , \i_m4stg_frac/addin_cout[67] ,
         \i_m4stg_frac/addin_cout[66] , \i_m4stg_frac/addin_cout[65] ,
         \i_m4stg_frac/addin_cout[64] , \i_m4stg_frac/addin_cout[63] ,
         \i_m4stg_frac/addin_cout[62] , \i_m4stg_frac/addin_cout[61] ,
         \i_m4stg_frac/addin_cout[60] , \i_m4stg_frac/addin_cout[59] ,
         \i_m4stg_frac/addin_cout[58] , \i_m4stg_frac/addin_cout[57] ,
         \i_m4stg_frac/addin_cout[56] , \i_m4stg_frac/addin_cout[55] ,
         \i_m4stg_frac/addin_cout[54] , \i_m4stg_frac/addin_cout[53] ,
         \i_m4stg_frac/addin_cout[52] , \i_m4stg_frac/addin_cout[51] ,
         \i_m4stg_frac/addin_cout[50] , \i_m4stg_frac/addin_cout[49] ,
         \i_m4stg_frac/addin_cout[48] , \i_m4stg_frac/addin_cout[47] ,
         \i_m4stg_frac/addin_cout[46] , \i_m4stg_frac/addin_cout[45] ,
         \i_m4stg_frac/addin_cout[44] , \i_m4stg_frac/addin_cout[43] ,
         \i_m4stg_frac/addin_cout[42] , \i_m4stg_frac/addin_cout[41] ,
         \i_m4stg_frac/addin_cout[40] , \i_m4stg_frac/addin_cout[39] ,
         \i_m4stg_frac/addin_cout[38] , \i_m4stg_frac/addin_cout[37] ,
         \i_m4stg_frac/addin_cout[36] , \i_m4stg_frac/addin_cout[35] ,
         \i_m4stg_frac/addin_cout[34] , \i_m4stg_frac/addin_cout[33] ,
         \i_m4stg_frac/addin_cout[32] , \i_m4stg_frac/addin_cout[31] ,
         \i_m4stg_frac/addin_cout[30] , \i_m4stg_frac/addin_cout[29] ,
         \i_m4stg_frac/addin_cout[28] , \i_m4stg_frac/addin_cout[27] ,
         \i_m4stg_frac/addin_cout[26] , \i_m4stg_frac/addin_cout[25] ,
         \i_m4stg_frac/addin_cout[24] , \i_m4stg_frac/addin_cout[23] ,
         \i_m4stg_frac/addin_cout[22] , \i_m4stg_frac/addin_cout[21] ,
         \i_m4stg_frac/addin_cout[20] , \i_m4stg_frac/addin_cout[19] ,
         \i_m4stg_frac/addin_cout[18] , \i_m4stg_frac/addin_cout[17] ,
         \i_m4stg_frac/addin_cout[16] , \i_m4stg_frac/addin_cout[14] ,
         \i_m4stg_frac/addin_cout[13] , \i_m4stg_frac/addin_cout[12] ,
         \i_m4stg_frac/addin_cout[11] , \i_m4stg_frac/addin_cout[10] ,
         \i_m4stg_frac/addin_cout[9] , \i_m4stg_frac/addin_cout[8] ,
         \i_m4stg_frac/addin_cout[7] , \i_m4stg_frac/addin_cout[6] ,
         \i_m4stg_frac/addin_cout[5] , \i_m4stg_frac/addin_cout[4] ,
         \i_m4stg_frac/addin_cout[3] , \i_m4stg_frac/addin_cout[2] ,
         \i_m4stg_frac/ps[98] , \i_m4stg_frac/ps[97] , \i_m4stg_frac/ps[96] ,
         \i_m4stg_frac/ps[95] , \i_m4stg_frac/ps[94] , \i_m4stg_frac/ps[93] ,
         \i_m4stg_frac/ps[92] , \i_m4stg_frac/ps[91] , \i_m4stg_frac/ps[90] ,
         \i_m4stg_frac/ps[89] , \i_m4stg_frac/ps[88] , \i_m4stg_frac/ps[87] ,
         \i_m4stg_frac/ps[86] , \i_m4stg_frac/ps[85] , \i_m4stg_frac/ps[84] ,
         \i_m4stg_frac/ps[83] , \i_m4stg_frac/ps[82] , \i_m4stg_frac/ps[81] ,
         \i_m4stg_frac/ps[80] , \i_m4stg_frac/ps[79] , \i_m4stg_frac/ps[78] ,
         \i_m4stg_frac/ps[77] , \i_m4stg_frac/ps[76] , \i_m4stg_frac/ps[75] ,
         \i_m4stg_frac/ps[74] , \i_m4stg_frac/ps[73] , \i_m4stg_frac/ps[72] ,
         \i_m4stg_frac/ps[71] , \i_m4stg_frac/ps[70] , \i_m4stg_frac/ps[69] ,
         \i_m4stg_frac/ps[68] , \i_m4stg_frac/ps[67] , \i_m4stg_frac/ps[66] ,
         \i_m4stg_frac/ps[65] , \i_m4stg_frac/ps[64] , \i_m4stg_frac/ps[63] ,
         \i_m4stg_frac/ps[62] , \i_m4stg_frac/ps[61] , \i_m4stg_frac/ps[60] ,
         \i_m4stg_frac/ps[59] , \i_m4stg_frac/ps[58] , \i_m4stg_frac/ps[57] ,
         \i_m4stg_frac/ps[56] , \i_m4stg_frac/ps[55] , \i_m4stg_frac/ps[54] ,
         \i_m4stg_frac/ps[53] , \i_m4stg_frac/ps[52] , \i_m4stg_frac/ps[51] ,
         \i_m4stg_frac/ps[50] , \i_m4stg_frac/ps[49] , \i_m4stg_frac/ps[48] ,
         \i_m4stg_frac/ps[47] , \i_m4stg_frac/ps[46] , \i_m4stg_frac/ps[45] ,
         \i_m4stg_frac/ps[44] , \i_m4stg_frac/ps[43] , \i_m4stg_frac/ps[42] ,
         \i_m4stg_frac/ps[41] , \i_m4stg_frac/ps[40] , \i_m4stg_frac/ps[39] ,
         \i_m4stg_frac/ps[38] , \i_m4stg_frac/ps[37] , \i_m4stg_frac/ps[36] ,
         \i_m4stg_frac/ps[35] , \i_m4stg_frac/ps[34] , \i_m4stg_frac/ps[33] ,
         \i_m4stg_frac/ps[32] , \i_m4stg_frac/pc[97] , \i_m4stg_frac/pc[96] ,
         \i_m4stg_frac/pc[95] , \i_m4stg_frac/pc[94] , \i_m4stg_frac/pc[93] ,
         \i_m4stg_frac/pc[92] , \i_m4stg_frac/pc[91] , \i_m4stg_frac/pc[90] ,
         \i_m4stg_frac/pc[89] , \i_m4stg_frac/pc[88] , \i_m4stg_frac/pc[87] ,
         \i_m4stg_frac/pc[86] , \i_m4stg_frac/pc[85] , \i_m4stg_frac/pc[84] ,
         \i_m4stg_frac/pc[83] , \i_m4stg_frac/pc[82] , \i_m4stg_frac/pc[81] ,
         \i_m4stg_frac/pc[80] , \i_m4stg_frac/pc[79] , \i_m4stg_frac/pc[78] ,
         \i_m4stg_frac/pc[77] , \i_m4stg_frac/pc[76] , \i_m4stg_frac/pc[75] ,
         \i_m4stg_frac/pc[74] , \i_m4stg_frac/pc[73] , \i_m4stg_frac/pc[72] ,
         \i_m4stg_frac/pc[71] , \i_m4stg_frac/pc[70] , \i_m4stg_frac/pc[69] ,
         \i_m4stg_frac/pc[68] , \i_m4stg_frac/pc[67] , \i_m4stg_frac/pc[66] ,
         \i_m4stg_frac/pc[65] , \i_m4stg_frac/pc[64] , \i_m4stg_frac/pc[63] ,
         \i_m4stg_frac/pc[62] , \i_m4stg_frac/pc[61] , \i_m4stg_frac/pc[60] ,
         \i_m4stg_frac/pc[59] , \i_m4stg_frac/pc[58] , \i_m4stg_frac/pc[57] ,
         \i_m4stg_frac/pc[56] , \i_m4stg_frac/pc[55] , \i_m4stg_frac/pc[54] ,
         \i_m4stg_frac/pc[53] , \i_m4stg_frac/pc[52] , \i_m4stg_frac/pc[51] ,
         \i_m4stg_frac/pc[50] , \i_m4stg_frac/pc[49] , \i_m4stg_frac/pc[48] ,
         \i_m4stg_frac/pc[47] , \i_m4stg_frac/pc[46] , \i_m4stg_frac/pc[45] ,
         \i_m4stg_frac/pc[44] , \i_m4stg_frac/pc[43] , \i_m4stg_frac/pc[42] ,
         \i_m4stg_frac/pc[41] , \i_m4stg_frac/pc[40] , \i_m4stg_frac/pc[39] ,
         \i_m4stg_frac/pc[38] , \i_m4stg_frac/pc[37] , \i_m4stg_frac/pc[36] ,
         \i_m4stg_frac/pc[35] , \i_m4stg_frac/pc[34] , \i_m4stg_frac/pc[33] ,
         \i_m4stg_frac/pc[32] , \i_m4stg_frac/pc[31] , \i_m4stg_frac/a1s[79] ,
         \i_m4stg_frac/a1s[78] , \i_m4stg_frac/a1s[77] ,
         \i_m4stg_frac/a1s[76] , \i_m4stg_frac/a1s[75] ,
         \i_m4stg_frac/a1s[74] , \i_m4stg_frac/a1s[73] ,
         \i_m4stg_frac/a1s[72] , \i_m4stg_frac/a1s[71] ,
         \i_m4stg_frac/a1s[70] , \i_m4stg_frac/a1s[69] ,
         \i_m4stg_frac/a1s[68] , \i_m4stg_frac/a1s[67] ,
         \i_m4stg_frac/a1s[66] , \i_m4stg_frac/a1s[65] ,
         \i_m4stg_frac/a1s[64] , \i_m4stg_frac/a1s[63] ,
         \i_m4stg_frac/a1s[62] , \i_m4stg_frac/a1s[61] ,
         \i_m4stg_frac/a1s[60] , \i_m4stg_frac/a1s[59] ,
         \i_m4stg_frac/a1s[58] , \i_m4stg_frac/a1s[57] ,
         \i_m4stg_frac/a1s[56] , \i_m4stg_frac/a1s[55] ,
         \i_m4stg_frac/a1s[54] , \i_m4stg_frac/a1s[53] ,
         \i_m4stg_frac/a1s[52] , \i_m4stg_frac/a1s[51] ,
         \i_m4stg_frac/a1c[79] , \i_m4stg_frac/a1c[78] ,
         \i_m4stg_frac/a1c[77] , \i_m4stg_frac/a1c[76] ,
         \i_m4stg_frac/a1c[75] , \i_m4stg_frac/a1c[74] ,
         \i_m4stg_frac/a1c[73] , \i_m4stg_frac/a1c[72] ,
         \i_m4stg_frac/a1c[71] , \i_m4stg_frac/a1c[70] ,
         \i_m4stg_frac/a1c[69] , \i_m4stg_frac/a1c[68] ,
         \i_m4stg_frac/a1c[67] , \i_m4stg_frac/a1c[66] ,
         \i_m4stg_frac/a1c[65] , \i_m4stg_frac/a1c[64] ,
         \i_m4stg_frac/a1c[63] , \i_m4stg_frac/a1c[62] ,
         \i_m4stg_frac/a1c[61] , \i_m4stg_frac/a1c[60] ,
         \i_m4stg_frac/a1c[59] , \i_m4stg_frac/a1c[58] ,
         \i_m4stg_frac/a1c[57] , \i_m4stg_frac/a1c[56] ,
         \i_m4stg_frac/a1c[55] , \i_m4stg_frac/a1c[54] ,
         \i_m4stg_frac/a1c[53] , \i_m4stg_frac/a1c[52] ,
         \i_m4stg_frac/a1c[51] , \i_m4stg_frac/a1c[50] ,
         \i_m4stg_frac/a1c[49] , \i_m4stg_frac/a1c[48] ,
         \i_m4stg_frac/a1c[47] , \i_m4stg_frac/a1c[46] ,
         \i_m4stg_frac/a1c[45] , \i_m4stg_frac/a1c[44] ,
         \i_m4stg_frac/a1c[43] , \i_m4stg_frac/a1c[42] ,
         \i_m4stg_frac/a1c[41] , \i_m4stg_frac/a1c[40] ,
         \i_m4stg_frac/a1c[39] , \i_m4stg_frac/a1c[38] ,
         \i_m4stg_frac/a1c[37] , \i_m4stg_frac/a1c[36] ,
         \i_m4stg_frac/a1c[35] , \i_m4stg_frac/a1c[34] ,
         \i_m4stg_frac/a1c[33] , \i_m4stg_frac/a1c[32] ,
         \i_m4stg_frac/a1c[31] , \i_m4stg_frac/a1c[30] ,
         \i_m4stg_frac/a1c[29] , \i_m4stg_frac/a1c[28] ,
         \i_m4stg_frac/a1c[27] , \i_m4stg_frac/a1c[26] ,
         \i_m4stg_frac/a1c[25] , \i_m4stg_frac/a1c[24] ,
         \i_m4stg_frac/a1c[23] , \i_m4stg_frac/a1c[22] ,
         \i_m4stg_frac/a1c[21] , \i_m4stg_frac/a1c[20] ,
         \i_m4stg_frac/a1c[19] , \i_m4stg_frac/a1c[18] ,
         \i_m4stg_frac/a1c[17] , \i_m4stg_frac/a1c[16] ,
         \i_m4stg_frac/a1c[15] , \i_m4stg_frac/a1c[14] ,
         \i_m4stg_frac/a1c[13] , \i_m4stg_frac/a1c[12] ,
         \i_m4stg_frac/a1c[11] , \i_m4stg_frac/a1c[10] , \i_m4stg_frac/a1c[9] ,
         \i_m4stg_frac/a1c[8] , \i_m4stg_frac/a1c[7] , \i_m4stg_frac/a1c[6] ,
         \i_m4stg_frac/a1c[5] , \i_m4stg_frac/a1c[4] ,
         \i_m4stg_frac/a1sum[81] , \i_m4stg_frac/a1sum[79] ,
         \i_m4stg_frac/a1sum[78] , \i_m4stg_frac/a1sum[77] ,
         \i_m4stg_frac/a1sum[76] , \i_m4stg_frac/a1sum[75] ,
         \i_m4stg_frac/a1sum[74] , \i_m4stg_frac/a1sum[73] ,
         \i_m4stg_frac/a1sum[72] , \i_m4stg_frac/a1sum[71] ,
         \i_m4stg_frac/a1sum[70] , \i_m4stg_frac/a1sum[69] ,
         \i_m4stg_frac/a1sum[68] , \i_m4stg_frac/a1sum[67] ,
         \i_m4stg_frac/a1sum[66] , \i_m4stg_frac/a1sum[65] ,
         \i_m4stg_frac/a1sum[64] , \i_m4stg_frac/a1sum[63] ,
         \i_m4stg_frac/a1sum[62] , \i_m4stg_frac/a1sum[61] ,
         \i_m4stg_frac/a1sum[60] , \i_m4stg_frac/a1sum[59] ,
         \i_m4stg_frac/a1sum[58] , \i_m4stg_frac/a1sum[57] ,
         \i_m4stg_frac/a1sum[56] , \i_m4stg_frac/a1sum[55] ,
         \i_m4stg_frac/a1sum[54] , \i_m4stg_frac/a1sum[53] ,
         \i_m4stg_frac/a1sum[52] , \i_m4stg_frac/a1sum[51] ,
         \i_m4stg_frac/a1sum[50] , \i_m4stg_frac/a1sum[49] ,
         \i_m4stg_frac/a1sum[48] , \i_m4stg_frac/a1sum[47] ,
         \i_m4stg_frac/a1sum[46] , \i_m4stg_frac/a1sum[45] ,
         \i_m4stg_frac/a1sum[44] , \i_m4stg_frac/a1sum[43] ,
         \i_m4stg_frac/a1sum[42] , \i_m4stg_frac/a1sum[41] ,
         \i_m4stg_frac/a1sum[40] , \i_m4stg_frac/a1sum[39] ,
         \i_m4stg_frac/a1sum[38] , \i_m4stg_frac/a1sum[37] ,
         \i_m4stg_frac/a1sum[36] , \i_m4stg_frac/a1sum[35] ,
         \i_m4stg_frac/a1sum[34] , \i_m4stg_frac/a1sum[33] ,
         \i_m4stg_frac/a1sum[32] , \i_m4stg_frac/a1sum[31] ,
         \i_m4stg_frac/a1sum[30] , \i_m4stg_frac/a1sum[29] ,
         \i_m4stg_frac/a1sum[28] , \i_m4stg_frac/a1sum[27] ,
         \i_m4stg_frac/a1sum[26] , \i_m4stg_frac/a1sum[25] ,
         \i_m4stg_frac/a1sum[24] , \i_m4stg_frac/a1sum[23] ,
         \i_m4stg_frac/a1sum[22] , \i_m4stg_frac/a1sum[21] ,
         \i_m4stg_frac/a1sum[20] , \i_m4stg_frac/a1sum[19] ,
         \i_m4stg_frac/a1sum[18] , \i_m4stg_frac/a1sum[17] ,
         \i_m4stg_frac/a1sum[16] , \i_m4stg_frac/a1sum[15] ,
         \i_m4stg_frac/a1sum[14] , \i_m4stg_frac/a1sum[13] ,
         \i_m4stg_frac/a1sum[12] , \i_m4stg_frac/a1sum[11] ,
         \i_m4stg_frac/a1sum[10] , \i_m4stg_frac/a1sum[9] ,
         \i_m4stg_frac/a1sum[8] , \i_m4stg_frac/a1sum[7] ,
         \i_m4stg_frac/a1sum[6] , \i_m4stg_frac/a1sum[5] ,
         \i_m4stg_frac/a1sum[4] , \i_m4stg_frac/a1sum[3] ,
         \i_m4stg_frac/a1sum[2] , \i_m4stg_frac/a1sum[1] ,
         \i_m4stg_frac/a1sum[0] , \i_m4stg_frac/a1cout[79] ,
         \i_m4stg_frac/a1cout[78] , \i_m4stg_frac/a1cout[77] ,
         \i_m4stg_frac/a1cout[76] , \i_m4stg_frac/a1cout[75] ,
         \i_m4stg_frac/a1cout[74] , \i_m4stg_frac/a1cout[73] ,
         \i_m4stg_frac/a1cout[72] , \i_m4stg_frac/a1cout[71] ,
         \i_m4stg_frac/a1cout[70] , \i_m4stg_frac/a1cout[69] ,
         \i_m4stg_frac/a1cout[68] , \i_m4stg_frac/a1cout[67] ,
         \i_m4stg_frac/a1cout[66] , \i_m4stg_frac/a1cout[65] ,
         \i_m4stg_frac/a1cout[64] , \i_m4stg_frac/a1cout[63] ,
         \i_m4stg_frac/a1cout[62] , \i_m4stg_frac/a1cout[61] ,
         \i_m4stg_frac/a1cout[60] , \i_m4stg_frac/a1cout[59] ,
         \i_m4stg_frac/a1cout[58] , \i_m4stg_frac/a1cout[57] ,
         \i_m4stg_frac/a1cout[56] , \i_m4stg_frac/a1cout[55] ,
         \i_m4stg_frac/a1cout[54] , \i_m4stg_frac/a1cout[53] ,
         \i_m4stg_frac/a1cout[52] , \i_m4stg_frac/a1cout[51] ,
         \i_m4stg_frac/a1cout[50] , \i_m4stg_frac/a1cout[49] ,
         \i_m4stg_frac/a1cout[48] , \i_m4stg_frac/a1cout[47] ,
         \i_m4stg_frac/a1cout[46] , \i_m4stg_frac/a1cout[45] ,
         \i_m4stg_frac/a1cout[44] , \i_m4stg_frac/a1cout[43] ,
         \i_m4stg_frac/a1cout[42] , \i_m4stg_frac/a1cout[41] ,
         \i_m4stg_frac/a1cout[40] , \i_m4stg_frac/a1cout[39] ,
         \i_m4stg_frac/a1cout[38] , \i_m4stg_frac/a1cout[37] ,
         \i_m4stg_frac/a1cout[36] , \i_m4stg_frac/a1cout[35] ,
         \i_m4stg_frac/a1cout[34] , \i_m4stg_frac/a1cout[33] ,
         \i_m4stg_frac/a1cout[32] , \i_m4stg_frac/a1cout[31] ,
         \i_m4stg_frac/a1cout[30] , \i_m4stg_frac/a1cout[29] ,
         \i_m4stg_frac/a1cout[28] , \i_m4stg_frac/a1cout[27] ,
         \i_m4stg_frac/a1cout[26] , \i_m4stg_frac/a1cout[25] ,
         \i_m4stg_frac/a1cout[24] , \i_m4stg_frac/a1cout[23] ,
         \i_m4stg_frac/a1cout[22] , \i_m4stg_frac/a1cout[21] ,
         \i_m4stg_frac/a1cout[20] , \i_m4stg_frac/a1cout[19] ,
         \i_m4stg_frac/a1cout[18] , \i_m4stg_frac/a1cout[17] ,
         \i_m4stg_frac/a1cout[16] , \i_m4stg_frac/a1cout[15] ,
         \i_m4stg_frac/a1cout[14] , \i_m4stg_frac/a1cout[13] ,
         \i_m4stg_frac/a1cout[12] , \i_m4stg_frac/a1cout[11] ,
         \i_m4stg_frac/a1cout[10] , \i_m4stg_frac/a1cout[9] ,
         \i_m4stg_frac/a1cout[8] , \i_m4stg_frac/a1cout[7] ,
         \i_m4stg_frac/a1cout[6] , \i_m4stg_frac/a1cout[5] ,
         \i_m4stg_frac/a1cout[4] , \i_m4stg_frac/a0s[16] ,
         \i_m4stg_frac/a0s[17] , \i_m4stg_frac/a0s[18] ,
         \i_m4stg_frac/a0s[19] , \i_m4stg_frac/a0s[20] ,
         \i_m4stg_frac/a0s[21] , \i_m4stg_frac/a0s[22] ,
         \i_m4stg_frac/a0s[23] , \i_m4stg_frac/a0s[24] ,
         \i_m4stg_frac/a0s[25] , \i_m4stg_frac/a0s[26] ,
         \i_m4stg_frac/a0s[27] , \i_m4stg_frac/a0s[28] ,
         \i_m4stg_frac/a0s[29] , \i_m4stg_frac/a0s[30] ,
         \i_m4stg_frac/a0s[31] , \i_m4stg_frac/a0s[32] ,
         \i_m4stg_frac/a0s[33] , \i_m4stg_frac/a0s[34] ,
         \i_m4stg_frac/a0s[35] , \i_m4stg_frac/a0s[36] ,
         \i_m4stg_frac/a0s[37] , \i_m4stg_frac/a0s[38] ,
         \i_m4stg_frac/a0s[39] , \i_m4stg_frac/a0s[40] ,
         \i_m4stg_frac/a0s[41] , \i_m4stg_frac/a0s[42] ,
         \i_m4stg_frac/a0s[43] , \i_m4stg_frac/a0s[44] ,
         \i_m4stg_frac/a0s[45] , \i_m4stg_frac/a0s[46] ,
         \i_m4stg_frac/a0s[47] , \i_m4stg_frac/a0s[48] ,
         \i_m4stg_frac/a0s[49] , \i_m4stg_frac/a0s[50] ,
         \i_m4stg_frac/a0s[51] , \i_m4stg_frac/a0s[52] ,
         \i_m4stg_frac/a0s[53] , \i_m4stg_frac/a0s[54] ,
         \i_m4stg_frac/a0s[55] , \i_m4stg_frac/a0s[56] ,
         \i_m4stg_frac/a0s[57] , \i_m4stg_frac/a0s[58] ,
         \i_m4stg_frac/a0s[59] , \i_m4stg_frac/a0s[60] ,
         \i_m4stg_frac/a0s[61] , \i_m4stg_frac/a0s[62] ,
         \i_m4stg_frac/a0s[63] , \i_m4stg_frac/a0s[64] ,
         \i_m4stg_frac/a0s[65] , \i_m4stg_frac/a0s[66] ,
         \i_m4stg_frac/a0s[68] , \i_m4stg_frac/a0s[69] ,
         \i_m4stg_frac/a0s[70] , \i_m4stg_frac/a0s[71] ,
         \i_m4stg_frac/a0s[72] , \i_m4stg_frac/a0s[73] ,
         \i_m4stg_frac/a0s[74] , \i_m4stg_frac/a0s[75] ,
         \i_m4stg_frac/a0s[76] , \i_m4stg_frac/a0s[77] ,
         \i_m4stg_frac/a0s[78] , \i_m4stg_frac/a0s[79] ,
         \i_m4stg_frac/a0s[80] , \i_m4stg_frac/a0c[79] ,
         \i_m4stg_frac/a0c[78] , \i_m4stg_frac/a0c[77] ,
         \i_m4stg_frac/a0c[76] , \i_m4stg_frac/a0c[75] ,
         \i_m4stg_frac/a0c[74] , \i_m4stg_frac/a0c[73] ,
         \i_m4stg_frac/a0c[72] , \i_m4stg_frac/a0c[71] ,
         \i_m4stg_frac/a0c[70] , \i_m4stg_frac/a0c[69] ,
         \i_m4stg_frac/a0c[68] , \i_m4stg_frac/a0c[67] ,
         \i_m4stg_frac/a0c[65] , \i_m4stg_frac/a0c[64] ,
         \i_m4stg_frac/a0c[63] , \i_m4stg_frac/a0c[62] ,
         \i_m4stg_frac/a0c[61] , \i_m4stg_frac/a0c[60] ,
         \i_m4stg_frac/a0c[59] , \i_m4stg_frac/a0c[58] ,
         \i_m4stg_frac/a0c[57] , \i_m4stg_frac/a0c[56] ,
         \i_m4stg_frac/a0c[55] , \i_m4stg_frac/a0c[54] ,
         \i_m4stg_frac/a0c[53] , \i_m4stg_frac/a0c[52] ,
         \i_m4stg_frac/a0c[51] , \i_m4stg_frac/a0c[50] ,
         \i_m4stg_frac/a0c[49] , \i_m4stg_frac/a0c[48] ,
         \i_m4stg_frac/a0c[47] , \i_m4stg_frac/a0c[46] ,
         \i_m4stg_frac/a0c[45] , \i_m4stg_frac/a0c[44] ,
         \i_m4stg_frac/a0c[43] , \i_m4stg_frac/a0c[42] ,
         \i_m4stg_frac/a0c[41] , \i_m4stg_frac/a0c[40] ,
         \i_m4stg_frac/a0c[39] , \i_m4stg_frac/a0c[38] ,
         \i_m4stg_frac/a0c[37] , \i_m4stg_frac/a0c[36] ,
         \i_m4stg_frac/a0c[35] , \i_m4stg_frac/a0c[34] ,
         \i_m4stg_frac/a0c[33] , \i_m4stg_frac/a0c[32] ,
         \i_m4stg_frac/a0c[31] , \i_m4stg_frac/a0c[30] ,
         \i_m4stg_frac/a0c[29] , \i_m4stg_frac/a0c[28] ,
         \i_m4stg_frac/a0c[27] , \i_m4stg_frac/a0c[26] ,
         \i_m4stg_frac/a0c[25] , \i_m4stg_frac/a0c[24] ,
         \i_m4stg_frac/a0c[23] , \i_m4stg_frac/a0c[22] ,
         \i_m4stg_frac/a0c[21] , \i_m4stg_frac/a0c[20] ,
         \i_m4stg_frac/a0c[19] , \i_m4stg_frac/a0c[18] ,
         \i_m4stg_frac/a0c[17] , \i_m4stg_frac/a0c[16] ,
         \i_m4stg_frac/a0c[15] , \i_m4stg_frac/a0c[12] ,
         \i_m4stg_frac/a0c[11] , \i_m4stg_frac/a0c[10] , \i_m4stg_frac/a0c[9] ,
         \i_m4stg_frac/a0c[8] , \i_m4stg_frac/a0c[7] , \i_m4stg_frac/a0c[4] ,
         \i_m4stg_frac/a0sum[79] , \i_m4stg_frac/a0sum[78] ,
         \i_m4stg_frac/a0sum[77] , \i_m4stg_frac/a0sum[76] ,
         \i_m4stg_frac/a0sum[75] , \i_m4stg_frac/a0sum[74] ,
         \i_m4stg_frac/a0sum[73] , \i_m4stg_frac/a0sum[72] ,
         \i_m4stg_frac/a0sum[71] , \i_m4stg_frac/a0sum[70] ,
         \i_m4stg_frac/a0sum[69] , \i_m4stg_frac/a0sum[68] ,
         \i_m4stg_frac/a0sum[67] , \i_m4stg_frac/a0sum[66] ,
         \i_m4stg_frac/a0sum[65] , \i_m4stg_frac/a0sum[64] ,
         \i_m4stg_frac/a0sum[63] , \i_m4stg_frac/a0sum[62] ,
         \i_m4stg_frac/a0sum[61] , \i_m4stg_frac/a0sum[60] ,
         \i_m4stg_frac/a0sum[59] , \i_m4stg_frac/a0sum[58] ,
         \i_m4stg_frac/a0sum[57] , \i_m4stg_frac/a0sum[56] ,
         \i_m4stg_frac/a0sum[55] , \i_m4stg_frac/a0sum[54] ,
         \i_m4stg_frac/a0sum[53] , \i_m4stg_frac/a0sum[52] ,
         \i_m4stg_frac/a0sum[51] , \i_m4stg_frac/a0sum[50] ,
         \i_m4stg_frac/a0sum[49] , \i_m4stg_frac/a0sum[48] ,
         \i_m4stg_frac/a0sum[47] , \i_m4stg_frac/a0sum[46] ,
         \i_m4stg_frac/a0sum[45] , \i_m4stg_frac/a0sum[44] ,
         \i_m4stg_frac/a0sum[43] , \i_m4stg_frac/a0sum[42] ,
         \i_m4stg_frac/a0sum[41] , \i_m4stg_frac/a0sum[40] ,
         \i_m4stg_frac/a0sum[39] , \i_m4stg_frac/a0sum[38] ,
         \i_m4stg_frac/a0sum[37] , \i_m4stg_frac/a0sum[36] ,
         \i_m4stg_frac/a0sum[35] , \i_m4stg_frac/a0sum[34] ,
         \i_m4stg_frac/a0sum[33] , \i_m4stg_frac/a0sum[32] ,
         \i_m4stg_frac/a0sum[31] , \i_m4stg_frac/a0sum[30] ,
         \i_m4stg_frac/a0sum[29] , \i_m4stg_frac/a0sum[28] ,
         \i_m4stg_frac/a0sum[27] , \i_m4stg_frac/a0sum[26] ,
         \i_m4stg_frac/a0sum[25] , \i_m4stg_frac/a0sum[24] ,
         \i_m4stg_frac/a0sum[23] , \i_m4stg_frac/a0sum[22] ,
         \i_m4stg_frac/a0sum[21] , \i_m4stg_frac/a0sum[20] ,
         \i_m4stg_frac/a0sum[19] , \i_m4stg_frac/a0sum[18] ,
         \i_m4stg_frac/a0sum[17] , \i_m4stg_frac/a0sum[16] ,
         \i_m4stg_frac/a0sum[15] , \i_m4stg_frac/a0sum[14] ,
         \i_m4stg_frac/a0sum[13] , \i_m4stg_frac/a0sum[12] ,
         \i_m4stg_frac/a0sum[11] , \i_m4stg_frac/a0sum[10] ,
         \i_m4stg_frac/a0sum[9] , \i_m4stg_frac/a0sum[8] ,
         \i_m4stg_frac/a0sum[7] , \i_m4stg_frac/a0sum[6] ,
         \i_m4stg_frac/a0sum[5] , \i_m4stg_frac/a0sum[4] ,
         \i_m4stg_frac/a0sum[3] , \i_m4stg_frac/a0sum[2] ,
         \i_m4stg_frac/a0sum[1] , \i_m4stg_frac/a0sum[0] ,
         \i_m4stg_frac/a0cout[79] , \i_m4stg_frac/a0cout[78] ,
         \i_m4stg_frac/a0cout[77] , \i_m4stg_frac/a0cout[76] ,
         \i_m4stg_frac/a0cout[75] , \i_m4stg_frac/a0cout[74] ,
         \i_m4stg_frac/a0cout[73] , \i_m4stg_frac/a0cout[72] ,
         \i_m4stg_frac/a0cout[71] , \i_m4stg_frac/a0cout[70] ,
         \i_m4stg_frac/a0cout[69] , \i_m4stg_frac/a0cout[68] ,
         \i_m4stg_frac/a0cout[67] , \i_m4stg_frac/a0cout[66] ,
         \i_m4stg_frac/a0cout[65] , \i_m4stg_frac/a0cout[64] ,
         \i_m4stg_frac/a0cout[63] , \i_m4stg_frac/a0cout[62] ,
         \i_m4stg_frac/a0cout[61] , \i_m4stg_frac/a0cout[60] ,
         \i_m4stg_frac/a0cout[59] , \i_m4stg_frac/a0cout[58] ,
         \i_m4stg_frac/a0cout[57] , \i_m4stg_frac/a0cout[56] ,
         \i_m4stg_frac/a0cout[55] , \i_m4stg_frac/a0cout[54] ,
         \i_m4stg_frac/a0cout[53] , \i_m4stg_frac/a0cout[52] ,
         \i_m4stg_frac/a0cout[51] , \i_m4stg_frac/a0cout[50] ,
         \i_m4stg_frac/a0cout[49] , \i_m4stg_frac/a0cout[48] ,
         \i_m4stg_frac/a0cout[47] , \i_m4stg_frac/a0cout[46] ,
         \i_m4stg_frac/a0cout[45] , \i_m4stg_frac/a0cout[44] ,
         \i_m4stg_frac/a0cout[43] , \i_m4stg_frac/a0cout[42] ,
         \i_m4stg_frac/a0cout[41] , \i_m4stg_frac/a0cout[40] ,
         \i_m4stg_frac/a0cout[39] , \i_m4stg_frac/a0cout[38] ,
         \i_m4stg_frac/a0cout[37] , \i_m4stg_frac/a0cout[36] ,
         \i_m4stg_frac/a0cout[35] , \i_m4stg_frac/a0cout[34] ,
         \i_m4stg_frac/a0cout[33] , \i_m4stg_frac/a0cout[32] ,
         \i_m4stg_frac/a0cout[31] , \i_m4stg_frac/a0cout[30] ,
         \i_m4stg_frac/a0cout[29] , \i_m4stg_frac/a0cout[28] ,
         \i_m4stg_frac/a0cout[27] , \i_m4stg_frac/a0cout[26] ,
         \i_m4stg_frac/a0cout[25] , \i_m4stg_frac/a0cout[24] ,
         \i_m4stg_frac/a0cout[23] , \i_m4stg_frac/a0cout[22] ,
         \i_m4stg_frac/a0cout[21] , \i_m4stg_frac/a0cout[20] ,
         \i_m4stg_frac/a0cout[19] , \i_m4stg_frac/a0cout[18] ,
         \i_m4stg_frac/a0cout[17] , \i_m4stg_frac/a0cout[16] ,
         \i_m4stg_frac/a0cout[15] , \i_m4stg_frac/a0cout[14] ,
         \i_m4stg_frac/a0cout[13] , \i_m4stg_frac/a0cout[12] ,
         \i_m4stg_frac/a0cout[11] , \i_m4stg_frac/a0cout[10] ,
         \i_m4stg_frac/a0cout[9] , \i_m4stg_frac/a0cout[8] ,
         \i_m4stg_frac/a0cout[7] , \i_m4stg_frac/a0cout[6] ,
         \i_m4stg_frac/a0cout[5] , \i_m4stg_frac/a0cout[4] ,
         \i_m4stg_frac/b15[2] , \i_m4stg_frac/b12[2] , \i_m4stg_frac/b11[0] ,
         \i_m4stg_frac/b9[2] , \i_m4stg_frac/b8[0] , \i_m4stg_frac/b7[2] ,
         \i_m4stg_frac/b6[0] , \i_m4stg_frac/b4[2] , \i_m4stg_frac/b3[0] ,
         \i_m4stg_frac/b1[2] , \i_m4stg_frac/b0[0] , \i_m4stg_frac/cyc3 ,
         \i_m4stg_frac/cyc1 , n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631;
  wire   [6:0] m3bstg_ld0_inv;
  wire   [12:0] m3stg_exp;
  wire   [12:0] m4stg_exp;
  wire   [12:0] m5stg_exp;
  wire   [52:0] m2stg_frac1_array_in;
  wire   [52:0] m2stg_frac2_array_in;
  wire   [6:0] m3stg_ld0_inv;
  wire   [105:0] m4stg_frac;
  assign so = 1'b0;
  assign mul_exc_out[1] = 1'b0;

  LATCHX1 \fpu_mul_exp_dp/ckbuf_mul_exp_dp/clken_reg  ( .CLK(n709), .D(
        \fpu_mul_exp_dp/ckbuf_mul_exp_dp/N1 ), .Q(
        \fpu_mul_exp_dp/ckbuf_mul_exp_dp/clken ), .QN(n189) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_inc_exp/q_reg[4]  ( .D(m4stg_shl_55), 
        .RSTB(n1360), .SETB(1'b1), .CLK(n1613), .Q(
        \fpu_mul_exp_dp/m5stg_shl_55 ) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_inc_exp/q_reg[0]  ( .D(m4stg_inc_exp_105), 
        .RSTB(n1358), .SETB(1'b1), .CLK(n1613), .Q(
        \fpu_mul_exp_dp/m5stg_inc_exp_105 ) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_inc_exp/q_reg[1]  ( .D(m4stg_inc_exp_55), 
        .RSTB(n1357), .SETB(1'b1), .CLK(n1613), .Q(
        \fpu_mul_exp_dp/m5stg_inc_exp_55 ) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_inc_exp/q_reg[2]  ( .D(m4stg_inc_exp_54), 
        .RSTB(n1358), .SETB(1'b1), .CLK(n1612), .Q(
        \fpu_mul_exp_dp/m5stg_inc_exp_54 ) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[7]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[7] ), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[7] ), .QN(n180) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[8]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[8] ), .SETB(1'b1), .CLK(n1613), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[8] ), .QN(n178) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[9]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[9] ), .SETB(1'b1), .CLK(n1613), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[9] ), .QN(n176) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[10]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[10] ), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[10] ), .QN(n174) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[11]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[11] ), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[11] ), .QN(n172) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[12]  ( .D(n604), .RSTB(n456), 
        .SETB(1'b1), .CLK(n1614), .Q(\fpu_mul_exp_dp/m5stg_exp_pre1[12] ) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[0]  ( .D(n604), .RSTB(n438), 
        .SETB(1'b1), .CLK(n1613), .Q(\fpu_mul_exp_dp/m5stg_exp_pre1[0] ), .QN(
        n168) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[1]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[1] ), .SETB(1'b1), .CLK(n1613), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[1] ), .QN(n166) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[2]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[2] ), .SETB(1'b1), .CLK(n1613), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[2] ), .QN(n164) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[3]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[3] ), .SETB(1'b1), .CLK(n1612), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[3] ), .QN(n162) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[4]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[4] ), .SETB(1'b1), .CLK(n1612), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[4] ), .QN(n160) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[5]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[5] ), .SETB(1'b1), .CLK(n1613), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[5] ), .QN(n158) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre1/q_reg[6]  ( .D(n604), .RSTB(
        \fpu_mul_exp_dp/m4stg_exp_plus1[6] ), .SETB(1'b1), .CLK(n1613), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre1[6] ), .QN(n156) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[12]  ( .D(m5stg_exp[12]), 
        .RSTB(n603), .SETB(n1359), .CLK(n1613), .Q(n877), .QN(n455) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[12]  ( .D(n325), .CLK(n1621), .Q(
        n1288) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[12]  ( .D(n312), .CLK(n1621), .Q(
        n1000), .QN(n148) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[12]  ( .D(n299), .CLK(n1621), .Q(
        \fpu_mul_exp_dp/m3stg_expa[12] ), .QN(n147) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[12]  ( .D(n286), .CLK(n1621), .Q(
        n1119), .QN(n146) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[11]  ( .D(n326), .CLK(n1615), .Q(
        n1349), .QN(n145) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[11]  ( .D(n313), .CLK(n1621), .Q(
        \fpu_mul_exp_dp/m3bstg_exp[11] ), .QN(n144) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[11]  ( .D(n300), .CLK(n1621), .Q(
        \fpu_mul_exp_dp/m3stg_expa[11] ), .QN(n143) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[11]  ( .D(n287), .CLK(n1622), .Q(
        m3stg_exp[11]), .QN(n142) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[10]  ( .D(n327), .CLK(n1616), .Q(
        n1287) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[10]  ( .D(n314), .CLK(n1616), .Q(
        n997), .QN(n140) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[10]  ( .D(n301), .CLK(n1616), .Q(
        n1152), .QN(n448) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[10]  ( .D(n288), .CLK(n1615), .Q(
        m3stg_exp[10]), .QN(n138) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[9]  ( .D(n328), .CLK(n1615), .Q(
        n1348), .QN(n137) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[9]  ( .D(n315), .CLK(n1620), .Q(
        \fpu_mul_exp_dp/m3bstg_exp[9] ), .QN(n136) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[9]  ( .D(n302), .CLK(n1620), .Q(
        \fpu_mul_exp_dp/m3stg_expa[9] ), .QN(n135) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[9]  ( .D(n289), .CLK(n1620), .Q(
        m3stg_exp[9]), .QN(n134) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[8]  ( .D(n329), .CLK(n1620), .Q(
        n1286) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[8]  ( .D(n316), .CLK(n1620), .Q(
        n999), .QN(n132) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[8]  ( .D(n303), .CLK(n1620), .Q(
        \fpu_mul_exp_dp/m3stg_expa[8] ), .QN(n453) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[8]  ( .D(n290), .CLK(n1620), .Q(
        n1203), .QN(n130) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[7]  ( .D(n330), .CLK(n1616), .Q(
        n1285) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[7]  ( .D(n317), .CLK(n1616), .Q(
        n972) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[7]  ( .D(n304), .CLK(n1616), .Q(
        n1153) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[7]  ( .D(n291), .CLK(n1619), .Q(n900) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[6]  ( .D(n331), .CLK(n1619), .Q(
        n1237) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[6]  ( .D(n318), .CLK(n1619), .Q(
        n971) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[6]  ( .D(n305), .CLK(n1619), .Q(
        n1122) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[6]  ( .D(n292), .CLK(n1619), .Q(
        n1114), .QN(n122) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[5]  ( .D(n332), .CLK(n1616), .Q(
        n1236) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[5]  ( .D(n319), .CLK(n1620), .Q(
        n996), .QN(n120) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[5]  ( .D(n306), .CLK(n1620), .Q(
        n1213), .QN(n119) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[5]  ( .D(n293), .CLK(n1620), .Q(
        m3stg_exp[5]), .QN(n118) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[4]  ( .D(n333), .CLK(n1620), .Q(
        n1235) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[4]  ( .D(n320), .CLK(n1620), .Q(
        n970) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[4]  ( .D(n307), .CLK(n1620), .Q(
        n1211), .QN(n115) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[4]  ( .D(n294), .CLK(n1620), .Q(n888), .QN(n114) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[3]  ( .D(n334), .CLK(n1615), .Q(
        n1239) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[3]  ( .D(n321), .CLK(n1615), .Q(
        n1001), .QN(n112) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[3]  ( .D(n308), .CLK(n1615), .Q(
        n1214), .QN(n111) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[3]  ( .D(n295), .CLK(n1619), .Q(
        m3stg_exp[3]), .QN(n110) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[2]  ( .D(n335), .CLK(n1619), .Q(
        n1234) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[2]  ( .D(n322), .CLK(n1619), .Q(
        n969) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[2]  ( .D(n309), .CLK(n1619), .Q(
        n1212), .QN(n107) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[2]  ( .D(n296), .CLK(n1619), .Q(
        n1166), .QN(n106) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[1]  ( .D(n336), .CLK(n1617), .Q(
        n1233) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[1]  ( .D(n323), .CLK(n1619), .Q(
        n998), .QN(n104) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[1]  ( .D(n310), .CLK(n1619), .Q(
        \fpu_mul_exp_dp/m3stg_expa[1] ), .QN(n103) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[1]  ( .D(n297), .CLK(n1619), .Q(
        n1115), .QN(n452) );
  DFFX1 \fpu_mul_exp_dp/i_m3astg_exp/q_reg[0]  ( .D(n337), .CLK(n1615), .Q(
        n1238) );
  DFFX1 \fpu_mul_exp_dp/i_m3bstg_exp/q_reg[0]  ( .D(n324), .CLK(n1617), .Q(
        n968) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_expa/q_reg[0]  ( .D(n311), .CLK(n1619), .Q(
        n1154) );
  DFFX1 \fpu_mul_exp_dp/i_m3stg_exp/q_reg[0]  ( .D(n298), .CLK(n1618), .Q(n895), .QN(n98) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[9]  ( .D(n341), .CLK(n1616), .Q(
        n1210), .QN(n441) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[7]  ( .D(n342), .CLK(n1616), .Q(
        n1140), .QN(n454) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[8]  ( .D(n1608), .RSTB(
        m2stg_exp_017f), .SETB(n94), .CLK(n1615), .Q(
        \fpu_mul_exp_dp/m2stg_exp[8] ), .QN(n449) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[6]  ( .D(n343), .CLK(n1616), .Q(n993) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[5]  ( .D(n344), .CLK(n1617), .Q(n992) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[4]  ( .D(n345), .CLK(n1616), .Q(n991) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[3]  ( .D(n346), .CLK(n1615), .Q(n995) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[2]  ( .D(n347), .CLK(n1617), .Q(n990) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[1]  ( .D(n348), .CLK(n1617), .Q(n989) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[0]  ( .D(n349), .CLK(n1615), .Q(n994) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[0]  ( .D(n350), .CLK(n1617), .Q(
        n1226) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[1]  ( .D(n351), .CLK(n1618), .Q(
        n1225) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[2]  ( .D(n352), .CLK(n1618), .Q(
        n1232) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[3]  ( .D(n353), .CLK(n1618), .Q(
        n963) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[4]  ( .D(n354), .CLK(n1618), .Q(
        n904) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[5]  ( .D(n355), .CLK(n1617), .Q(
        n962) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[6]  ( .D(n356), .CLK(n1617), .Q(
        n903) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[7]  ( .D(n357), .CLK(n1617), .Q(
        n965) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[8]  ( .D(n358), .CLK(n1618), .Q(
        n1177) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[9]  ( .D(n359), .CLK(n1616), .Q(
        n1175) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in1/q_reg[10]  ( .D(n360), .CLK(n1617), 
        .Q(n1178) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[0]  ( .D(n361), .CLK(n1617), .Q(
        n1227) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[1]  ( .D(n362), .CLK(n1618), .Q(
        n1228) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[2]  ( .D(n363), .CLK(n1618), .Q(
        n1231) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[3]  ( .D(n364), .CLK(n1618), .Q(
        n964) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[4]  ( .D(n365), .CLK(n1617), .Q(
        n905) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[5]  ( .D(n366), .CLK(n1618), .Q(
        n961) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[6]  ( .D(n367), .CLK(n1617), .Q(
        n902) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[7]  ( .D(n368), .CLK(n1618), .Q(
        n975) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[8]  ( .D(n369), .CLK(n1618), .Q(
        n1176) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[9]  ( .D(n370), .CLK(n1618), .Q(
        n1179) );
  DFFX1 \fpu_mul_exp_dp/i_m1stg_exp_in2/q_reg[10]  ( .D(n371), .CLK(n1618), 
        .Q(n1194) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[11]  ( .D(n274), .CLK(n1621), .Q(
        m4stg_exp[11]), .QN(n443) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[11]  ( .D(n1608), .RSTB(
        m4stg_exp[11]), .SETB(1'b1), .CLK(n1615), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[11] ), .QN(n63) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[11]  ( .D(m5stg_exp[11]), 
        .RSTB(n603), .SETB(n1357), .CLK(n1612), .Q(n212), .QN(n61) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[10]  ( .D(n275), .CLK(n1621), .Q(
        m4stg_exp[10]), .QN(n60) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[10]  ( .D(n1608), .RSTB(
        m4stg_exp[10]), .SETB(1'b1), .CLK(n1615), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[10] ), .QN(n59) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[10]  ( .D(n603), .RSTB(
        m5stg_exp[10]), .SETB(n1359), .CLK(n1612), .Q(n211), .QN(n57) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[9]  ( .D(n276), .CLK(n1621), .Q(
        m4stg_exp[9]), .QN(n445) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[9]  ( .D(n1608), .RSTB(
        m4stg_exp[9]), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[9] ), .QN(n55) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[9]  ( .D(n603), .RSTB(
        m5stg_exp[9]), .SETB(n1358), .CLK(n1612), .Q(n210), .QN(n53) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[8]  ( .D(n277), .CLK(n1621), .Q(
        m4stg_exp[8]), .QN(n52) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[8]  ( .D(n1608), .RSTB(
        m4stg_exp[8]), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[8] ), .QN(n51) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[8]  ( .D(n603), .RSTB(
        m5stg_exp[8]), .SETB(n1360), .CLK(n1612), .Q(n209), .QN(n49) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[7]  ( .D(n278), .CLK(n1621), .Q(
        m4stg_exp[7]), .QN(n447) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[7]  ( .D(n604), .RSTB(
        m4stg_exp[7]), .SETB(1'b1), .CLK(n1611), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[7] ), .QN(n47) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[7]  ( .D(m5stg_exp[7]), 
        .RSTB(n603), .SETB(n1358), .CLK(n1612), .Q(n208), .QN(n45) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[6]  ( .D(n279), .CLK(n1621), .Q(
        m4stg_exp[6]), .QN(n44) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[6]  ( .D(n604), .RSTB(
        m4stg_exp[6]), .SETB(1'b1), .CLK(n1611), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[6] ), .QN(n43) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[5]  ( .D(n280), .CLK(n1621), .Q(
        m4stg_exp[5]), .QN(n444) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[5]  ( .D(n1608), .RSTB(
        m4stg_exp[5]), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[5] ), .QN(n40) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[5]  ( .D(n603), .RSTB(
        m5stg_exp[5]), .SETB(n1358), .CLK(n1611), .Q(n206), .QN(n38) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[4]  ( .D(n281), .CLK(n1621), .Q(
        m4stg_exp[4]), .QN(n37) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[4]  ( .D(n1608), .RSTB(
        m4stg_exp[4]), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[4] ), .QN(n36) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[4]  ( .D(n603), .RSTB(
        m5stg_exp[4]), .SETB(n1360), .CLK(n1611), .Q(n205), .QN(n34) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[3]  ( .D(n282), .CLK(n1622), .Q(
        m4stg_exp[3]), .QN(n446) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[3]  ( .D(n604), .RSTB(
        m4stg_exp[3]), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[3] ), .QN(n32) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[3]  ( .D(n603), .RSTB(
        m5stg_exp[3]), .SETB(n1357), .CLK(n1612), .Q(n204), .QN(n30) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[2]  ( .D(n283), .CLK(n1622), .Q(
        m4stg_exp[2]), .QN(n29) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[2]  ( .D(n604), .RSTB(
        m4stg_exp[2]), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[2] ), .QN(n28) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[2]  ( .D(n603), .RSTB(
        m5stg_exp[2]), .SETB(n1360), .CLK(n1612), .Q(n203), .QN(n26) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[1]  ( .D(n284), .CLK(n1622), .Q(
        m4stg_exp[1]), .QN(n442) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[1]  ( .D(n604), .RSTB(
        m4stg_exp[1]), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[1] ), .QN(n24) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[1]  ( .D(n603), .RSTB(
        m5stg_exp[1]), .SETB(n1357), .CLK(n1612), .Q(n202), .QN(n22) );
  DFFX1 \fpu_mul_exp_dp/i_m4stg_exp/q_reg[0]  ( .D(n285), .CLK(n1622), .Q(
        m4stg_exp[0]), .QN(n438) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre2/q_reg[0]  ( .D(n604), .RSTB(
        m4stg_exp[0]), .SETB(1'b1), .CLK(n1614), .Q(
        \fpu_mul_exp_dp/m5stg_exp_pre2[0] ), .QN(n20) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[0]  ( .D(n603), .RSTB(
        m5stg_exp[0]), .SETB(n1359), .CLK(n1612), .Q(n201), .QN(n18) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[12]  ( .D(n338), .CLK(n1617), .Q(
        \fpu_mul_exp_dp/m2stg_exp[12] ), .QN(n17) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[11]  ( .D(n339), .CLK(n1616), .Q(
        n878), .QN(n1277) );
  DFFX1 \fpu_mul_exp_dp/i_m2stg_exp/q_reg[10]  ( .D(n340), .CLK(n1616), .Q(
        n876), .QN(n439) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_inc_exp/q_reg[3]  ( .D(m4stg_shl_54), 
        .RSTB(n1359), .SETB(1'b1), .CLK(n1613), .Q(
        \fpu_mul_exp_dp/m5stg_shl_54 ) );
  DFFSSRX1 \fpu_mul_exp_dp/i_m5stg_exp_pre3/q_reg[6]  ( .D(n603), .RSTB(
        m5stg_exp[6]), .SETB(n1360), .CLK(n1611), .Q(n207), .QN(n12) );
  DFFX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[0]  ( .D(n272), .CLK(n1615), .Q(
        mul_exp_out[0]) );
  DFFSSRX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[1]  ( .D(m5stg_exp[1]), .RSTB(
        n594), .SETB(n196), .CLK(n1611), .Q(mul_exp_out[1]), .QN(n10) );
  DFFSSRX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[2]  ( .D(m5stg_exp[2]), .RSTB(
        n594), .SETB(n195), .CLK(n1611), .Q(mul_exp_out[2]), .QN(n9) );
  DFFSSRX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[3]  ( .D(m5stg_exp[3]), .RSTB(
        n594), .SETB(n194), .CLK(n1611), .Q(mul_exp_out[3]), .QN(n8) );
  DFFSSRX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[4]  ( .D(m5stg_exp[4]), .RSTB(
        n594), .SETB(n193), .CLK(n1611), .Q(mul_exp_out[4]), .QN(n7) );
  DFFSSRX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[5]  ( .D(m5stg_exp[5]), .RSTB(
        n594), .SETB(n192), .CLK(n1611), .Q(mul_exp_out[5]), .QN(n6) );
  DFFSSRX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[6]  ( .D(m5stg_exp[6]), .RSTB(
        n594), .SETB(n191), .CLK(n1611), .Q(mul_exp_out[6]), .QN(n5) );
  DFFSSRX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[7]  ( .D(m5stg_exp[7]), .RSTB(
        n594), .SETB(n190), .CLK(n1611), .Q(mul_exp_out[7]), .QN(n4) );
  DFFX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[8]  ( .D(n271), .CLK(n1622), .Q(
        mul_exp_out[8]) );
  DFFX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[9]  ( .D(n270), .CLK(n1622), .Q(
        mul_exp_out[9]) );
  DFFX1 \fpu_mul_exp_dp/i_mul_exp_out/q_reg[10]  ( .D(n269), .CLK(n1622), .Q(
        mul_exp_out[10]) );
  DFFX1 \fpu_mul_ctl/i_m4stg_right_shift/q_reg[0]  ( .D(\fpu_mul_ctl/n384 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/m4stg_right_shift ), .QN(m4stg_inc_exp_55)
         );
  DFFX1 \fpu_mul_ctl/i_m4stg_expadd_eq_0/q_reg[0]  ( .D(\fpu_mul_ctl/n385 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/m4stg_expadd_eq_0 ), .QN(\fpu_mul_ctl/n1 )
         );
  DFFX1 \fpu_mul_ctl/i_m3bstg_ld0_inv/q_reg[6]  ( .D(\fpu_mul_ctl/n386 ), 
        .CLK(rclk), .Q(m3bstg_ld0_inv[6]) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_ld0_inv/q_reg[5]  ( .D(\fpu_mul_ctl/n387 ), 
        .CLK(rclk), .Q(m3bstg_ld0_inv[5]) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_ld0_inv/q_reg[4]  ( .D(\fpu_mul_ctl/n388 ), 
        .CLK(rclk), .Q(m3bstg_ld0_inv[4]) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_ld0_inv/q_reg[3]  ( .D(\fpu_mul_ctl/n389 ), 
        .CLK(rclk), .Q(m3bstg_ld0_inv[3]) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_ld0_inv/q_reg[2]  ( .D(\fpu_mul_ctl/n390 ), 
        .CLK(rclk), .Q(m3bstg_ld0_inv[2]) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_ld0_inv/q_reg[1]  ( .D(\fpu_mul_ctl/n391 ), 
        .CLK(rclk), .Q(m3bstg_ld0_inv[1]) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_ld0_inv/q_reg[0]  ( .D(\fpu_mul_ctl/n392 ), 
        .CLK(rclk), .Q(m3bstg_ld0_inv[0]) );
  DFFX1 \fpu_mul_ctl/i_m3astg_ld0_inv/q_reg[6]  ( .D(\fpu_mul_ctl/n393 ), 
        .CLK(rclk), .Q(n1296) );
  DFFX1 \fpu_mul_ctl/i_m3astg_ld0_inv/q_reg[5]  ( .D(\fpu_mul_ctl/n394 ), 
        .CLK(rclk), .Q(n1295) );
  DFFX1 \fpu_mul_ctl/i_m3astg_ld0_inv/q_reg[4]  ( .D(\fpu_mul_ctl/n395 ), 
        .CLK(rclk), .Q(n1294) );
  DFFX1 \fpu_mul_ctl/i_m3astg_ld0_inv/q_reg[3]  ( .D(\fpu_mul_ctl/n396 ), 
        .CLK(rclk), .Q(n1293) );
  DFFX1 \fpu_mul_ctl/i_m3astg_ld0_inv/q_reg[2]  ( .D(\fpu_mul_ctl/n397 ), 
        .CLK(rclk), .Q(n1292) );
  DFFX1 \fpu_mul_ctl/i_m3astg_ld0_inv/q_reg[1]  ( .D(\fpu_mul_ctl/n398 ), 
        .CLK(rclk), .Q(n1291) );
  DFFX1 \fpu_mul_ctl/i_m3astg_ld0_inv/q_reg[0]  ( .D(\fpu_mul_ctl/n399 ), 
        .CLK(rclk), .Q(n1290) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_2/q_reg[5]  ( .D(\fpu_mul_ctl/n400 ), .CLK(
        rclk), .Q(n1162), .QN(\fpu_mul_ctl/n16 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_2/q_reg[4]  ( .D(\fpu_mul_ctl/n401 ), .CLK(
        rclk), .Q(n1322), .QN(\fpu_mul_ctl/n17 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_2/q_reg[3]  ( .D(\fpu_mul_ctl/n402 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/m2stg_ld0_2[3] ), .QN(\fpu_mul_ctl/n18 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_2/q_reg[2]  ( .D(\fpu_mul_ctl/n403 ), .CLK(
        rclk), .Q(n1321), .QN(\fpu_mul_ctl/n19 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_2/q_reg[1]  ( .D(\fpu_mul_ctl/n404 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/m2stg_ld0_2[1] ), .QN(\fpu_mul_ctl/n20 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_2/q_reg[0]  ( .D(\fpu_mul_ctl/n405 ), .CLK(
        rclk), .Q(n1181) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_1/q_reg[5]  ( .D(\fpu_mul_ctl/n406 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/m2stg_ld0_1[5] ), .QN(\fpu_mul_ctl/n22 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_1/q_reg[4]  ( .D(\fpu_mul_ctl/n407 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/m2stg_ld0_1[4] ), .QN(\fpu_mul_ctl/n23 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_1/q_reg[3]  ( .D(\fpu_mul_ctl/n408 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/m2stg_ld0_1[3] ), .QN(\fpu_mul_ctl/n24 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_1/q_reg[2]  ( .D(\fpu_mul_ctl/n409 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/m2stg_ld0_1[2] ), .QN(\fpu_mul_ctl/n25 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_1/q_reg[1]  ( .D(\fpu_mul_ctl/n410 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/m2stg_ld0_1[1] ), .QN(\fpu_mul_ctl/n26 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_ld0_1/q_reg[0]  ( .D(\fpu_mul_ctl/n411 ), .CLK(
        rclk), .Q(n974) );
  DFFX1 \fpu_mul_ctl/i_mul_nx_out/q_reg[0]  ( .D(\fpu_mul_ctl/n412 ), .CLK(
        rclk), .Q(n1345), .QN(\fpu_mul_ctl/n28 ) );
  DFFX1 \fpu_mul_ctl/i_mul_uf_out/q_reg[0]  ( .D(\fpu_mul_ctl/n413 ), .CLK(
        rclk), .Q(mul_exc_out[2]) );
  DFFX1 \fpu_mul_ctl/i_mul_of_out_cout/q_reg[0]  ( .D(\fpu_mul_ctl/n414 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/mul_of_out_cout ), .QN(\fpu_mul_ctl/n30 )
         );
  DFFX1 \fpu_mul_ctl/i_mul_of_out_tmp2/q_reg[0]  ( .D(\fpu_mul_ctl/n415 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/mul_of_out_tmp2 ), .QN(\fpu_mul_ctl/n31 )
         );
  DFFX1 \fpu_mul_ctl/i_mul_of_out_tmp1/q_reg[0]  ( .D(\fpu_mul_ctl/n416 ), 
        .CLK(rclk), .Q(n1346), .QN(\fpu_mul_ctl/n32 ) );
  DFFX1 \fpu_mul_ctl/i_mul_nv_out/q_reg[0]  ( .D(\fpu_mul_ctl/n417 ), .CLK(
        rclk), .Q(mul_exc_out[4]) );
  DFFX1 \fpu_mul_ctl/i_mul_sign_out/q_reg[0]  ( .D(\fpu_mul_ctl/n418 ), .CLK(
        rclk), .Q(mul_sign_out) );
  DFFX1 \fpu_mul_ctl/i_m5stg_of_mask/q_reg[0]  ( .D(\fpu_mul_ctl/n419 ), .CLK(
        rclk), .Q(n981), .QN(\fpu_mul_ctl/n271 ) );
  DFFX1 \fpu_mul_ctl/i_m5stg_nv/q_reg[0]  ( .D(\fpu_mul_ctl/n420 ), .CLK(rclk), 
        .Q(n1276) );
  DFFX1 \fpu_mul_ctl/i_m5stg_sign/q_reg[0]  ( .D(\fpu_mul_ctl/n421 ), .CLK(
        rclk), .Q(n988), .QN(\fpu_mul_ctl/n733 ) );
  DFFX1 \fpu_mul_ctl/i_m4stg_of_mask/q_reg[0]  ( .D(\fpu_mul_ctl/n422 ), .CLK(
        rclk), .Q(n1275) );
  DFFX1 \fpu_mul_ctl/i_m4stg_nv/q_reg[0]  ( .D(\fpu_mul_ctl/n423 ), .CLK(rclk), 
        .Q(n1028) );
  DFFX1 \fpu_mul_ctl/i_m4stg_sign/q_reg[0]  ( .D(\fpu_mul_ctl/n424 ), .CLK(
        rclk), .Q(n1274) );
  DFFX1 \fpu_mul_ctl/i_m3stg_of_mask/q_reg[0]  ( .D(\fpu_mul_ctl/n425 ), .CLK(
        rclk), .Q(n1027) );
  DFFX1 \fpu_mul_ctl/i_m3stg_nv/q_reg[0]  ( .D(\fpu_mul_ctl/n426 ), .CLK(rclk), 
        .Q(n1273) );
  DFFX1 \fpu_mul_ctl/i_m3stg_sign/q_reg[0]  ( .D(\fpu_mul_ctl/n427 ), .CLK(
        rclk), .Q(n1026) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_of_mask/q_reg[0]  ( .D(\fpu_mul_ctl/n428 ), 
        .CLK(rclk), .Q(n1272) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_nv/q_reg[0]  ( .D(\fpu_mul_ctl/n429 ), .CLK(rclk), .Q(n1025) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_sign/q_reg[0]  ( .D(\fpu_mul_ctl/n430 ), .CLK(
        rclk), .Q(n1271) );
  DFFX1 \fpu_mul_ctl/i_m3astg_of_mask/q_reg[0]  ( .D(\fpu_mul_ctl/n431 ), 
        .CLK(rclk), .Q(n1024) );
  DFFX1 \fpu_mul_ctl/i_m3astg_nv/q_reg[0]  ( .D(\fpu_mul_ctl/n432 ), .CLK(rclk), .Q(n1289) );
  DFFX1 \fpu_mul_ctl/i_m3astg_sign/q_reg[0]  ( .D(\fpu_mul_ctl/n433 ), .CLK(
        rclk), .Q(n1023) );
  DFFX1 \fpu_mul_ctl/i_m2stg_of_mask/q_reg[0]  ( .D(\fpu_mul_ctl/n434 ), .CLK(
        rclk), .Q(n1281) );
  DFFX1 \fpu_mul_ctl/i_m2stg_sign2/q_reg[0]  ( .D(\fpu_mul_ctl/n435 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/m2stg_sign2 ), .QN(\fpu_mul_ctl/n50 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_sign1/q_reg[0]  ( .D(\fpu_mul_ctl/n436 ), .CLK(
        rclk), .Q(n980), .QN(\fpu_mul_ctl/n51 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_sign2/q_reg[0]  ( .D(\fpu_mul_ctl/n437 ), .CLK(
        rclk), .Q(n1335), .QN(\fpu_mul_ctl/n52 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_sign1/q_reg[0]  ( .D(\fpu_mul_ctl/n438 ), .CLK(
        rclk), .Q(n1270) );
  DFFSSRX1 \fpu_mul_ctl/i_mul_pipe_active/q_reg[0]  ( .D(\fpu_mul_ctl/n379 ), 
        .RSTB(\fpu_mul_ctl/n380 ), .SETB(\fpu_mul_ctl/n735 ), .CLK(rclk), .QN(
        mul_pipe_active) );
  DFFX1 \fpu_mul_ctl/i_m6stg_id/q_reg[9]  ( .D(\fpu_mul_ctl/n448 ), .CLK(rclk), 
        .Q(n1262) );
  DFFX1 \fpu_mul_ctl/i_m6stg_id/q_reg[8]  ( .D(\fpu_mul_ctl/n439 ), .CLK(rclk), 
        .Q(n1269) );
  DFFX1 \fpu_mul_ctl/i_m6stg_id/q_reg[7]  ( .D(\fpu_mul_ctl/n440 ), .CLK(rclk), 
        .Q(n1268) );
  DFFX1 \fpu_mul_ctl/i_m6stg_id/q_reg[6]  ( .D(\fpu_mul_ctl/n441 ), .CLK(rclk), 
        .Q(n1267) );
  DFFX1 \fpu_mul_ctl/i_m6stg_id/q_reg[5]  ( .D(\fpu_mul_ctl/n442 ), .CLK(rclk), 
        .Q(n1266) );
  DFFX1 \fpu_mul_ctl/i_m6stg_id/q_reg[4]  ( .D(\fpu_mul_ctl/n443 ), .CLK(rclk), 
        .Q(n1265) );
  DFFX1 \fpu_mul_ctl/i_m6stg_id/q_reg[3]  ( .D(\fpu_mul_ctl/n444 ), .CLK(rclk), 
        .Q(n1264) );
  DFFX1 \fpu_mul_ctl/i_m6stg_id/q_reg[2]  ( .D(\fpu_mul_ctl/n445 ), .CLK(rclk), 
        .Q(n1263) );
  DFFX1 \fpu_mul_ctl/i_m6stg_id/q_reg[1]  ( .D(\fpu_mul_ctl/n446 ), .CLK(rclk), 
        .Q(n1217) );
  DFFX1 \fpu_mul_ctl/i_m6stg_id/q_reg[0]  ( .D(\fpu_mul_ctl/n447 ), .CLK(rclk), 
        .Q(n1216) );
  DFFX1 \fpu_mul_ctl/i_m1stg_mul/q_reg[0]  ( .D(\fpu_mul_ctl/i_m1stg_mul/N3 ), 
        .CLK(rclk), .Q(n1215) );
  DFFX1 \fpu_mul_ctl/i_m5stg_opdec/q_reg[0]  ( .D(\fpu_mul_ctl/n454 ), .CLK(
        rclk), .Q(m5stg_fmuld) );
  DFFX1 \fpu_mul_ctl/i_m5stg_fmulda/q_reg[0]  ( .D(\fpu_mul_ctl/n458 ), .CLK(
        rclk), .Q(m5stg_fmulda) );
  DFFX1 \fpu_mul_ctl/i_m4stg_opdec/q_reg[0]  ( .D(\fpu_mul_ctl/n459 ), .CLK(
        rclk), .Q(n966) );
  DFFX1 \fpu_mul_ctl/i_m3stg_opdec/q_reg[0]  ( .D(\fpu_mul_ctl/n463 ), .CLK(
        rclk), .Q(n1258) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_opdec/q_reg[0]  ( .D(\fpu_mul_ctl/n467 ), .CLK(
        rclk), .Q(n1019) );
  DFFX1 \fpu_mul_ctl/i_m3astg_opdec/q_reg[0]  ( .D(\fpu_mul_ctl/n471 ), .CLK(
        rclk), .Q(n1255) );
  DFFX1 \fpu_mul_ctl/i_m2stg_opdec/q_reg[1]  ( .D(\fpu_mul_ctl/n475 ), .CLK(
        rclk), .Q(m2stg_fmuld) );
  DFFX1 \fpu_mul_ctl/i_m5stg_opdec/q_reg[3]  ( .D(\fpu_mul_ctl/n451 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/m5stg_opdec[4] ) );
  DFFX1 \fpu_mul_ctl/i_m4stg_opdec/q_reg[3]  ( .D(\fpu_mul_ctl/n455 ), .CLK(
        rclk), .Q(n1138) );
  DFFX1 \fpu_mul_ctl/i_m3stg_opdec/q_reg[3]  ( .D(\fpu_mul_ctl/n460 ), .CLK(
        rclk), .Q(n883) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_opdec/q_reg[3]  ( .D(\fpu_mul_ctl/n464 ), .CLK(
        rclk), .Q(n901) );
  DFFX1 \fpu_mul_ctl/i_m3astg_opdec/q_reg[3]  ( .D(\fpu_mul_ctl/n468 ), .CLK(
        rclk), .Q(n1139) );
  DFFX1 \fpu_mul_ctl/i_m2stg_opdec/q_reg[4]  ( .D(\fpu_mul_ctl/n472 ), .CLK(
        rclk), .Q(n954) );
  DFFX1 \fpu_mul_ctl/i_m6stg_opdec/q_reg[1]  ( .D(\fpu_mul_ctl/n449 ), .CLK(
        rclk), .Q(m6stg_fmul_dbl_dst) );
  DFFX1 \fpu_mul_ctl/i_m5stg_opdec/q_reg[2]  ( .D(\fpu_mul_ctl/n452 ), .CLK(
        rclk), .Q(n1261) );
  DFFX1 \fpu_mul_ctl/i_m4stg_opdec/q_reg[2]  ( .D(\fpu_mul_ctl/n456 ), .CLK(
        rclk), .Q(n1022) );
  DFFX1 \fpu_mul_ctl/i_m3stg_opdec/q_reg[2]  ( .D(\fpu_mul_ctl/n461 ), .CLK(
        rclk), .Q(n1259) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_opdec/q_reg[2]  ( .D(\fpu_mul_ctl/n465 ), .CLK(
        rclk), .Q(n1020) );
  DFFX1 \fpu_mul_ctl/i_m3astg_opdec/q_reg[2]  ( .D(\fpu_mul_ctl/n469 ), .CLK(
        rclk), .Q(n1256) );
  DFFX1 \fpu_mul_ctl/i_m2stg_opdec/q_reg[3]  ( .D(\fpu_mul_ctl/n473 ), .CLK(
        rclk), .Q(n1017) );
  DFFX1 \fpu_mul_ctl/i_m2stg_opdec/q_reg[0]  ( .D(\fpu_mul_ctl/n476 ), .CLK(
        rclk), .Q(m2stg_fsmuld) );
  DFFX1 \fpu_mul_ctl/i_m6stg_opdec/q_reg[0]  ( .D(\fpu_mul_ctl/n450 ), .CLK(
        rclk), .Q(m6stg_fmuls) );
  DFFX1 \fpu_mul_ctl/i_m5stg_opdec/q_reg[1]  ( .D(\fpu_mul_ctl/n453 ), .CLK(
        rclk), .Q(m5stg_fmuls), .QN(n1219) );
  DFFX1 \fpu_mul_ctl/i_m4stg_opdec/q_reg[1]  ( .D(\fpu_mul_ctl/n457 ), .CLK(
        rclk), .Q(n1260) );
  DFFX1 \fpu_mul_ctl/i_m3stg_opdec/q_reg[1]  ( .D(\fpu_mul_ctl/n462 ), .CLK(
        rclk), .Q(n1021) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_opdec/q_reg[1]  ( .D(\fpu_mul_ctl/n466 ), .CLK(
        rclk), .Q(n1257) );
  DFFX1 \fpu_mul_ctl/i_m3astg_opdec/q_reg[1]  ( .D(\fpu_mul_ctl/n470 ), .CLK(
        rclk), .Q(n1018) );
  DFFX1 \fpu_mul_ctl/i_m2stg_opdec/q_reg[2]  ( .D(\fpu_mul_ctl/n474 ), .CLK(
        rclk), .Q(m2stg_fmuls), .QN(n1218) );
  DFFX1 \fpu_mul_ctl/i_m1stg_op/q_reg[7]  ( .D(\fpu_mul_ctl/i_m1stg_op/N10 ), 
        .CLK(rclk), .Q(n1350), .QN(\fpu_mul_ctl/n93 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_op/q_reg[0]  ( .D(\fpu_mul_ctl/i_m1stg_op/N3 ), 
        .CLK(rclk), .Q(n1206), .QN(\fpu_mul_ctl/n270 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_op/q_reg[1]  ( .D(\fpu_mul_ctl/i_m1stg_op/N4 ), 
        .CLK(rclk), .Q(n1282), .QN(\fpu_mul_ctl/n269 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_op/q_reg[2]  ( .D(\fpu_mul_ctl/i_m1stg_op/N5 ), 
        .CLK(rclk), .Q(n1351), .QN(\fpu_mul_ctl/n94 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_op/q_reg[3]  ( .D(\fpu_mul_ctl/i_m1stg_op/N6 ), 
        .CLK(rclk), .Q(n1342), .QN(\fpu_mul_ctl/n95 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_op/q_reg[4]  ( .D(\fpu_mul_ctl/i_m1stg_op/N7 ), 
        .CLK(rclk), .Q(n1347), .QN(\fpu_mul_ctl/n96 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_op/q_reg[5]  ( .D(\fpu_mul_ctl/i_m1stg_op/N8 ), 
        .CLK(rclk), .Q(n1055), .QN(\fpu_mul_ctl/n257 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_op/q_reg[6]  ( .D(\fpu_mul_ctl/i_m1stg_op/N9 ), 
        .CLK(rclk), .Q(n1343), .QN(\fpu_mul_ctl/n97 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_snan_in1/q_reg[0]  ( .D(\fpu_mul_ctl/n531 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/n730 ), .QN(n1332) );
  DFFX1 \fpu_mul_ctl/i_m2stg_qnan_in1/q_reg[0]  ( .D(\fpu_mul_ctl/n529 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/n731 ), .QN(\fpu_mul_ctl/n266 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_inf_in/q_reg[0]  ( .D(\fpu_mul_ctl/n534 ), .CLK(
        rclk), .Q(n1341), .QN(\fpu_mul_ctl/n98 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_inf_in1/q_reg[0]  ( .D(\fpu_mul_ctl/n535 ), .CLK(
        rclk), .Q(n1029) );
  DFFX1 \fpu_mul_ctl/i_mul_frac_in1_51/q_reg[0]  ( .D(\fpu_mul_ctl/n561 ), 
        .CLK(rclk), .Q(n893), .QN(\fpu_mul_ctl/n272 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_zero_in/q_reg[0]  ( .D(\fpu_mul_ctl/n545 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/m2stg_zero_in ), .QN(\fpu_mul_ctl/n100 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_zero_in1/q_reg[0]  ( .D(\fpu_mul_ctl/n547 ), 
        .CLK(rclk), .Q(n1030) );
  DFFX1 \fpu_mul_ctl/i_mul_frac_in1_54/q_reg[0]  ( .D(\fpu_mul_ctl/n560 ), 
        .CLK(rclk), .Q(n894), .QN(\fpu_mul_ctl/n273 ) );
  DFFX1 \fpu_mul_ctl/i_mul_frac_in1_53_0_neq_0/q_reg[0]  ( .D(
        \fpu_mul_ctl/n559 ), .CLK(rclk), .Q(n1336), .QN(\fpu_mul_ctl/n102 ) );
  DFFX1 \fpu_mul_ctl/i_mul_frac_in1_50_0_neq_0/q_reg[0]  ( .D(
        \fpu_mul_ctl/n558 ), .CLK(rclk), .Q(n1204), .QN(\fpu_mul_ctl/n103 ) );
  DFFX1 \fpu_mul_ctl/i_mul_frac_in1_53_32_neq_0/q_reg[0]  ( .D(
        \fpu_mul_ctl/n557 ), .CLK(rclk), .Q(n1205), .QN(\fpu_mul_ctl/n104 ) );
  DFFX1 \fpu_mul_ctl/i_mul_exp_in1_exp_eq_0/q_reg[0]  ( .D(\fpu_mul_ctl/n556 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/n263 ), .QN(n1163) );
  DFFX1 \fpu_mul_ctl/i_mul_exp_in1_exp_neq_ffs/q_reg[0]  ( .D(
        \fpu_mul_ctl/n555 ), .CLK(rclk), .Q(n1037), .QN(\fpu_mul_ctl/n256 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_snan_in2/q_reg[0]  ( .D(\fpu_mul_ctl/n530 ), 
        .CLK(rclk), .Q(n1164), .QN(\fpu_mul_ctl/n262 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_qnan_in2/q_reg[0]  ( .D(\fpu_mul_ctl/n528 ), 
        .CLK(rclk), .Q(n1328), .QN(\fpu_mul_ctl/n106 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_nan_in2/q_reg[0]  ( .D(\fpu_mul_ctl/n536 ), .CLK(
        rclk), .Q(n1344), .QN(\fpu_mul_ctl/n107 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_inf_in2/q_reg[0]  ( .D(\fpu_mul_ctl/n533 ), .CLK(
        rclk), .Q(n1297) );
  DFFX1 \fpu_mul_ctl/i_mul_frac_in2_51/q_reg[0]  ( .D(\fpu_mul_ctl/n554 ), 
        .CLK(rclk), .Q(n1170), .QN(\fpu_mul_ctl/n267 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_zero_in2/q_reg[0]  ( .D(\fpu_mul_ctl/n546 ), 
        .CLK(rclk), .Q(n1284) );
  DFFX1 \fpu_mul_ctl/i_mul_frac_in2_54/q_reg[0]  ( .D(\fpu_mul_ctl/n553 ), 
        .CLK(rclk), .Q(n1167), .QN(\fpu_mul_ctl/n268 ) );
  DFFX1 \fpu_mul_ctl/i_mul_frac_in2_53_0_neq_0/q_reg[0]  ( .D(
        \fpu_mul_ctl/n552 ), .CLK(rclk), .Q(n1337), .QN(\fpu_mul_ctl/n110 ) );
  DFFX1 \fpu_mul_ctl/i_mul_frac_in2_50_0_neq_0/q_reg[0]  ( .D(
        \fpu_mul_ctl/n551 ), .CLK(rclk), .Q(n1198), .QN(\fpu_mul_ctl/n111 ) );
  DFFX1 \fpu_mul_ctl/i_mul_frac_in2_53_32_neq_0/q_reg[0]  ( .D(
        \fpu_mul_ctl/n550 ), .CLK(rclk), .Q(n1197), .QN(\fpu_mul_ctl/n112 ) );
  DFFX1 \fpu_mul_ctl/i_mul_exp_in2_exp_eq_0/q_reg[0]  ( .D(\fpu_mul_ctl/n549 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/n264 ), .QN(n1058) );
  DFFX1 \fpu_mul_ctl/i_mul_exp_in2_exp_neq_ffs/q_reg[0]  ( .D(
        \fpu_mul_ctl/n548 ), .CLK(rclk), .Q(\fpu_mul_ctl/n253 ), .QN(n885) );
  DFFX1 \fpu_mul_ctl/i_m1stg_sngop/q_reg[0]  ( .D(\fpu_mul_ctl/n544 ), .CLK(
        rclk), .Q(m1stg_sngop) );
  DFFX1 \fpu_mul_ctl/i_m1stg_sngopa/q_reg[3]  ( .D(\fpu_mul_ctl/n543 ), .CLK(
        rclk), .Q(n1298) );
  DFFX1 \fpu_mul_ctl/i_m1stg_sngopa/q_reg[2]  ( .D(\fpu_mul_ctl/n542 ), .CLK(
        rclk), .Q(n1056), .QN(\fpu_mul_ctl/n259 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_sngopa/q_reg[1]  ( .D(\fpu_mul_ctl/n541 ), .CLK(
        rclk), .Q(n923), .QN(\fpu_mul_ctl/n116 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_sngopa/q_reg[0]  ( .D(\fpu_mul_ctl/n540 ), .CLK(
        rclk), .Q(n910), .QN(\fpu_mul_ctl/n117 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_dblop/q_reg[0]  ( .D(\fpu_mul_ctl/n539 ), .CLK(
        rclk), .Q(m1stg_dblop), .QN(n1031) );
  DFFX1 \fpu_mul_ctl/i_m1stg_dblopa/q_reg[3]  ( .D(\fpu_mul_ctl/n538 ), .CLK(
        rclk), .Q(n1299) );
  DFFX1 \fpu_mul_ctl/i_m1stg_dblopa/q_reg[2]  ( .D(\fpu_mul_ctl/n537 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/n265 ), .QN(n1338) );
  DFFX1 \fpu_mul_ctl/i_m1stg_dblopa/q_reg[1]  ( .D(\fpu_mul_ctl/n532 ), .CLK(
        rclk), .Q(n922), .QN(\fpu_mul_ctl/n120 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_dblopa/q_reg[0]  ( .D(\fpu_mul_ctl/n527 ), .CLK(
        rclk), .Q(n886) );
  DFFX1 \fpu_mul_ctl/i_m1stg_dblop_inv/q_reg[0]  ( .D(\fpu_mul_ctl/n526 ), 
        .CLK(rclk), .Q(m1stg_dblop_inv), .QN(n1032) );
  DFFX1 \fpu_mul_ctl/i_m5stg_rnd_mode/q_reg[1]  ( .D(\fpu_mul_ctl/n483 ), 
        .CLK(rclk), .Q(n926), .QN(\fpu_mul_ctl/n123 ) );
  DFFX1 \fpu_mul_ctl/i_m4stg_rnd_mode/q_reg[1]  ( .D(\fpu_mul_ctl/n490 ), 
        .CLK(rclk), .Q(n1250) );
  DFFX1 \fpu_mul_ctl/i_m3stg_rnd_mode/q_reg[1]  ( .D(\fpu_mul_ctl/n497 ), 
        .CLK(rclk), .Q(n1012) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_rnd_mode/q_reg[1]  ( .D(\fpu_mul_ctl/n504 ), 
        .CLK(rclk), .Q(n1245) );
  DFFX1 \fpu_mul_ctl/i_m3astg_rnd_mode/q_reg[1]  ( .D(\fpu_mul_ctl/n511 ), 
        .CLK(rclk), .Q(n1007) );
  DFFX1 \fpu_mul_ctl/i_m2stg_rnd_mode/q_reg[1]  ( .D(\fpu_mul_ctl/n518 ), 
        .CLK(rclk), .Q(n1240) );
  DFFX1 \fpu_mul_ctl/i_m1stg_rnd_mode/q_reg[1]  ( .D(\fpu_mul_ctl/n525 ), 
        .CLK(rclk), .Q(n1002) );
  DFFX1 \fpu_mul_ctl/i_m5stg_rnd_mode/q_reg[0]  ( .D(\fpu_mul_ctl/n482 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/m5stg_rnd_mode[0] ), .QN(
        \fpu_mul_ctl/n732 ) );
  DFFX1 \fpu_mul_ctl/i_m4stg_rnd_mode/q_reg[0]  ( .D(\fpu_mul_ctl/n489 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/m4stg_rnd_mode[0] ), .QN(
        \fpu_mul_ctl/n130 ) );
  DFFX1 \fpu_mul_ctl/i_m3stg_rnd_mode/q_reg[0]  ( .D(\fpu_mul_ctl/n496 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/m3stg_rnd_mode[0] ), .QN(
        \fpu_mul_ctl/n131 ) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_rnd_mode/q_reg[0]  ( .D(\fpu_mul_ctl/n503 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/m3bstg_rnd_mode[0] ), .QN(
        \fpu_mul_ctl/n132 ) );
  DFFX1 \fpu_mul_ctl/i_m3astg_rnd_mode/q_reg[0]  ( .D(\fpu_mul_ctl/n510 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/m3astg_rnd_mode[0] ), .QN(
        \fpu_mul_ctl/n133 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_rnd_mode/q_reg[0]  ( .D(\fpu_mul_ctl/n517 ), 
        .CLK(rclk), .Q(\fpu_mul_ctl/m2stg_rnd_mode[0] ), .QN(
        \fpu_mul_ctl/n134 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_rnd_mode/q_reg[0]  ( .D(\fpu_mul_ctl/n524 ), 
        .CLK(rclk), .Q(n1333), .QN(\fpu_mul_ctl/n135 ) );
  DFFX1 \fpu_mul_ctl/i_m5stg_id/q_reg[4]  ( .D(\fpu_mul_ctl/n481 ), .CLK(rclk), 
        .Q(\fpu_mul_ctl/m5stg_id[4] ), .QN(\fpu_mul_ctl/n136 ) );
  DFFX1 \fpu_mul_ctl/i_m4stg_id/q_reg[4]  ( .D(\fpu_mul_ctl/n488 ), .CLK(rclk), 
        .Q(\fpu_mul_ctl/m4stg_id[4] ), .QN(\fpu_mul_ctl/n137 ) );
  DFFX1 \fpu_mul_ctl/i_m3stg_id/q_reg[4]  ( .D(\fpu_mul_ctl/n495 ), .CLK(rclk), 
        .Q(\fpu_mul_ctl/m3stg_id[4] ), .QN(\fpu_mul_ctl/n138 ) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_id/q_reg[4]  ( .D(\fpu_mul_ctl/n502 ), .CLK(rclk), .Q(\fpu_mul_ctl/m3bstg_id[4] ), .QN(\fpu_mul_ctl/n139 ) );
  DFFX1 \fpu_mul_ctl/i_m3astg_id/q_reg[4]  ( .D(\fpu_mul_ctl/n509 ), .CLK(rclk), .Q(\fpu_mul_ctl/m3astg_id[4] ), .QN(\fpu_mul_ctl/n140 ) );
  DFFX1 \fpu_mul_ctl/i_m2stg_id/q_reg[4]  ( .D(\fpu_mul_ctl/n516 ), .CLK(rclk), 
        .Q(\fpu_mul_ctl/m2stg_id[4] ), .QN(\fpu_mul_ctl/n141 ) );
  DFFX1 \fpu_mul_ctl/i_m1stg_id/q_reg[4]  ( .D(\fpu_mul_ctl/n523 ), .CLK(rclk), 
        .Q(n1334), .QN(\fpu_mul_ctl/n142 ) );
  DFFX1 \fpu_mul_ctl/i_m5stg_id/q_reg[3]  ( .D(\fpu_mul_ctl/n480 ), .CLK(rclk), 
        .Q(n931), .QN(\fpu_mul_ctl/n143 ) );
  DFFX1 \fpu_mul_ctl/i_m4stg_id/q_reg[3]  ( .D(\fpu_mul_ctl/n487 ), .CLK(rclk), 
        .Q(n1251) );
  DFFX1 \fpu_mul_ctl/i_m3stg_id/q_reg[3]  ( .D(\fpu_mul_ctl/n494 ), .CLK(rclk), 
        .Q(n1013) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_id/q_reg[3]  ( .D(\fpu_mul_ctl/n501 ), .CLK(rclk), .Q(n1246) );
  DFFX1 \fpu_mul_ctl/i_m3astg_id/q_reg[3]  ( .D(\fpu_mul_ctl/n508 ), .CLK(rclk), .Q(n1008) );
  DFFX1 \fpu_mul_ctl/i_m2stg_id/q_reg[3]  ( .D(\fpu_mul_ctl/n515 ), .CLK(rclk), 
        .Q(n1241) );
  DFFX1 \fpu_mul_ctl/i_m1stg_id/q_reg[3]  ( .D(\fpu_mul_ctl/n522 ), .CLK(rclk), 
        .Q(n1003) );
  DFFX1 \fpu_mul_ctl/i_m5stg_id/q_reg[2]  ( .D(\fpu_mul_ctl/n479 ), .CLK(rclk), 
        .Q(n982), .QN(\fpu_mul_ctl/n260 ) );
  DFFX1 \fpu_mul_ctl/i_m4stg_id/q_reg[2]  ( .D(\fpu_mul_ctl/n486 ), .CLK(rclk), 
        .Q(n1252) );
  DFFX1 \fpu_mul_ctl/i_m3stg_id/q_reg[2]  ( .D(\fpu_mul_ctl/n493 ), .CLK(rclk), 
        .Q(n1014) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_id/q_reg[2]  ( .D(\fpu_mul_ctl/n500 ), .CLK(rclk), .Q(n1247) );
  DFFX1 \fpu_mul_ctl/i_m3astg_id/q_reg[2]  ( .D(\fpu_mul_ctl/n507 ), .CLK(rclk), .Q(n1009) );
  DFFX1 \fpu_mul_ctl/i_m2stg_id/q_reg[2]  ( .D(\fpu_mul_ctl/n514 ), .CLK(rclk), 
        .Q(n1242) );
  DFFX1 \fpu_mul_ctl/i_m1stg_id/q_reg[2]  ( .D(\fpu_mul_ctl/n521 ), .CLK(rclk), 
        .Q(n1004) );
  DFFX1 \fpu_mul_ctl/i_m5stg_id/q_reg[1]  ( .D(\fpu_mul_ctl/n478 ), .CLK(rclk), 
        .Q(n983), .QN(\fpu_mul_ctl/n156 ) );
  DFFX1 \fpu_mul_ctl/i_m4stg_id/q_reg[1]  ( .D(\fpu_mul_ctl/n485 ), .CLK(rclk), 
        .Q(n1253) );
  DFFX1 \fpu_mul_ctl/i_m3stg_id/q_reg[1]  ( .D(\fpu_mul_ctl/n492 ), .CLK(rclk), 
        .Q(n1015) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_id/q_reg[1]  ( .D(\fpu_mul_ctl/n499 ), .CLK(rclk), .Q(n1248) );
  DFFX1 \fpu_mul_ctl/i_m3astg_id/q_reg[1]  ( .D(\fpu_mul_ctl/n506 ), .CLK(rclk), .Q(n1010) );
  DFFX1 \fpu_mul_ctl/i_m2stg_id/q_reg[1]  ( .D(\fpu_mul_ctl/n513 ), .CLK(rclk), 
        .Q(n1243) );
  DFFX1 \fpu_mul_ctl/i_m1stg_id/q_reg[1]  ( .D(\fpu_mul_ctl/n520 ), .CLK(rclk), 
        .Q(n1005) );
  DFFX1 \fpu_mul_ctl/i_m5stg_id/q_reg[0]  ( .D(\fpu_mul_ctl/n477 ), .CLK(rclk), 
        .Q(n984), .QN(\fpu_mul_ctl/n163 ) );
  DFFX1 \fpu_mul_ctl/i_m4stg_id/q_reg[0]  ( .D(\fpu_mul_ctl/n484 ), .CLK(rclk), 
        .Q(n1254) );
  DFFX1 \fpu_mul_ctl/i_m3stg_id/q_reg[0]  ( .D(\fpu_mul_ctl/n491 ), .CLK(rclk), 
        .Q(n1016) );
  DFFX1 \fpu_mul_ctl/i_m3bstg_id/q_reg[0]  ( .D(\fpu_mul_ctl/n498 ), .CLK(rclk), .Q(n1249) );
  DFFX1 \fpu_mul_ctl/i_m3astg_id/q_reg[0]  ( .D(\fpu_mul_ctl/n505 ), .CLK(rclk), .Q(n1011) );
  DFFX1 \fpu_mul_ctl/i_m2stg_id/q_reg[0]  ( .D(\fpu_mul_ctl/n512 ), .CLK(rclk), 
        .Q(n1244) );
  DFFX1 \fpu_mul_ctl/i_m1stg_id/q_reg[0]  ( .D(\fpu_mul_ctl/n519 ), .CLK(rclk), 
        .Q(n1006) );
  DFFSSRX1 \fpu_mul_ctl/i_m6stg_opdec/q_reg[2]  ( .D(\fpu_mul_ctl/n735 ), 
        .RSTB(\fpu_mul_ctl/m5stg_opdec[4] ), .SETB(\fpu_mul_ctl/n105 ), .CLK(
        rclk), .Q(\fpu_mul_ctl/n261 ), .QN(n1223) );
  DFFARX1 \fpu_mul_ctl/dffrl_mul_ctl/q_reg[0]  ( .D(
        \fpu_mul_ctl/dffrl_mul_ctl/N4 ), .CLK(rclk), .RSTB(arst_l), .Q(n1209), 
        .QN(mul_rst_l) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[51]  ( .D(\fpu_mul_frac_dp/n922 ), .CLK(\fpu_mul_frac_dp/n832 ), .Q(mul_frac_out[51]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[50]  ( .D(\fpu_mul_frac_dp/n923 ), .CLK(n1581), .Q(mul_frac_out[50]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[49]  ( .D(\fpu_mul_frac_dp/n924 ), .CLK(n1582), .Q(mul_frac_out[49]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[48]  ( .D(\fpu_mul_frac_dp/n925 ), .CLK(n1583), .Q(mul_frac_out[48]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[47]  ( .D(\fpu_mul_frac_dp/n926 ), .CLK(n1560), .Q(mul_frac_out[47]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[46]  ( .D(\fpu_mul_frac_dp/n927 ), .CLK(n1560), .Q(mul_frac_out[46]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[45]  ( .D(\fpu_mul_frac_dp/n928 ), .CLK(n1560), .Q(mul_frac_out[45]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[44]  ( .D(\fpu_mul_frac_dp/n929 ), .CLK(n1560), .Q(mul_frac_out[44]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[43]  ( .D(\fpu_mul_frac_dp/n930 ), .CLK(n1560), .Q(mul_frac_out[43]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[42]  ( .D(\fpu_mul_frac_dp/n931 ), .CLK(n1560), .Q(mul_frac_out[42]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[41]  ( .D(\fpu_mul_frac_dp/n932 ), .CLK(n1560), .Q(mul_frac_out[41]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[40]  ( .D(\fpu_mul_frac_dp/n933 ), .CLK(n1560), .Q(mul_frac_out[40]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[39]  ( .D(\fpu_mul_frac_dp/n934 ), .CLK(n1560), .Q(mul_frac_out[39]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[38]  ( .D(\fpu_mul_frac_dp/n935 ), .CLK(n1560), .Q(mul_frac_out[38]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[37]  ( .D(\fpu_mul_frac_dp/n936 ), .CLK(n1560), .Q(mul_frac_out[37]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[36]  ( .D(\fpu_mul_frac_dp/n937 ), .CLK(n1560), .Q(mul_frac_out[36]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[35]  ( .D(\fpu_mul_frac_dp/n938 ), .CLK(n1559), .Q(mul_frac_out[35]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[34]  ( .D(\fpu_mul_frac_dp/n939 ), .CLK(n1559), .Q(mul_frac_out[34]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[33]  ( .D(\fpu_mul_frac_dp/n940 ), .CLK(n1559), .Q(mul_frac_out[33]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[32]  ( .D(\fpu_mul_frac_dp/n941 ), .CLK(n1559), .Q(mul_frac_out[32]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[31]  ( .D(\fpu_mul_frac_dp/n942 ), .CLK(n1559), .Q(mul_frac_out[31]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[30]  ( .D(\fpu_mul_frac_dp/n943 ), .CLK(n1559), .Q(mul_frac_out[30]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[29]  ( .D(\fpu_mul_frac_dp/n944 ), .CLK(n1559), .Q(mul_frac_out[29]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[28]  ( .D(\fpu_mul_frac_dp/n945 ), .CLK(n1557), .Q(mul_frac_out[28]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[27]  ( .D(\fpu_mul_frac_dp/n946 ), .CLK(n1557), .Q(mul_frac_out[27]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[26]  ( .D(\fpu_mul_frac_dp/n947 ), .CLK(n1557), .Q(mul_frac_out[26]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[25]  ( .D(\fpu_mul_frac_dp/n948 ), .CLK(n1557), .Q(mul_frac_out[25]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[24]  ( .D(\fpu_mul_frac_dp/n949 ), .CLK(n1557), .Q(mul_frac_out[24]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[23]  ( .D(\fpu_mul_frac_dp/n950 ), .CLK(n1557), .Q(mul_frac_out[23]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[22]  ( .D(\fpu_mul_frac_dp/n951 ), .CLK(n1557), .Q(mul_frac_out[22]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[21]  ( .D(\fpu_mul_frac_dp/n952 ), .CLK(n1557), .Q(mul_frac_out[21]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[20]  ( .D(\fpu_mul_frac_dp/n953 ), .CLK(n1557), .Q(mul_frac_out[20]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[19]  ( .D(\fpu_mul_frac_dp/n954 ), .CLK(n1557), .Q(mul_frac_out[19]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[18]  ( .D(\fpu_mul_frac_dp/n955 ), .CLK(n1557), .Q(mul_frac_out[18]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[17]  ( .D(\fpu_mul_frac_dp/n956 ), .CLK(n1557), .Q(mul_frac_out[17]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[16]  ( .D(\fpu_mul_frac_dp/n957 ), .CLK(n1558), .Q(mul_frac_out[16]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[15]  ( .D(\fpu_mul_frac_dp/n958 ), .CLK(n1558), .Q(mul_frac_out[15]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[14]  ( .D(\fpu_mul_frac_dp/n959 ), .CLK(n1558), .Q(mul_frac_out[14]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[13]  ( .D(\fpu_mul_frac_dp/n960 ), .CLK(n1558), .Q(mul_frac_out[13]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[12]  ( .D(\fpu_mul_frac_dp/n961 ), .CLK(n1558), .Q(mul_frac_out[12]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[11]  ( .D(\fpu_mul_frac_dp/n962 ), .CLK(n1558), .Q(mul_frac_out[11]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[10]  ( .D(\fpu_mul_frac_dp/n963 ), .CLK(n1558), .Q(mul_frac_out[10]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[9]  ( .D(\fpu_mul_frac_dp/n964 ), 
        .CLK(n1558), .Q(mul_frac_out[9]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[8]  ( .D(\fpu_mul_frac_dp/n965 ), 
        .CLK(n1558), .Q(mul_frac_out[8]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[7]  ( .D(\fpu_mul_frac_dp/n966 ), 
        .CLK(n1558), .Q(mul_frac_out[7]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[6]  ( .D(\fpu_mul_frac_dp/n967 ), 
        .CLK(n1558), .Q(mul_frac_out[6]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[5]  ( .D(\fpu_mul_frac_dp/n968 ), 
        .CLK(n1558), .Q(mul_frac_out[5]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[4]  ( .D(\fpu_mul_frac_dp/n969 ), 
        .CLK(n1559), .Q(mul_frac_out[4]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[3]  ( .D(\fpu_mul_frac_dp/n970 ), 
        .CLK(n1559), .Q(mul_frac_out[3]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[2]  ( .D(\fpu_mul_frac_dp/n971 ), 
        .CLK(n1559), .Q(mul_frac_out[2]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[1]  ( .D(\fpu_mul_frac_dp/n972 ), 
        .CLK(n1559), .Q(mul_frac_out[1]) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_out/q_reg[0]  ( .D(\fpu_mul_frac_dp/n973 ), 
        .CLK(n1559), .Q(mul_frac_out[0]) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[54]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N57 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[54] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[54]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N57 ), .CLK(n1578), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[54] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[53]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N56 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[53] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[53]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N56 ), .CLK(n1578), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[53] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[52]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N55 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[52] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[52]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N55 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[52] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[51]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N54 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[51] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[51]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N54 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[51] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[50]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N53 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[50] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[50]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N53 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[50] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[49]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N52 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[49] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[49]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N52 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[49] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[48]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N51 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[48] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[48]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N51 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[48] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[47]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N50 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[47] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[47]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N50 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[47] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[46]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N49 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[46] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[46]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N49 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[46] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[45]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N48 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[45] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[45]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N48 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[45] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[44]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N47 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[44] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[44]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N47 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[44] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[43]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N46 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[43] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[43]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N46 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[43] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[42]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N45 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[42] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[42]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N45 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[42] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[41]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N44 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[41] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[41]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N44 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[41] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[40]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N43 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[40] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[40]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N43 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[40] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[39]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N42 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[39] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[39]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N42 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[39] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[38]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N41 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[38] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[38]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N41 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[38] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[37]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N40 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[37] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[37]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N40 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[37] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[36]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N39 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[36] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[36]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N39 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[36] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[35]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N38 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[35] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[35]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N38 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[35] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[34]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N37 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[34] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[34]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N37 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[34] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[33]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N36 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[33] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[33]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N36 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[33] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[32]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N35 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[32] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[32]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N35 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[32] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[31]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N34 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[31] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[31]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N34 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[31] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[30]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N33 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[30] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[30]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N33 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[30] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[29]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N32 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[29] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[29]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N32 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[29] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[28]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N31 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[28] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[28]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N31 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[28] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[27]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N30 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[27] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[27]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N30 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[27] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[26]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N29 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[26] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[26]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N29 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[26] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[25]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N28 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[25] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[25]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N28 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[25] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[24]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N27 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[24] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[24]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N27 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[24] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[23]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N26 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[23] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[23]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N26 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[23] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[22]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N25 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[22] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[22]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N25 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[22] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[21]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N24 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[21] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[21]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N24 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[21] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[20]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N23 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[20] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[20]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N23 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[20] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[19]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N22 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[19] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[19]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N22 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[19] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[18]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N21 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[18] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[18]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N21 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[18] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[17]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N20 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[17] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[17]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N20 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[17] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[16]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N19 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[16] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[16]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N19 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[16] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[15]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N18 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[15] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[15]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N18 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[15] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[14]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N17 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[14] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[14]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N17 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[14] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[13]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N16 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[13] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[13]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N16 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[13] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[12]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N15 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[12] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[12]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N15 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[12] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[11]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N14 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[11] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[11]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N14 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[11] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[10]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N13 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[10] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[10]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N13 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[10] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[9]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N12 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[9] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[9]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N12 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[9] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[8]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N11 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[8] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[8]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N11 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[8] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[7]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N10 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[7] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[7]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N10 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[7] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[6]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N9 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[6] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[6]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N9 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[6] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[5]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N8 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[5] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[5]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N8 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[5] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[4]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N7 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[4] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[4]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N7 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[4] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[3]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N6 ), .CLK(\fpu_mul_frac_dp/n832 ), 
        .Q(\fpu_mul_frac_dp/m5stg_frac_pre1[3] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[3]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N6 ), .CLK(\fpu_mul_frac_dp/n832 ), 
        .Q(\fpu_mul_frac_dp/m5stg_frac_pre4[3] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[2]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N5 ), .CLK(\fpu_mul_frac_dp/n832 ), 
        .Q(\fpu_mul_frac_dp/m5stg_frac_pre1[2] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[2]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N5 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre4[2] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[1]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N4 ), .CLK(n1588), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre1[1] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[1]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N4 ), .CLK(\fpu_mul_frac_dp/n832 ), 
        .Q(\fpu_mul_frac_dp/m5stg_frac_pre4[1] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre1/q_reg[0]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N3 ), .CLK(\fpu_mul_frac_dp/n832 ), 
        .Q(\fpu_mul_frac_dp/m5stg_frac_pre1[0] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre4/q_reg[0]  ( .D(se_mul), .CLK(n1588), 
        .QN(\fpu_mul_frac_dp/m5stg_frac_pre4[0] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[54]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N57 ), .CLK(n1578), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[54] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[53]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N56 ), .CLK(n1578), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[53] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[52]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N55 ), .CLK(n1578), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[52] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[51]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N54 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[51] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[50]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N53 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[50] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[49]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N52 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[49] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[48]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N51 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[48] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[47]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N50 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[47] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[46]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N49 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[46] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[45]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N48 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[45] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[44]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N47 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[44] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[43]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N46 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[43] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[42]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N45 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[42] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[41]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N44 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[41] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[40]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N43 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[40] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[39]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N42 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[39] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[38]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N41 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[38] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[37]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N40 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[37] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[36]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N39 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[36] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[35]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N38 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[35] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[34]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N37 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[34] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[33]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N36 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[33] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[32]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N35 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[32] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[31]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N34 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[31] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[30]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N33 ), .CLK(n1564), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[30] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[29]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N32 ), .CLK(n1567), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[29] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[28]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N31 ), .CLK(n1570), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[28] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[27]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N30 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[27] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[26]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N29 ), .CLK(n1565), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[26] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[25]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N28 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[25] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[24]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N27 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[24] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[23]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N26 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[23] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[22]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N25 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[22] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[21]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N24 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[21] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[20]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N23 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[20] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[19]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N22 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[19] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[18]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N21 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[18] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[17]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N20 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[17] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[16]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N19 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[16] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[15]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N18 ), .CLK(n1571), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[15] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[14]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N17 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[14] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[13]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N16 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[13] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[12]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N15 ), .CLK(n1568), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[12] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[11]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N14 ), .CLK(n1572), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[11] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[10]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N13 ), .CLK(n1563), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[10] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[9]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N12 ), .CLK(n1566), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[9] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[8]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N11 ), .CLK(n1569), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[8] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[7]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N10 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[7] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[6]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N9 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[6] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[5]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N8 ), .CLK(n1562), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[5] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[4]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N7 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[4] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[3]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N6 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[3] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[2]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N5 ), .CLK(\fpu_mul_frac_dp/n832 ), 
        .Q(\fpu_mul_frac_dp/m5stg_frac_pre3[2] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[1]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N4 ), .CLK(n1561), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre3[1] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre3/q_reg[0]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N3 ), .CLK(\fpu_mul_frac_dp/n832 ), 
        .Q(\fpu_mul_frac_dp/m5stg_frac_pre3[0] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[54]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N57 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[54] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[53]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N56 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[53] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[52]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N55 ), .CLK(n1578), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[52] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[51]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N54 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[51] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[50]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N53 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[50] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[49]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N52 ), .CLK(n1573), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[49] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[48]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N51 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[48] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[47]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N50 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[47] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[46]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N49 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[46] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[45]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N48 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[45] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[44]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N47 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[44] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[43]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N46 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[43] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[42]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N45 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[42] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[41]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N44 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[41] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[40]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N43 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[40] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[39]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N42 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[39] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[38]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N41 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[38] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[37]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N40 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[37] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[36]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N39 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[36] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[35]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N38 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[35] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[34]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N37 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[34] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[33]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N36 ), .CLK(n1574), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[33] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[32]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N35 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[32] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[31]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N34 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[31] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[30]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N33 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[30] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[29]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N32 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[29] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[28]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N31 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[28] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[27]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N30 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[27] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[26]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N29 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[26] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[25]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N28 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[25] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[24]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N27 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[24] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[23]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N26 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[23] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[22]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N25 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[22] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[21]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N24 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[21] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[20]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N23 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[20] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[19]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N22 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[19] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[18]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N21 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[18] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[17]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N20 ), .CLK(n1575), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[17] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[16]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N19 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[16] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[15]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N18 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[15] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[14]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N17 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[14] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[13]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N16 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[13] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[12]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N15 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[12] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[11]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N14 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[11] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[10]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N13 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[10] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[9]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N12 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[9] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[8]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N11 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[8] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[7]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N10 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[7] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[6]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N9 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[6] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[5]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N8 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[5] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[4]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N7 ), .CLK(n1577), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[4] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[3]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N6 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[3] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[2]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N5 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[2] ) );
  DFFX1 \fpu_mul_frac_dp/i_m5stg_frac_pre2/q_reg[1]  ( .D(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N4 ), .CLK(n1576), .Q(
        \fpu_mul_frac_dp/m5stg_frac_pre2[1] ) );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[50]  ( .D(
        \fpu_mul_frac_dp/n974 ), .CLK(n1579), .Q(n1035), .QN(
        \fpu_mul_frac_dp/n766 ) );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[43]  ( .D(
        \fpu_mul_frac_dp/n975 ), .CLK(n1578), .Q(n1036), .QN(
        \fpu_mul_frac_dp/n767 ) );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[42]  ( .D(
        \fpu_mul_frac_dp/n976 ), .CLK(n1578), .Q(n908), .QN(
        \fpu_mul_frac_dp/n838 ) );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[41]  ( .D(
        \fpu_mul_frac_dp/n977 ), .CLK(n1578), .Q(n1033), .QN(
        \fpu_mul_frac_dp/n765 ) );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[40]  ( .D(
        \fpu_mul_frac_dp/n978 ), .CLK(n1578), .Q(n906), .QN(
        \fpu_mul_frac_dp/n833 ) );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[39]  ( .D(
        \fpu_mul_frac_dp/n979 ), .CLK(n1578), .Q(n879), .QN(
        \fpu_mul_frac_dp/n834 ) );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[38]  ( .D(
        \fpu_mul_frac_dp/n980 ), .CLK(n1578), .Q(n884), .QN(
        \fpu_mul_frac_dp/n831 ) );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[37]  ( .D(
        \fpu_mul_frac_dp/n981 ), .CLK(n1579), .Q(m3stg_ld0_inv[6]) );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[36]  ( .D(
        \fpu_mul_frac_dp/n982 ), .CLK(n1579), .Q(m3stg_ld0_inv[5]), .QN(n1279)
         );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[35]  ( .D(
        \fpu_mul_frac_dp/n983 ), .CLK(n1579), .Q(m3stg_ld0_inv[4]), .QN(n1059)
         );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[34]  ( .D(
        \fpu_mul_frac_dp/n984 ), .CLK(n1579), .Q(m3stg_ld0_inv[3]), .QN(n1280)
         );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[33]  ( .D(
        \fpu_mul_frac_dp/n985 ), .CLK(n1579), .Q(m3stg_ld0_inv[2]), .QN(n1150)
         );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[32]  ( .D(
        \fpu_mul_frac_dp/n986 ), .CLK(n1579), .Q(m3stg_ld0_inv[1]), .QN(n1051)
         );
  DFFX1 \fpu_mul_frac_dp/i_mstg_xtra_regs/q_reg[31]  ( .D(
        \fpu_mul_frac_dp/n987 ), .CLK(n1579), .Q(m3stg_ld0_inv[0]), .QN(n1340)
         );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[54]  ( .D(\fpu_mul_frac_dp/n988 ), .CLK(n1580), .Q(n1224), .QN(\fpu_mul_frac_dp/n286 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[53]  ( .D(\fpu_mul_frac_dp/n989 ), .CLK(n1580), .Q(n1151), .QN(\fpu_mul_frac_dp/n287 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[52]  ( .D(\fpu_mul_frac_dp/n990 ), .CLK(n1580), .Q(n942) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[51]  ( .D(\fpu_mul_frac_dp/n991 ), .CLK(n1580), .Q(n1132), .QN(\fpu_mul_frac_dp/n289 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[50]  ( .D(\fpu_mul_frac_dp/n992 ), .CLK(n1580), .Q(n916), .QN(\fpu_mul_frac_dp/n818 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[49]  ( .D(\fpu_mul_frac_dp/n993 ), .CLK(n1580), .Q(n891), .QN(\fpu_mul_frac_dp/n789 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[48]  ( .D(\fpu_mul_frac_dp/n994 ), .CLK(n1580), .Q(n1042), .QN(\fpu_mul_frac_dp/n761 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[47]  ( .D(\fpu_mul_frac_dp/n995 ), .CLK(n1580), .Q(n890), .QN(\fpu_mul_frac_dp/n753 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[46]  ( .D(\fpu_mul_frac_dp/n996 ), .CLK(n1579), .Q(n918), .QN(\fpu_mul_frac_dp/n811 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[45]  ( .D(\fpu_mul_frac_dp/n997 ), .CLK(n1579), .Q(n1044), .QN(\fpu_mul_frac_dp/n815 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[44]  ( .D(\fpu_mul_frac_dp/n998 ), .CLK(n1579), .Q(n880), .QN(\fpu_mul_frac_dp/n800 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[43]  ( .D(\fpu_mul_frac_dp/n999 ), .CLK(n1579), .Q(n917), .QN(\fpu_mul_frac_dp/n779 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[42]  ( .D(
        \fpu_mul_frac_dp/n1000 ), .CLK(n1588), .Q(n1047), .QN(
        \fpu_mul_frac_dp/n803 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[41]  ( .D(
        \fpu_mul_frac_dp/n1001 ), .CLK(n1588), .Q(n921), .QN(
        \fpu_mul_frac_dp/n782 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[40]  ( .D(
        \fpu_mul_frac_dp/n1002 ), .CLK(n1588), .Q(n1043), .QN(
        \fpu_mul_frac_dp/n300 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[39]  ( .D(
        \fpu_mul_frac_dp/n1003 ), .CLK(n1588), .Q(n889), .QN(
        \fpu_mul_frac_dp/n754 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[38]  ( .D(
        \fpu_mul_frac_dp/n1004 ), .CLK(n1588), .Q(n920), .QN(
        \fpu_mul_frac_dp/n812 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[37]  ( .D(
        \fpu_mul_frac_dp/n1005 ), .CLK(n1588), .Q(n1048), .QN(
        \fpu_mul_frac_dp/n303 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[36]  ( .D(
        \fpu_mul_frac_dp/n1006 ), .CLK(n1588), .Q(n909), .QN(
        \fpu_mul_frac_dp/n776 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[35]  ( .D(
        \fpu_mul_frac_dp/n1007 ), .CLK(n1588), .Q(n1046), .QN(
        \fpu_mul_frac_dp/n305 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[34]  ( .D(
        \fpu_mul_frac_dp/n1008 ), .CLK(n1588), .Q(n919), .QN(
        \fpu_mul_frac_dp/n306 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[33]  ( .D(
        \fpu_mul_frac_dp/n1009 ), .CLK(n1588), .Q(n1045), .QN(
        \fpu_mul_frac_dp/n307 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[32]  ( .D(
        \fpu_mul_frac_dp/n1010 ), .CLK(n1587), .Q(n887), .QN(
        \fpu_mul_frac_dp/n820 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[31]  ( .D(
        \fpu_mul_frac_dp/n1011 ), .CLK(n1587), .Q(n958), .QN(
        \fpu_mul_frac_dp/n309 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[30]  ( .D(
        \fpu_mul_frac_dp/n1012 ), .CLK(n1587), .Q(n1160), .QN(
        \fpu_mul_frac_dp/n310 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[29]  ( .D(
        \fpu_mul_frac_dp/n1013 ), .CLK(n1587), .Q(n959), .QN(
        \fpu_mul_frac_dp/n311 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[28]  ( .D(
        \fpu_mul_frac_dp/n1014 ), .CLK(n1587), .Q(\fpu_mul_frac_dp/n837 ), 
        .QN(\fpu_mul_frac_dp/n425 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[27]  ( .D(
        \fpu_mul_frac_dp/n1015 ), .CLK(n1587), .Q(n1148), .QN(
        \fpu_mul_frac_dp/n791 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[26]  ( .D(
        \fpu_mul_frac_dp/n1016 ), .CLK(n1587), .Q(n897), .QN(
        \fpu_mul_frac_dp/n819 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[25]  ( .D(
        \fpu_mul_frac_dp/n1017 ), .CLK(n1587), .Q(n957), .QN(
        \fpu_mul_frac_dp/n793 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[24]  ( .D(
        \fpu_mul_frac_dp/n1018 ), .CLK(n1587), .Q(n1157), .QN(
        \fpu_mul_frac_dp/n826 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[23]  ( .D(
        \fpu_mul_frac_dp/n1019 ), .CLK(n1587), .Q(n955), .QN(
        \fpu_mul_frac_dp/n775 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[22]  ( .D(
        \fpu_mul_frac_dp/n1020 ), .CLK(n1587), .Q(n1146), .QN(
        \fpu_mul_frac_dp/n809 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[21]  ( .D(
        \fpu_mul_frac_dp/n1021 ), .CLK(n1587), .Q(n940), .QN(
        \fpu_mul_frac_dp/n794 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[20]  ( .D(
        \fpu_mul_frac_dp/n1022 ), .CLK(n1586), .Q(n1156), .QN(
        \fpu_mul_frac_dp/n822 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[19]  ( .D(
        \fpu_mul_frac_dp/n1023 ), .CLK(n1586), .Q(n932), .QN(
        \fpu_mul_frac_dp/n780 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[18]  ( .D(
        \fpu_mul_frac_dp/n1024 ), .CLK(n1586), .Q(n1136), .QN(
        \fpu_mul_frac_dp/n804 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[17]  ( .D(
        \fpu_mul_frac_dp/n1025 ), .CLK(n1586), .Q(n930), .QN(
        \fpu_mul_frac_dp/n750 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[16]  ( .D(
        \fpu_mul_frac_dp/n1026 ), .CLK(n1586), .Q(n1141), .QN(
        \fpu_mul_frac_dp/n758 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[15]  ( .D(
        \fpu_mul_frac_dp/n1027 ), .CLK(n1586), .Q(n892), .QN(
        \fpu_mul_frac_dp/n783 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[14]  ( .D(
        \fpu_mul_frac_dp/n1028 ), .CLK(n1586), .Q(n1054), .QN(
        \fpu_mul_frac_dp/n817 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[13]  ( .D(
        \fpu_mul_frac_dp/n1029 ), .CLK(n1586), .Q(n927), .QN(
        \fpu_mul_frac_dp/n797 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[12]  ( .D(
        \fpu_mul_frac_dp/n1030 ), .CLK(n1586), .Q(n1113), .QN(
        \fpu_mul_frac_dp/n824 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[11]  ( .D(
        \fpu_mul_frac_dp/n1031 ), .CLK(n1586), .Q(n925), .QN(
        \fpu_mul_frac_dp/n788 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[10]  ( .D(
        \fpu_mul_frac_dp/n1032 ), .CLK(n1586), .Q(n881), .QN(
        \fpu_mul_frac_dp/n757 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[9]  ( .D(\fpu_mul_frac_dp/n1033 ), .CLK(n1586), .Q(n1137), .QN(\fpu_mul_frac_dp/n808 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[8]  ( .D(\fpu_mul_frac_dp/n1034 ), .CLK(n1585), .Q(n898), .QN(\fpu_mul_frac_dp/n777 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[7]  ( .D(\fpu_mul_frac_dp/n1035 ), .CLK(n1585), .Q(n953), .QN(\fpu_mul_frac_dp/n762 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[6]  ( .D(\fpu_mul_frac_dp/n1036 ), .CLK(n1585), .Q(n1149), .QN(\fpu_mul_frac_dp/n749 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[5]  ( .D(\fpu_mul_frac_dp/n1037 ), .CLK(n1585), .Q(n941), .QN(\fpu_mul_frac_dp/n801 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[4]  ( .D(\fpu_mul_frac_dp/n1038 ), .CLK(n1585), .Q(n1155), .QN(\fpu_mul_frac_dp/n784 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[3]  ( .D(\fpu_mul_frac_dp/n1039 ), .CLK(n1585), .Q(n896), .QN(\fpu_mul_frac_dp/n814 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[2]  ( .D(\fpu_mul_frac_dp/n1040 ), .CLK(n1585), .Q(n1147), .QN(\fpu_mul_frac_dp/n790 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[1]  ( .D(\fpu_mul_frac_dp/n1041 ), .CLK(n1585), .Q(n939), .QN(\fpu_mul_frac_dp/n816 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in2/q_reg[0]  ( .D(\fpu_mul_frac_dp/n1042 ), .CLK(n1585), .Q(n1158), .QN(\fpu_mul_frac_dp/n334 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[54]  ( .D(
        \fpu_mul_frac_dp/n1043 ), .CLK(n1585), .Q(n1200), .QN(
        \fpu_mul_frac_dp/n335 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[53]  ( .D(
        \fpu_mul_frac_dp/n1044 ), .CLK(n1585), .Q(n1315), .QN(
        \fpu_mul_frac_dp/n336 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[52]  ( .D(
        \fpu_mul_frac_dp/n1045 ), .CLK(n1585), .Q(n1318), .QN(
        \fpu_mul_frac_dp/n337 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[51]  ( .D(
        \fpu_mul_frac_dp/n1046 ), .CLK(n1584), .Q(n1124), .QN(
        \fpu_mul_frac_dp/n338 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[50]  ( .D(
        \fpu_mul_frac_dp/n1047 ), .CLK(n1584), .Q(n1301), .QN(
        \fpu_mul_frac_dp/n339 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[49]  ( .D(
        \fpu_mul_frac_dp/n1048 ), .CLK(n1584), .Q(n1306), .QN(
        \fpu_mul_frac_dp/n340 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[48]  ( .D(
        \fpu_mul_frac_dp/n1049 ), .CLK(n1584), .Q(n1195), .QN(
        \fpu_mul_frac_dp/n341 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[47]  ( .D(
        \fpu_mul_frac_dp/n1050 ), .CLK(n1584), .Q(n1193), .QN(
        \fpu_mul_frac_dp/n342 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[46]  ( .D(
        \fpu_mul_frac_dp/n1051 ), .CLK(n1584), .Q(n1300), .QN(
        \fpu_mul_frac_dp/n343 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[45]  ( .D(
        \fpu_mul_frac_dp/n1052 ), .CLK(n1584), .Q(n977), .QN(
        \fpu_mul_frac_dp/n344 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[44]  ( .D(
        \fpu_mul_frac_dp/n1053 ), .CLK(n1584), .Q(n973), .QN(
        \fpu_mul_frac_dp/n345 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[43]  ( .D(
        \fpu_mul_frac_dp/n1054 ), .CLK(n1584), .Q(n1305), .QN(
        \fpu_mul_frac_dp/n346 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[42]  ( .D(
        \fpu_mul_frac_dp/n1055 ), .CLK(n1584), .Q(n1304), .QN(
        \fpu_mul_frac_dp/n347 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[41]  ( .D(
        \fpu_mul_frac_dp/n1056 ), .CLK(n1584), .Q(n1309), .QN(
        \fpu_mul_frac_dp/n348 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[40]  ( .D(
        \fpu_mul_frac_dp/n1057 ), .CLK(n1584), .Q(n1308), .QN(
        \fpu_mul_frac_dp/n349 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[39]  ( .D(
        \fpu_mul_frac_dp/n1058 ), .CLK(n1583), .Q(n1187), .QN(
        \fpu_mul_frac_dp/n350 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[38]  ( .D(
        \fpu_mul_frac_dp/n1059 ), .CLK(n1583), .Q(n1303), .QN(
        \fpu_mul_frac_dp/n351 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[37]  ( .D(
        \fpu_mul_frac_dp/n1060 ), .CLK(n1583), .Q(n1307), .QN(
        \fpu_mul_frac_dp/n352 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[36]  ( .D(
        \fpu_mul_frac_dp/n1061 ), .CLK(n1583), .Q(n947), .QN(
        \fpu_mul_frac_dp/n353 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[35]  ( .D(
        \fpu_mul_frac_dp/n1062 ), .CLK(n1583), .Q(n1182), .QN(
        \fpu_mul_frac_dp/n354 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[34]  ( .D(
        \fpu_mul_frac_dp/n1063 ), .CLK(n1583), .Q(n1302), .QN(
        \fpu_mul_frac_dp/n355 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[33]  ( .D(
        \fpu_mul_frac_dp/n1064 ), .CLK(n1583), .Q(n1183), .QN(
        \fpu_mul_frac_dp/n356 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[32]  ( .D(
        \fpu_mul_frac_dp/n1065 ), .CLK(n1583), .Q(n967), .QN(
        \fpu_mul_frac_dp/n357 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[31]  ( .D(
        \fpu_mul_frac_dp/n1066 ), .CLK(n1583), .Q(n1319), .QN(
        \fpu_mul_frac_dp/n358 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[30]  ( .D(
        \fpu_mul_frac_dp/n1067 ), .CLK(n1583), .Q(n1320), .QN(
        \fpu_mul_frac_dp/n359 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[29]  ( .D(
        \fpu_mul_frac_dp/n1068 ), .CLK(n1583), .Q(n1326), .QN(
        \fpu_mul_frac_dp/n360 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[28]  ( .D(
        \fpu_mul_frac_dp/n1069 ), .CLK(n1583), .Q(\fpu_mul_frac_dp/n813 ), 
        .QN(n1207) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[27]  ( .D(
        \fpu_mul_frac_dp/n1070 ), .CLK(n1582), .Q(n986), .QN(
        \fpu_mul_frac_dp/n785 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[26]  ( .D(
        \fpu_mul_frac_dp/n1071 ), .CLK(n1582), .Q(n1220), .QN(
        \fpu_mul_frac_dp/n810 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[25]  ( .D(
        \fpu_mul_frac_dp/n1072 ), .CLK(n1582), .Q(n978), .QN(
        \fpu_mul_frac_dp/n796 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[24]  ( .D(
        \fpu_mul_frac_dp/n1073 ), .CLK(n1582), .Q(n1201), .QN(
        \fpu_mul_frac_dp/n823 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[23]  ( .D(
        \fpu_mul_frac_dp/n1074 ), .CLK(n1582), .Q(n987), .QN(
        \fpu_mul_frac_dp/n786 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[22]  ( .D(
        \fpu_mul_frac_dp/n1075 ), .CLK(n1582), .Q(n1221), .QN(
        \fpu_mul_frac_dp/n825 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[21]  ( .D(
        \fpu_mul_frac_dp/n1076 ), .CLK(n1582), .Q(n985), .QN(
        \fpu_mul_frac_dp/n763 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[20]  ( .D(
        \fpu_mul_frac_dp/n1077 ), .CLK(n1582), .Q(n1222), .QN(
        \fpu_mul_frac_dp/n829 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[19]  ( .D(
        \fpu_mul_frac_dp/n1078 ), .CLK(n1582), .Q(n882), .QN(
        \fpu_mul_frac_dp/n759 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[18]  ( .D(
        \fpu_mul_frac_dp/n1079 ), .CLK(n1582), .Q(n960), .QN(
        \fpu_mul_frac_dp/n805 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[17]  ( .D(
        \fpu_mul_frac_dp/n1080 ), .CLK(n1582), .Q(n899), .QN(
        \fpu_mul_frac_dp/n751 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[16]  ( .D(
        \fpu_mul_frac_dp/n1081 ), .CLK(n1582), .Q(n1159), .QN(
        \fpu_mul_frac_dp/n778 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[15]  ( .D(
        \fpu_mul_frac_dp/n1082 ), .CLK(n1581), .Q(n1202), .QN(
        \fpu_mul_frac_dp/n807 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[14]  ( .D(
        \fpu_mul_frac_dp/n1083 ), .CLK(n1581), .Q(n1310), .QN(
        \fpu_mul_frac_dp/n795 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[13]  ( .D(
        \fpu_mul_frac_dp/n1084 ), .CLK(n1581), .Q(n1314), .QN(
        \fpu_mul_frac_dp/n821 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[12]  ( .D(
        \fpu_mul_frac_dp/n1085 ), .CLK(n1581), .Q(\fpu_mul_frac_dp/n836 ), 
        .QN(n1283) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[11]  ( .D(
        \fpu_mul_frac_dp/n1086 ), .CLK(n1581), .Q(n1121), .QN(
        \fpu_mul_frac_dp/n760 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[10]  ( .D(
        \fpu_mul_frac_dp/n1087 ), .CLK(n1581), .Q(n1171), .QN(
        \fpu_mul_frac_dp/n802 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[9]  ( .D(\fpu_mul_frac_dp/n1088 ), .CLK(n1581), .Q(n952), .QN(\fpu_mul_frac_dp/n752 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[8]  ( .D(\fpu_mul_frac_dp/n1089 ), .CLK(n1581), .Q(n1186), .QN(\fpu_mul_frac_dp/n781 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[7]  ( .D(\fpu_mul_frac_dp/n1090 ), .CLK(n1581), .Q(n1317), .QN(\fpu_mul_frac_dp/n828 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[6]  ( .D(\fpu_mul_frac_dp/n1091 ), .CLK(n1581), .Q(n943), .QN(\fpu_mul_frac_dp/n787 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[5]  ( .D(\fpu_mul_frac_dp/n1092 ), .CLK(n1581), .Q(n1312), .QN(\fpu_mul_frac_dp/n756 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[4]  ( .D(\fpu_mul_frac_dp/n1093 ), .CLK(n1581), .Q(n1316), .QN(\fpu_mul_frac_dp/n806 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[3]  ( .D(\fpu_mul_frac_dp/n1094 ), .CLK(n1580), .Q(n1180), .QN(\fpu_mul_frac_dp/n764 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[2]  ( .D(\fpu_mul_frac_dp/n1095 ), .CLK(n1580), .Q(n1311), .QN(\fpu_mul_frac_dp/n792 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[1]  ( .D(\fpu_mul_frac_dp/n1096 ), .CLK(n1580), .Q(n956), .QN(\fpu_mul_frac_dp/n827 ) );
  DFFX1 \fpu_mul_frac_dp/i_mul_frac_in1/q_reg[0]  ( .D(\fpu_mul_frac_dp/n1097 ), .CLK(n1580), .Q(n1208), .QN(\fpu_mul_frac_dp/n382 ) );
  LATCHX1 \fpu_mul_frac_dp/ckbuf_mul_frac_dp/clken_reg  ( .CLK(n709), .D(
        \fpu_mul_frac_dp/ckbuf_mul_frac_dp/N1 ), .Q(
        \fpu_mul_frac_dp/ckbuf_mul_frac_dp/clken ), .QN(\fpu_mul_frac_dp/n383 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[67]  ( .D(\i_m4stg_frac/pcout_dff/N70 ), 
        .CLK(n1490), .Q(\i_m4stg_frac/pc[97] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[66]  ( .D(\i_m4stg_frac/pcout_dff/N69 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/pc[96] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[65]  ( .D(\i_m4stg_frac/pcout_dff/N68 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/pc[95] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[64]  ( .D(\i_m4stg_frac/pcout_dff/N67 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/pc[94] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[63]  ( .D(\i_m4stg_frac/pcout_dff/N66 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/pc[93] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[62]  ( .D(\i_m4stg_frac/pcout_dff/N65 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/pc[92] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[61]  ( .D(\i_m4stg_frac/pcout_dff/N64 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/pc[91] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[60]  ( .D(\i_m4stg_frac/pcout_dff/N63 ), 
        .CLK(n1489), .Q(\i_m4stg_frac/pc[90] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[59]  ( .D(\i_m4stg_frac/pcout_dff/N62 ), 
        .CLK(n1489), .Q(\i_m4stg_frac/pc[89] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[58]  ( .D(\i_m4stg_frac/pcout_dff/N61 ), 
        .CLK(n1500), .Q(\i_m4stg_frac/pc[88] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[57]  ( .D(\i_m4stg_frac/pcout_dff/N60 ), 
        .CLK(n1499), .Q(\i_m4stg_frac/pc[87] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[56]  ( .D(\i_m4stg_frac/pcout_dff/N59 ), 
        .CLK(n1486), .Q(\i_m4stg_frac/pc[86] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[55]  ( .D(\i_m4stg_frac/pcout_dff/N58 ), 
        .CLK(n1500), .Q(\i_m4stg_frac/pc[85] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[54]  ( .D(\i_m4stg_frac/pcout_dff/N57 ), 
        .CLK(n1501), .Q(\i_m4stg_frac/pc[84] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[53]  ( .D(\i_m4stg_frac/pcout_dff/N56 ), 
        .CLK(n1502), .Q(\i_m4stg_frac/pc[83] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[52]  ( .D(\i_m4stg_frac/pcout_dff/N55 ), 
        .CLK(n1503), .Q(\i_m4stg_frac/pc[82] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[51]  ( .D(\i_m4stg_frac/pcout_dff/N54 ), 
        .CLK(n1502), .Q(\i_m4stg_frac/pc[81] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[50]  ( .D(\i_m4stg_frac/pcout_dff/N53 ), 
        .CLK(n1501), .Q(\i_m4stg_frac/pc[80] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[49]  ( .D(\i_m4stg_frac/pcout_dff/N52 ), 
        .CLK(n1501), .Q(\i_m4stg_frac/pc[79] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[48]  ( .D(\i_m4stg_frac/pcout_dff/N51 ), 
        .CLK(n1502), .Q(\i_m4stg_frac/pc[78] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[47]  ( .D(\i_m4stg_frac/pcout_dff/N50 ), 
        .CLK(n1496), .Q(\i_m4stg_frac/pc[77] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[46]  ( .D(\i_m4stg_frac/pcout_dff/N49 ), 
        .CLK(n1493), .Q(\i_m4stg_frac/pc[76] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[45]  ( .D(\i_m4stg_frac/pcout_dff/N48 ), 
        .CLK(n1506), .Q(\i_m4stg_frac/pc[75] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[44]  ( .D(\i_m4stg_frac/pcout_dff/N47 ), 
        .CLK(n1506), .Q(\i_m4stg_frac/pc[74] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[43]  ( .D(\i_m4stg_frac/pcout_dff/N46 ), 
        .CLK(n1506), .Q(\i_m4stg_frac/pc[73] ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[42]  ( .D(\i_m4stg_frac/pcout_dff/N45 ), 
        .CLK(n1498), .Q(\i_m4stg_frac/pc[72] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[72]  ( .D(\i_m4stg_frac/n355 ), .CLK(
        n1498), .Q(\i_m4stg_frac/addin_cout[72] ), .QN(\i_m4stg_frac/n52 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[41]  ( .D(\i_m4stg_frac/pcout_dff/N44 ), 
        .CLK(n1498), .Q(\i_m4stg_frac/pc[71] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[71]  ( .D(\i_m4stg_frac/n357 ), .CLK(
        n1497), .Q(\i_m4stg_frac/addin_cout[71] ), .QN(\i_m4stg_frac/n54 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[40]  ( .D(\i_m4stg_frac/pcout_dff/N43 ), 
        .CLK(n1497), .Q(\i_m4stg_frac/pc[70] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[70]  ( .D(\i_m4stg_frac/n359 ), .CLK(
        n1497), .Q(\i_m4stg_frac/addin_cout[70] ), .QN(\i_m4stg_frac/n56 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[39]  ( .D(\i_m4stg_frac/pcout_dff/N42 ), 
        .CLK(n1496), .Q(\i_m4stg_frac/pc[69] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[69]  ( .D(\i_m4stg_frac/n495 ), .CLK(
        n1496), .Q(\i_m4stg_frac/addin_cout[69] ), .QN(\i_m4stg_frac/n58 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[38]  ( .D(\i_m4stg_frac/pcout_dff/N41 ), 
        .CLK(n1496), .Q(\i_m4stg_frac/pc[68] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[68]  ( .D(\i_m4stg_frac/n497 ), .CLK(
        n1495), .Q(\i_m4stg_frac/addin_cout[68] ), .QN(\i_m4stg_frac/n60 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[37]  ( .D(\i_m4stg_frac/pcout_dff/N40 ), 
        .CLK(n1495), .Q(\i_m4stg_frac/pc[67] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[67]  ( .D(\i_m4stg_frac/n499 ), .CLK(
        n1495), .Q(\i_m4stg_frac/addin_cout[67] ), .QN(\i_m4stg_frac/n62 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[36]  ( .D(\i_m4stg_frac/pcout_dff/N39 ), 
        .CLK(n1494), .Q(\i_m4stg_frac/pc[66] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[66]  ( .D(\i_m4stg_frac/n501 ), .CLK(
        n1494), .Q(\i_m4stg_frac/addin_cout[66] ), .QN(\i_m4stg_frac/n64 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[35]  ( .D(\i_m4stg_frac/pcout_dff/N38 ), 
        .CLK(n1493), .Q(\i_m4stg_frac/pc[65] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[65]  ( .D(\i_m4stg_frac/n503 ), .CLK(
        n1493), .Q(\i_m4stg_frac/addin_cout[65] ), .QN(\i_m4stg_frac/n66 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[34]  ( .D(\i_m4stg_frac/pcout_dff/N37 ), 
        .CLK(n1492), .Q(\i_m4stg_frac/pc[64] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[64]  ( .D(\i_m4stg_frac/n505 ), .CLK(
        n1492), .Q(\i_m4stg_frac/addin_cout[64] ), .QN(\i_m4stg_frac/n68 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[33]  ( .D(\i_m4stg_frac/pcout_dff/N36 ), 
        .CLK(n1492), .Q(\i_m4stg_frac/pc[63] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[63]  ( .D(\i_m4stg_frac/n507 ), .CLK(
        n1492), .Q(\i_m4stg_frac/addin_cout[63] ), .QN(\i_m4stg_frac/n70 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[32]  ( .D(\i_m4stg_frac/pcout_dff/N35 ), 
        .CLK(n1491), .Q(\i_m4stg_frac/pc[62] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[62]  ( .D(\i_m4stg_frac/n509 ), .CLK(
        n1491), .Q(\i_m4stg_frac/addin_cout[62] ), .QN(\i_m4stg_frac/n72 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[31]  ( .D(\i_m4stg_frac/pcout_dff/N34 ), 
        .CLK(n1491), .Q(\i_m4stg_frac/pc[61] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[61]  ( .D(\i_m4stg_frac/n511 ), .CLK(
        n1491), .Q(\i_m4stg_frac/addin_cout[61] ), .QN(\i_m4stg_frac/n74 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[30]  ( .D(\i_m4stg_frac/pcout_dff/N33 ), 
        .CLK(n1499), .Q(\i_m4stg_frac/pc[60] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[60]  ( .D(\i_m4stg_frac/n513 ), .CLK(
        n1499), .Q(\i_m4stg_frac/addin_cout[60] ), .QN(\i_m4stg_frac/n76 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[29]  ( .D(\i_m4stg_frac/pcout_dff/N32 ), 
        .CLK(n1499), .Q(\i_m4stg_frac/pc[59] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[59]  ( .D(\i_m4stg_frac/n515 ), .CLK(
        n1499), .Q(\i_m4stg_frac/addin_cout[59] ), .QN(\i_m4stg_frac/n78 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[28]  ( .D(\i_m4stg_frac/pcout_dff/N31 ), 
        .CLK(n1485), .Q(\i_m4stg_frac/pc[58] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[58]  ( .D(\i_m4stg_frac/n517 ), .CLK(
        n1485), .Q(\i_m4stg_frac/addin_cout[58] ), .QN(\i_m4stg_frac/n80 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[27]  ( .D(\i_m4stg_frac/pcout_dff/N30 ), 
        .CLK(n1484), .Q(\i_m4stg_frac/pc[57] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[57]  ( .D(\i_m4stg_frac/n519 ), .CLK(
        n1485), .Q(\i_m4stg_frac/addin_cout[57] ), .QN(\i_m4stg_frac/n82 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[26]  ( .D(\i_m4stg_frac/pcout_dff/N29 ), 
        .CLK(n1483), .Q(\i_m4stg_frac/pc[56] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[56]  ( .D(\i_m4stg_frac/n521 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_cout[56] ), .QN(\i_m4stg_frac/n84 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[25]  ( .D(\i_m4stg_frac/pcout_dff/N28 ), 
        .CLK(n1483), .Q(\i_m4stg_frac/pc[55] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[55]  ( .D(\i_m4stg_frac/n523 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_cout[55] ), .QN(\i_m4stg_frac/n86 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[24]  ( .D(\i_m4stg_frac/pcout_dff/N27 ), 
        .CLK(n1485), .Q(\i_m4stg_frac/pc[54] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[54]  ( .D(\i_m4stg_frac/n525 ), .CLK(
        n1485), .Q(\i_m4stg_frac/addin_cout[54] ), .QN(\i_m4stg_frac/n88 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[23]  ( .D(\i_m4stg_frac/pcout_dff/N26 ), 
        .CLK(n1500), .Q(\i_m4stg_frac/pc[53] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[53]  ( .D(\i_m4stg_frac/n527 ), .CLK(
        n1500), .Q(\i_m4stg_frac/addin_cout[53] ), .QN(\i_m4stg_frac/n90 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[22]  ( .D(\i_m4stg_frac/pcout_dff/N25 ), 
        .CLK(n1501), .Q(\i_m4stg_frac/pc[52] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[52]  ( .D(\i_m4stg_frac/n529 ), .CLK(
        n1501), .Q(\i_m4stg_frac/addin_cout[52] ), .QN(\i_m4stg_frac/n92 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[21]  ( .D(\i_m4stg_frac/pcout_dff/N24 ), 
        .CLK(n1502), .Q(\i_m4stg_frac/pc[51] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[51]  ( .D(\i_m4stg_frac/n531 ), .CLK(
        n1502), .Q(\i_m4stg_frac/addin_cout[51] ), .QN(\i_m4stg_frac/n94 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[20]  ( .D(\i_m4stg_frac/pcout_dff/N23 ), 
        .CLK(n1502), .Q(\i_m4stg_frac/pc[50] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[50]  ( .D(\i_m4stg_frac/n533 ), .CLK(
        n1503), .Q(\i_m4stg_frac/addin_cout[50] ), .QN(\i_m4stg_frac/n96 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[19]  ( .D(\i_m4stg_frac/pcout_dff/N22 ), 
        .CLK(n1494), .Q(\i_m4stg_frac/pc[49] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[49]  ( .D(\i_m4stg_frac/n535 ), .CLK(
        n1495), .Q(\i_m4stg_frac/addin_cout[49] ), .QN(\i_m4stg_frac/n98 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[18]  ( .D(\i_m4stg_frac/pcout_dff/N21 ), 
        .CLK(n1492), .Q(\i_m4stg_frac/pc[48] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[48]  ( .D(\i_m4stg_frac/n537 ), .CLK(
        n1493), .Q(\i_m4stg_frac/addin_cout[48] ), .QN(\i_m4stg_frac/n100 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[17]  ( .D(\i_m4stg_frac/pcout_dff/N20 ), 
        .CLK(n1506), .Q(\i_m4stg_frac/pc[47] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[47]  ( .D(\i_m4stg_frac/n539 ), .CLK(
        n1506), .Q(\i_m4stg_frac/addin_cout[47] ), .QN(\i_m4stg_frac/n102 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[16]  ( .D(\i_m4stg_frac/pcout_dff/N19 ), 
        .CLK(n1505), .Q(\i_m4stg_frac/pc[46] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[46]  ( .D(\i_m4stg_frac/n541 ), .CLK(
        n1505), .Q(\i_m4stg_frac/addin_cout[46] ), .QN(\i_m4stg_frac/n104 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[15]  ( .D(\i_m4stg_frac/pcout_dff/N18 ), 
        .CLK(n1504), .Q(\i_m4stg_frac/pc[45] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[45]  ( .D(\i_m4stg_frac/n543 ), .CLK(
        n1504), .Q(\i_m4stg_frac/addin_cout[45] ), .QN(\i_m4stg_frac/n106 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[14]  ( .D(\i_m4stg_frac/pcout_dff/N17 ), 
        .CLK(n1504), .Q(\i_m4stg_frac/pc[44] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[44]  ( .D(\i_m4stg_frac/n545 ), .CLK(
        n1504), .Q(\i_m4stg_frac/addin_cout[44] ), .QN(\i_m4stg_frac/n108 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[13]  ( .D(\i_m4stg_frac/pcout_dff/N16 ), 
        .CLK(n1503), .Q(\i_m4stg_frac/pc[43] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[43]  ( .D(\i_m4stg_frac/n547 ), .CLK(
        n1504), .Q(\i_m4stg_frac/addin_cout[43] ), .QN(\i_m4stg_frac/n110 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[12]  ( .D(\i_m4stg_frac/pcout_dff/N15 ), 
        .CLK(n1505), .Q(\i_m4stg_frac/pc[42] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[42]  ( .D(\i_m4stg_frac/n549 ), .CLK(
        n1505), .Q(\i_m4stg_frac/addin_cout[42] ), .QN(\i_m4stg_frac/n112 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[11]  ( .D(\i_m4stg_frac/pcout_dff/N14 ), 
        .CLK(n1491), .Q(\i_m4stg_frac/pc[41] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[41]  ( .D(\i_m4stg_frac/n551 ), .CLK(
        n1495), .Q(\i_m4stg_frac/addin_cout[41] ), .QN(\i_m4stg_frac/n114 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[10]  ( .D(\i_m4stg_frac/pcout_dff/N13 ), 
        .CLK(n1496), .Q(\i_m4stg_frac/pc[40] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[40]  ( .D(\i_m4stg_frac/n553 ), .CLK(
        n1497), .Q(\i_m4stg_frac/addin_cout[40] ), .QN(\i_m4stg_frac/n116 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[9]  ( .D(\i_m4stg_frac/pcout_dff/N12 ), 
        .CLK(n1498), .Q(\i_m4stg_frac/pc[39] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[39]  ( .D(\i_m4stg_frac/n555 ), .CLK(
        n1498), .Q(\i_m4stg_frac/addin_cout[39] ), .QN(\i_m4stg_frac/n118 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[8]  ( .D(\i_m4stg_frac/pcout_dff/N11 ), 
        .CLK(n1497), .Q(\i_m4stg_frac/pc[38] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[38]  ( .D(\i_m4stg_frac/n557 ), .CLK(
        n1497), .Q(\i_m4stg_frac/addin_cout[38] ), .QN(\i_m4stg_frac/n120 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[7]  ( .D(\i_m4stg_frac/pcout_dff/N10 ), 
        .CLK(n1496), .Q(\i_m4stg_frac/pc[37] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[37]  ( .D(\i_m4stg_frac/n559 ), .CLK(
        n1496), .Q(\i_m4stg_frac/addin_cout[37] ), .QN(\i_m4stg_frac/n122 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[6]  ( .D(\i_m4stg_frac/pcout_dff/N9 ), 
        .CLK(n1495), .Q(\i_m4stg_frac/pc[36] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[36]  ( .D(\i_m4stg_frac/n561 ), .CLK(
        n1495), .Q(\i_m4stg_frac/addin_cout[36] ), .QN(\i_m4stg_frac/n124 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[5]  ( .D(\i_m4stg_frac/pcout_dff/N8 ), 
        .CLK(n1494), .Q(\i_m4stg_frac/pc[35] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[35]  ( .D(\i_m4stg_frac/n563 ), .CLK(
        n1494), .Q(\i_m4stg_frac/addin_cout[35] ), .QN(\i_m4stg_frac/n126 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[4]  ( .D(\i_m4stg_frac/pcout_dff/N7 ), 
        .CLK(n1494), .Q(\i_m4stg_frac/pc[34] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[34]  ( .D(\i_m4stg_frac/n565 ), .CLK(
        n1494), .Q(\i_m4stg_frac/addin_cout[34] ), .QN(\i_m4stg_frac/n128 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[3]  ( .D(\i_m4stg_frac/pcout_dff/N6 ), 
        .CLK(n1493), .Q(\i_m4stg_frac/pc[33] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[33]  ( .D(\i_m4stg_frac/n567 ), .CLK(
        n1493), .Q(\i_m4stg_frac/addin_cout[33] ), .QN(\i_m4stg_frac/n130 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[2]  ( .D(\i_m4stg_frac/pcout_dff/N5 ), 
        .CLK(n1499), .Q(\i_m4stg_frac/pc[32] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[32]  ( .D(\i_m4stg_frac/n569 ), .CLK(
        n1499), .Q(\i_m4stg_frac/addin_cout[32] ), .QN(\i_m4stg_frac/n132 ) );
  DFFX1 \i_m4stg_frac/pcout_dff/q_reg[1]  ( .D(\i_m4stg_frac/pcout_dff/N4 ), 
        .CLK(n1486), .Q(\i_m4stg_frac/pc[31] ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[31]  ( .D(\i_m4stg_frac/n571 ), .CLK(
        n1486), .Q(\i_m4stg_frac/addin_cout[31] ), .QN(\i_m4stg_frac/n134 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[30]  ( .D(\i_m4stg_frac/n573 ), .CLK(
        n1485), .Q(\i_m4stg_frac/addin_cout[30] ), .QN(\i_m4stg_frac/n136 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[29]  ( .D(\i_m4stg_frac/n575 ), .CLK(
        n1485), .Q(\i_m4stg_frac/addin_cout[29] ), .QN(\i_m4stg_frac/n137 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[28]  ( .D(\i_m4stg_frac/n577 ), .CLK(
        n1483), .Q(\i_m4stg_frac/addin_cout[28] ), .QN(\i_m4stg_frac/n138 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[27]  ( .D(\i_m4stg_frac/n579 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_cout[27] ), .QN(\i_m4stg_frac/n139 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[26]  ( .D(\i_m4stg_frac/n581 ), .CLK(
        n1483), .Q(\i_m4stg_frac/addin_cout[26] ), .QN(\i_m4stg_frac/n140 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[25]  ( .D(\i_m4stg_frac/n583 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_cout[25] ), .QN(\i_m4stg_frac/n141 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[24]  ( .D(\i_m4stg_frac/n585 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_cout[24] ), .QN(\i_m4stg_frac/n142 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[23]  ( .D(\i_m4stg_frac/n587 ), .CLK(
        n1483), .Q(\i_m4stg_frac/addin_cout[23] ), .QN(\i_m4stg_frac/n143 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[22]  ( .D(\i_m4stg_frac/n589 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_cout[22] ), .QN(\i_m4stg_frac/n144 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[21]  ( .D(\i_m4stg_frac/n443 ), .CLK(
        n1500), .Q(\i_m4stg_frac/addin_cout[21] ), .QN(\i_m4stg_frac/n145 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[20]  ( .D(\i_m4stg_frac/n591 ), .CLK(
        n1501), .Q(\i_m4stg_frac/addin_cout[20] ), .QN(\i_m4stg_frac/n146 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[19]  ( .D(\i_m4stg_frac/n593 ), .CLK(
        n1502), .Q(\i_m4stg_frac/addin_cout[19] ), .QN(\i_m4stg_frac/n147 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[18]  ( .D(\i_m4stg_frac/n595 ), .CLK(
        n1503), .Q(\i_m4stg_frac/addin_cout[18] ), .QN(\i_m4stg_frac/n148 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[17]  ( .D(\i_m4stg_frac/n597 ), .CLK(
        n1505), .Q(\i_m4stg_frac/addin_cout[17] ), .QN(\i_m4stg_frac/n149 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[16]  ( .D(\i_m4stg_frac/a2cot_dff/N19 ), 
        .CLK(n1504), .Q(\i_m4stg_frac/addin_cout[16] ), .QN(
        \i_m4stg_frac/n150 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[14]  ( .D(\i_m4stg_frac/n599 ), .CLK(
        n1503), .Q(\i_m4stg_frac/addin_cout[14] ), .QN(\i_m4stg_frac/n152 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[13]  ( .D(\i_m4stg_frac/n601 ), .CLK(
        n1503), .Q(\i_m4stg_frac/addin_cout[13] ), .QN(\i_m4stg_frac/n153 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[12]  ( .D(\i_m4stg_frac/n603 ), .CLK(
        n1503), .Q(\i_m4stg_frac/addin_cout[12] ), .QN(\i_m4stg_frac/n154 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[11]  ( .D(\i_m4stg_frac/n605 ), .CLK(
        n1504), .Q(\i_m4stg_frac/addin_cout[11] ), .QN(\i_m4stg_frac/n155 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[10]  ( .D(\i_m4stg_frac/n607 ), .CLK(
        n1505), .Q(\i_m4stg_frac/addin_cout[10] ), .QN(\i_m4stg_frac/n156 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[9]  ( .D(\i_m4stg_frac/n635 ), .CLK(
        n1491), .Q(\i_m4stg_frac/addin_cout[9] ), .QN(\i_m4stg_frac/n157 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[8]  ( .D(\i_m4stg_frac/n637 ), .CLK(
        n1497), .Q(\i_m4stg_frac/addin_cout[8] ), .QN(\i_m4stg_frac/n158 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[7]  ( .D(\i_m4stg_frac/n621 ), .CLK(
        n1498), .Q(\i_m4stg_frac/addin_cout[7] ), .QN(\i_m4stg_frac/n159 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[6]  ( .D(\i_m4stg_frac/n493 ), .CLK(
        n1497), .Q(\i_m4stg_frac/addin_cout[6] ), .QN(\i_m4stg_frac/n160 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[5]  ( .D(\i_m4stg_frac/n445 ), .CLK(
        n1496), .Q(\i_m4stg_frac/addin_cout[5] ), .QN(\i_m4stg_frac/n161 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[4]  ( .D(\i_m4stg_frac/n361 ), .CLK(
        n1495), .Q(\i_m4stg_frac/addin_cout[4] ), .QN(\i_m4stg_frac/n162 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[3]  ( .D(\i_m4stg_frac/n363 ), .CLK(
        n1499), .Q(\i_m4stg_frac/addin_cout[3] ), .QN(\i_m4stg_frac/n163 ) );
  DFFX1 \i_m4stg_frac/a2cot_dff/q_reg[2]  ( .D(\i_m4stg_frac/n365 ), .CLK(
        n1486), .Q(\i_m4stg_frac/addin_cout[2] ), .QN(\i_m4stg_frac/n164 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[67]  ( .D(\i_m4stg_frac/psum_dff/N70 ), 
        .CLK(n1490), .Q(\i_m4stg_frac/ps[98] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[66]  ( .D(\i_m4stg_frac/psum_dff/N69 ), 
        .CLK(n1490), .Q(\i_m4stg_frac/ps[97] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[65]  ( .D(\i_m4stg_frac/psum_dff/N68 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/ps[96] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[64]  ( .D(\i_m4stg_frac/psum_dff/N67 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/ps[95] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[63]  ( .D(\i_m4stg_frac/psum_dff/N66 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/ps[94] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[62]  ( .D(\i_m4stg_frac/psum_dff/N65 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/ps[93] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[61]  ( .D(\i_m4stg_frac/psum_dff/N64 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/ps[92] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[60]  ( .D(\i_m4stg_frac/psum_dff/N63 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/ps[91] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[59]  ( .D(\i_m4stg_frac/psum_dff/N62 ), 
        .CLK(n1488), .Q(\i_m4stg_frac/ps[90] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[58]  ( .D(\i_m4stg_frac/psum_dff/N61 ), 
        .CLK(n1489), .Q(\i_m4stg_frac/ps[89] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[57]  ( .D(\i_m4stg_frac/psum_dff/N60 ), 
        .CLK(n1499), .Q(\i_m4stg_frac/ps[88] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[56]  ( .D(\i_m4stg_frac/psum_dff/N59 ), 
        .CLK(n1486), .Q(\i_m4stg_frac/ps[87] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[55]  ( .D(\i_m4stg_frac/psum_dff/N58 ), 
        .CLK(n1485), .Q(\i_m4stg_frac/ps[86] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[54]  ( .D(\i_m4stg_frac/psum_dff/N57 ), 
        .CLK(n1500), .Q(\i_m4stg_frac/ps[85] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[53]  ( .D(\i_m4stg_frac/psum_dff/N56 ), 
        .CLK(n1501), .Q(\i_m4stg_frac/ps[84] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[52]  ( .D(\i_m4stg_frac/psum_dff/N55 ), 
        .CLK(n1502), .Q(\i_m4stg_frac/ps[83] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[51]  ( .D(\i_m4stg_frac/psum_dff/N54 ), 
        .CLK(n1503), .Q(\i_m4stg_frac/ps[82] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[50]  ( .D(\i_m4stg_frac/psum_dff/N53 ), 
        .CLK(n1502), .Q(\i_m4stg_frac/ps[81] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[49]  ( .D(\i_m4stg_frac/psum_dff/N52 ), 
        .CLK(n1501), .Q(\i_m4stg_frac/ps[80] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[48]  ( .D(\i_m4stg_frac/psum_dff/N51 ), 
        .CLK(n1501), .Q(\i_m4stg_frac/ps[79] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[47]  ( .D(\i_m4stg_frac/psum_dff/N50 ), 
        .CLK(n1502), .Q(\i_m4stg_frac/ps[78] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[46]  ( .D(\i_m4stg_frac/psum_dff/N49 ), 
        .CLK(n1494), .Q(\i_m4stg_frac/ps[77] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[45]  ( .D(\i_m4stg_frac/psum_dff/N48 ), 
        .CLK(n1492), .Q(\i_m4stg_frac/ps[76] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[44]  ( .D(\i_m4stg_frac/psum_dff/N47 ), 
        .CLK(n1506), .Q(\i_m4stg_frac/ps[75] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[43]  ( .D(\i_m4stg_frac/psum_dff/N46 ), 
        .CLK(n1505), .Q(\i_m4stg_frac/ps[74] ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[42]  ( .D(\i_m4stg_frac/psum_dff/N45 ), 
        .CLK(n1492), .Q(\i_m4stg_frac/ps[73] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[73]  ( .D(\i_m4stg_frac/n623 ), .CLK(
        n1492), .Q(\i_m4stg_frac/addin_sum[73] ), .QN(\i_m4stg_frac/n217 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[41]  ( .D(\i_m4stg_frac/psum_dff/N44 ), 
        .CLK(n1486), .Q(\i_m4stg_frac/ps[72] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[72]  ( .D(\i_m4stg_frac/n625 ), .CLK(
        n1498), .Q(\i_m4stg_frac/addin_sum[72] ), .QN(\i_m4stg_frac/n219 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[40]  ( .D(\i_m4stg_frac/psum_dff/N43 ), 
        .CLK(n1498), .Q(\i_m4stg_frac/ps[71] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[71]  ( .D(\i_m4stg_frac/n627 ), .CLK(
        n1498), .Q(\i_m4stg_frac/addin_sum[71] ), .QN(\i_m4stg_frac/n221 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[39]  ( .D(\i_m4stg_frac/psum_dff/N42 ), 
        .CLK(n1497), .Q(\i_m4stg_frac/ps[70] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[70]  ( .D(\i_m4stg_frac/n629 ), .CLK(
        n1497), .Q(\i_m4stg_frac/addin_sum[70] ), .QN(\i_m4stg_frac/n223 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[38]  ( .D(\i_m4stg_frac/psum_dff/N41 ), 
        .CLK(n1496), .Q(\i_m4stg_frac/ps[69] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[69]  ( .D(\i_m4stg_frac/n441 ), .CLK(
        n1496), .Q(\i_m4stg_frac/addin_sum[69] ), .QN(\i_m4stg_frac/n225 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[37]  ( .D(\i_m4stg_frac/psum_dff/N40 ), 
        .CLK(n1495), .Q(\i_m4stg_frac/ps[68] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[68]  ( .D(\i_m4stg_frac/n367 ), .CLK(
        n1495), .Q(\i_m4stg_frac/addin_sum[68] ), .QN(\i_m4stg_frac/n227 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[36]  ( .D(\i_m4stg_frac/psum_dff/N39 ), 
        .CLK(n1494), .Q(\i_m4stg_frac/ps[67] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[67]  ( .D(\i_m4stg_frac/n369 ), .CLK(
        n1494), .Q(\i_m4stg_frac/addin_sum[67] ), .QN(\i_m4stg_frac/n229 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[35]  ( .D(\i_m4stg_frac/psum_dff/N38 ), 
        .CLK(n1493), .Q(\i_m4stg_frac/ps[66] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[66]  ( .D(\i_m4stg_frac/n371 ), .CLK(
        n1493), .Q(\i_m4stg_frac/addin_sum[66] ), .QN(\i_m4stg_frac/n231 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[34]  ( .D(\i_m4stg_frac/psum_dff/N37 ), 
        .CLK(n1493), .Q(\i_m4stg_frac/ps[65] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[65]  ( .D(\i_m4stg_frac/n373 ), .CLK(
        n1493), .Q(\i_m4stg_frac/addin_sum[65] ), .QN(\i_m4stg_frac/n233 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[33]  ( .D(\i_m4stg_frac/psum_dff/N36 ), 
        .CLK(n1492), .Q(\i_m4stg_frac/ps[64] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[64]  ( .D(\i_m4stg_frac/n375 ), .CLK(
        n1492), .Q(\i_m4stg_frac/addin_sum[64] ), .QN(\i_m4stg_frac/n235 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[32]  ( .D(\i_m4stg_frac/psum_dff/N35 ), 
        .CLK(n1492), .Q(\i_m4stg_frac/ps[63] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[63]  ( .D(\i_m4stg_frac/n377 ), .CLK(
        n1492), .Q(\i_m4stg_frac/addin_sum[63] ), .QN(\i_m4stg_frac/n237 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[31]  ( .D(\i_m4stg_frac/psum_dff/N34 ), 
        .CLK(n1491), .Q(\i_m4stg_frac/ps[62] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[62]  ( .D(\i_m4stg_frac/n379 ), .CLK(
        n1491), .Q(\i_m4stg_frac/addin_sum[62] ), .QN(\i_m4stg_frac/n239 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[30]  ( .D(\i_m4stg_frac/psum_dff/N33 ), 
        .CLK(n1491), .Q(\i_m4stg_frac/ps[61] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[61]  ( .D(\i_m4stg_frac/n381 ), .CLK(
        n1491), .Q(\i_m4stg_frac/addin_sum[61] ), .QN(\i_m4stg_frac/n241 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[29]  ( .D(\i_m4stg_frac/psum_dff/N32 ), 
        .CLK(n1500), .Q(\i_m4stg_frac/ps[60] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[60]  ( .D(\i_m4stg_frac/n383 ), .CLK(
        n1500), .Q(\i_m4stg_frac/addin_sum[60] ), .QN(\i_m4stg_frac/n243 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[28]  ( .D(\i_m4stg_frac/psum_dff/N31 ), 
        .CLK(n1499), .Q(\i_m4stg_frac/ps[59] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[59]  ( .D(\i_m4stg_frac/n385 ), .CLK(
        n1499), .Q(\i_m4stg_frac/addin_sum[59] ), .QN(\i_m4stg_frac/n245 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[27]  ( .D(\i_m4stg_frac/psum_dff/N30 ), 
        .CLK(n1486), .Q(\i_m4stg_frac/ps[58] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[58]  ( .D(\i_m4stg_frac/n387 ), .CLK(
        n1485), .Q(\i_m4stg_frac/addin_sum[58] ), .QN(\i_m4stg_frac/n247 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[26]  ( .D(\i_m4stg_frac/psum_dff/N29 ), 
        .CLK(n1484), .Q(\i_m4stg_frac/ps[57] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[57]  ( .D(\i_m4stg_frac/n389 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_sum[57] ), .QN(\i_m4stg_frac/n249 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[25]  ( .D(\i_m4stg_frac/psum_dff/N28 ), 
        .CLK(n1484), .Q(\i_m4stg_frac/ps[56] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[56]  ( .D(\i_m4stg_frac/n391 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_sum[56] ), .QN(\i_m4stg_frac/n251 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[24]  ( .D(\i_m4stg_frac/psum_dff/N27 ), 
        .CLK(n1483), .Q(\i_m4stg_frac/ps[55] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[55]  ( .D(\i_m4stg_frac/n393 ), .CLK(
        n1485), .Q(\i_m4stg_frac/addin_sum[55] ), .QN(\i_m4stg_frac/n253 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[23]  ( .D(\i_m4stg_frac/psum_dff/N26 ), 
        .CLK(n1485), .Q(\i_m4stg_frac/ps[54] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[54]  ( .D(\i_m4stg_frac/n395 ), .CLK(
        n1485), .Q(\i_m4stg_frac/addin_sum[54] ), .QN(\i_m4stg_frac/n255 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[22]  ( .D(\i_m4stg_frac/psum_dff/N25 ), 
        .CLK(n1500), .Q(\i_m4stg_frac/ps[53] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[53]  ( .D(\i_m4stg_frac/n397 ), .CLK(
        n1500), .Q(\i_m4stg_frac/addin_sum[53] ), .QN(\i_m4stg_frac/n257 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[21]  ( .D(\i_m4stg_frac/psum_dff/N24 ), 
        .CLK(n1501), .Q(\i_m4stg_frac/ps[52] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[52]  ( .D(\i_m4stg_frac/n399 ), .CLK(
        n1501), .Q(\i_m4stg_frac/addin_sum[52] ), .QN(\i_m4stg_frac/n259 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[20]  ( .D(\i_m4stg_frac/psum_dff/N23 ), 
        .CLK(n1502), .Q(\i_m4stg_frac/ps[51] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[51]  ( .D(\i_m4stg_frac/n401 ), .CLK(
        n1502), .Q(\i_m4stg_frac/addin_sum[51] ), .QN(\i_m4stg_frac/n261 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[19]  ( .D(\i_m4stg_frac/psum_dff/N22 ), 
        .CLK(n1503), .Q(\i_m4stg_frac/ps[50] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[50]  ( .D(\i_m4stg_frac/n403 ), .CLK(
        n1503), .Q(\i_m4stg_frac/addin_sum[50] ), .QN(\i_m4stg_frac/n263 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[18]  ( .D(\i_m4stg_frac/psum_dff/N21 ), 
        .CLK(n1495), .Q(\i_m4stg_frac/ps[49] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[49]  ( .D(\i_m4stg_frac/n405 ), .CLK(
        n1496), .Q(\i_m4stg_frac/addin_sum[49] ), .QN(\i_m4stg_frac/n265 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[17]  ( .D(\i_m4stg_frac/psum_dff/N20 ), 
        .CLK(n1493), .Q(\i_m4stg_frac/ps[48] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[48]  ( .D(\i_m4stg_frac/n407 ), .CLK(
        n1493), .Q(\i_m4stg_frac/addin_sum[48] ), .QN(\i_m4stg_frac/n267 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[16]  ( .D(\i_m4stg_frac/psum_dff/N19 ), 
        .CLK(n1506), .Q(\i_m4stg_frac/ps[47] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[47]  ( .D(\i_m4stg_frac/n409 ), .CLK(
        n1506), .Q(\i_m4stg_frac/addin_sum[47] ), .QN(\i_m4stg_frac/n269 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[15]  ( .D(\i_m4stg_frac/psum_dff/N18 ), 
        .CLK(n1505), .Q(\i_m4stg_frac/ps[46] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[46]  ( .D(\i_m4stg_frac/n411 ), .CLK(
        n1506), .Q(\i_m4stg_frac/addin_sum[46] ), .QN(\i_m4stg_frac/n271 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[14]  ( .D(\i_m4stg_frac/psum_dff/N17 ), 
        .CLK(n1505), .Q(\i_m4stg_frac/ps[45] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[45]  ( .D(\i_m4stg_frac/n413 ), .CLK(
        n1505), .Q(\i_m4stg_frac/addin_sum[45] ), .QN(\i_m4stg_frac/n273 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[13]  ( .D(\i_m4stg_frac/psum_dff/N16 ), 
        .CLK(n1504), .Q(\i_m4stg_frac/ps[44] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[44]  ( .D(\i_m4stg_frac/n415 ), .CLK(
        n1504), .Q(\i_m4stg_frac/addin_sum[44] ), .QN(\i_m4stg_frac/n275 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[12]  ( .D(\i_m4stg_frac/psum_dff/N15 ), 
        .CLK(n1504), .Q(\i_m4stg_frac/ps[43] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[43]  ( .D(\i_m4stg_frac/n417 ), .CLK(
        n1504), .Q(\i_m4stg_frac/addin_sum[43] ), .QN(\i_m4stg_frac/n277 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[11]  ( .D(\i_m4stg_frac/psum_dff/N14 ), 
        .CLK(n1505), .Q(\i_m4stg_frac/ps[42] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[42]  ( .D(\i_m4stg_frac/n419 ), .CLK(
        n1505), .Q(\i_m4stg_frac/addin_sum[42] ), .QN(\i_m4stg_frac/n279 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[10]  ( .D(\i_m4stg_frac/psum_dff/N13 ), 
        .CLK(n1492), .Q(\i_m4stg_frac/ps[41] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[41]  ( .D(\i_m4stg_frac/n421 ), .CLK(
        n1492), .Q(\i_m4stg_frac/addin_sum[41] ), .QN(\i_m4stg_frac/n281 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[9]  ( .D(\i_m4stg_frac/psum_dff/N12 ), 
        .CLK(n1498), .Q(\i_m4stg_frac/ps[40] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[40]  ( .D(\i_m4stg_frac/n423 ), .CLK(
        n1498), .Q(\i_m4stg_frac/addin_sum[40] ), .QN(\i_m4stg_frac/n283 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[8]  ( .D(\i_m4stg_frac/psum_dff/N11 ), 
        .CLK(n1498), .Q(\i_m4stg_frac/ps[39] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[39]  ( .D(\i_m4stg_frac/n425 ), .CLK(
        n1498), .Q(\i_m4stg_frac/addin_sum[39] ), .QN(\i_m4stg_frac/n285 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[7]  ( .D(\i_m4stg_frac/psum_dff/N10 ), 
        .CLK(n1497), .Q(\i_m4stg_frac/ps[38] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[38]  ( .D(\i_m4stg_frac/n427 ), .CLK(
        n1497), .Q(\i_m4stg_frac/addin_sum[38] ), .QN(\i_m4stg_frac/n287 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[6]  ( .D(\i_m4stg_frac/psum_dff/N9 ), 
        .CLK(n1496), .Q(\i_m4stg_frac/ps[37] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[37]  ( .D(\i_m4stg_frac/n429 ), .CLK(
        n1496), .Q(\i_m4stg_frac/addin_sum[37] ), .QN(\i_m4stg_frac/n289 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[5]  ( .D(\i_m4stg_frac/psum_dff/N8 ), 
        .CLK(n1495), .Q(\i_m4stg_frac/ps[36] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[36]  ( .D(\i_m4stg_frac/n431 ), .CLK(
        n1495), .Q(\i_m4stg_frac/addin_sum[36] ), .QN(\i_m4stg_frac/n291 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[4]  ( .D(\i_m4stg_frac/psum_dff/N7 ), 
        .CLK(n1494), .Q(\i_m4stg_frac/ps[35] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[35]  ( .D(\i_m4stg_frac/n433 ), .CLK(
        n1494), .Q(\i_m4stg_frac/addin_sum[35] ), .QN(\i_m4stg_frac/n293 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[3]  ( .D(\i_m4stg_frac/psum_dff/N6 ), 
        .CLK(n1494), .Q(\i_m4stg_frac/ps[34] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[34]  ( .D(\i_m4stg_frac/n435 ), .CLK(
        n1494), .Q(\i_m4stg_frac/addin_sum[34] ), .QN(\i_m4stg_frac/n295 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[2]  ( .D(\i_m4stg_frac/psum_dff/N5 ), 
        .CLK(n1493), .Q(\i_m4stg_frac/ps[33] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[33]  ( .D(\i_m4stg_frac/n437 ), .CLK(
        n1493), .Q(\i_m4stg_frac/addin_sum[33] ), .QN(\i_m4stg_frac/n297 ) );
  DFFX1 \i_m4stg_frac/psum_dff/q_reg[1]  ( .D(\i_m4stg_frac/psum_dff/N4 ), 
        .CLK(n1499), .Q(\i_m4stg_frac/ps[32] ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[32]  ( .D(\i_m4stg_frac/n439 ), .CLK(
        n1499), .Q(\i_m4stg_frac/addin_sum[32] ), .QN(\i_m4stg_frac/n299 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[31]  ( .D(\i_m4stg_frac/n453 ), .CLK(
        n1502), .Q(\i_m4stg_frac/addin_sum[31] ), .QN(\i_m4stg_frac/n301 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[30]  ( .D(\i_m4stg_frac/n455 ), .CLK(
        n1485), .Q(\i_m4stg_frac/addin_sum[30] ), .QN(\i_m4stg_frac/n302 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[29]  ( .D(\i_m4stg_frac/n457 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_sum[29] ), .QN(\i_m4stg_frac/n303 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[28]  ( .D(\i_m4stg_frac/n459 ), .CLK(
        n1483), .Q(\i_m4stg_frac/addin_sum[28] ), .QN(\i_m4stg_frac/n304 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[27]  ( .D(\i_m4stg_frac/n461 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_sum[27] ), .QN(\i_m4stg_frac/n305 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[26]  ( .D(\i_m4stg_frac/n463 ), .CLK(
        n1483), .Q(\i_m4stg_frac/addin_sum[26] ), .QN(\i_m4stg_frac/n306 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[25]  ( .D(\i_m4stg_frac/n465 ), .CLK(
        n1483), .Q(\i_m4stg_frac/addin_sum[25] ), .QN(\i_m4stg_frac/n307 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[24]  ( .D(\i_m4stg_frac/n467 ), .CLK(
        n1483), .Q(\i_m4stg_frac/addin_sum[24] ), .QN(\i_m4stg_frac/n308 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[23]  ( .D(\i_m4stg_frac/n469 ), .CLK(
        n1484), .Q(\i_m4stg_frac/addin_sum[23] ), .QN(\i_m4stg_frac/n309 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[22]  ( .D(\i_m4stg_frac/n471 ), .CLK(
        n1485), .Q(\i_m4stg_frac/addin_sum[22] ), .QN(\i_m4stg_frac/n310 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[21]  ( .D(\i_m4stg_frac/n609 ), .CLK(
        n1500), .Q(\i_m4stg_frac/addin_sum[21] ), .QN(\i_m4stg_frac/n311 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[20]  ( .D(\i_m4stg_frac/n492 ), .CLK(
        n1501), .Q(\i_m4stg_frac/addin_sum[20] ), .QN(\i_m4stg_frac/n312 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[19]  ( .D(\i_m4stg_frac/n473 ), .CLK(
        n1502), .Q(\i_m4stg_frac/addin_sum[19] ), .QN(\i_m4stg_frac/n313 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[18]  ( .D(\i_m4stg_frac/n475 ), .CLK(
        n1503), .Q(\i_m4stg_frac/addin_sum[18] ), .QN(\i_m4stg_frac/n314 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[17]  ( .D(\i_m4stg_frac/n477 ), .CLK(
        n1505), .Q(\i_m4stg_frac/addin_sum[17] ), .QN(\i_m4stg_frac/n315 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[16]  ( .D(\i_m4stg_frac/n479 ), .CLK(
        n1504), .Q(\i_m4stg_frac/addin_sum[16] ), .QN(\i_m4stg_frac/n316 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[15]  ( .D(\i_m4stg_frac/n611 ), .CLK(
        n1504), .Q(\i_m4stg_frac/addin_sum[15] ), .QN(\i_m4stg_frac/n317 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[14]  ( .D(\i_m4stg_frac/n447 ), .CLK(
        n1503), .Q(\i_m4stg_frac/addin_sum[14] ), .QN(\i_m4stg_frac/n318 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[13]  ( .D(\i_m4stg_frac/n481 ), .CLK(
        n1503), .Q(\i_m4stg_frac/addin_sum[13] ), .QN(\i_m4stg_frac/n319 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[12]  ( .D(\i_m4stg_frac/n483 ), .CLK(
        n1503), .Q(\i_m4stg_frac/addin_sum[12] ), .QN(\i_m4stg_frac/n320 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[11]  ( .D(\i_m4stg_frac/n485 ), .CLK(
        n1504), .Q(\i_m4stg_frac/addin_sum[11] ), .QN(\i_m4stg_frac/n321 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[10]  ( .D(\i_m4stg_frac/n449 ), .CLK(
        n1505), .Q(\i_m4stg_frac/addin_sum[10] ), .QN(\i_m4stg_frac/n322 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[9]  ( .D(\i_m4stg_frac/n451 ), .CLK(
        n1491), .Q(\i_m4stg_frac/addin_sum[9] ), .QN(\i_m4stg_frac/n323 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[8]  ( .D(\i_m4stg_frac/n487 ), .CLK(
        n1497), .Q(\i_m4stg_frac/addin_sum[8] ), .QN(\i_m4stg_frac/n324 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[7]  ( .D(\i_m4stg_frac/n489 ), .CLK(
        n1498), .Q(\i_m4stg_frac/addin_sum[7] ), .QN(\i_m4stg_frac/n325 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[6]  ( .D(\i_m4stg_frac/n491 ), .CLK(
        n1497), .Q(\i_m4stg_frac/addin_sum[6] ), .QN(\i_m4stg_frac/n326 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[5]  ( .D(\i_m4stg_frac/n631 ), .CLK(
        n1496), .Q(\i_m4stg_frac/addin_sum[5] ), .QN(\i_m4stg_frac/n327 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[4]  ( .D(\i_m4stg_frac/n633 ), .CLK(
        n1495), .Q(\i_m4stg_frac/addin_sum[4] ), .QN(\i_m4stg_frac/n328 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[3]  ( .D(\i_m4stg_frac/n613 ), .CLK(
        n1499), .Q(\i_m4stg_frac/addin_sum[3] ), .QN(\i_m4stg_frac/n329 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[2]  ( .D(\i_m4stg_frac/n615 ), .CLK(
        n1486), .Q(n1165) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[1]  ( .D(\i_m4stg_frac/n617 ), .CLK(
        n1486), .Q(\i_m4stg_frac/addin_sum[1] ), .QN(\i_m4stg_frac/n331 ) );
  DFFX1 \i_m4stg_frac/a2sum_dff/q_reg[0]  ( .D(\i_m4stg_frac/n619 ), .CLK(
        n1486), .Q(\i_m4stg_frac/addin_sum[0] ), .QN(\i_m4stg_frac/n332 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[75]  ( .D(\i_m4stg_frac/a1cout[79] ), 
        .RSTB(n1525), .SETB(1'b1), .CLK(n1460), .Q(\i_m4stg_frac/a1c[79] ), 
        .QN(\i_m4stg_frac/n338 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[74]  ( .D(\i_m4stg_frac/a1cout[78] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1462), .Q(\i_m4stg_frac/a1c[78] ), 
        .QN(\i_m4stg_frac/n340 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[73]  ( .D(\i_m4stg_frac/a1cout[77] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1462), .Q(\i_m4stg_frac/a1c[77] ), 
        .QN(\i_m4stg_frac/n342 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[72]  ( .D(\i_m4stg_frac/a1cout[76] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1c[76] ), 
        .QN(\i_m4stg_frac/n344 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[71]  ( .D(\i_m4stg_frac/a1cout[75] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1c[75] ), 
        .QN(\i_m4stg_frac/n346 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[70]  ( .D(\i_m4stg_frac/a1cout[74] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1c[74] ), 
        .QN(\i_m4stg_frac/n348 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[69]  ( .D(\i_m4stg_frac/a1cout[73] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1c[73] ), 
        .QN(\i_m4stg_frac/n350 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[68]  ( .D(\i_m4stg_frac/a1cout[72] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1c[72] ), 
        .QN(\i_m4stg_frac/n352 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[67]  ( .D(\i_m4stg_frac/a1cout[71] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1c[71] ), 
        .QN(\i_m4stg_frac/n354 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[66]  ( .D(\i_m4stg_frac/a1cout[70] ), 
        .RSTB(n1534), .SETB(1'b1), .CLK(n1482), .Q(\i_m4stg_frac/a1c[70] ), 
        .QN(\i_m4stg_frac/n356 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[65]  ( .D(\i_m4stg_frac/a1cout[69] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1480), .Q(\i_m4stg_frac/a1c[69] ), 
        .QN(\i_m4stg_frac/n358 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[64]  ( .D(\i_m4stg_frac/a1cout[68] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1481), .Q(\i_m4stg_frac/a1c[68] ), 
        .QN(\i_m4stg_frac/n360 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[63]  ( .D(\i_m4stg_frac/a1cout[67] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1480), .Q(\i_m4stg_frac/a1c[67] ), 
        .QN(\i_m4stg_frac/n362 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[62]  ( .D(\i_m4stg_frac/a1cout[66] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1473), .Q(\i_m4stg_frac/a1c[66] ), 
        .QN(\i_m4stg_frac/n364 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[61]  ( .D(\i_m4stg_frac/a1cout[65] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1c[65] ), 
        .QN(\i_m4stg_frac/n366 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[60]  ( .D(\i_m4stg_frac/a1cout[64] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1c[64] ), 
        .QN(\i_m4stg_frac/n368 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[59]  ( .D(\i_m4stg_frac/a1cout[63] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1c[63] ), 
        .QN(\i_m4stg_frac/n370 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[58]  ( .D(\i_m4stg_frac/a1cout[62] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1c[62] ), 
        .QN(\i_m4stg_frac/n372 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[57]  ( .D(\i_m4stg_frac/a1cout[61] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1c[61] ), 
        .QN(\i_m4stg_frac/n374 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[56]  ( .D(\i_m4stg_frac/a1cout[60] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1c[60] ), 
        .QN(\i_m4stg_frac/n376 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[55]  ( .D(\i_m4stg_frac/a1cout[59] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1450), .Q(\i_m4stg_frac/a1c[59] ), 
        .QN(\i_m4stg_frac/n378 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[54]  ( .D(\i_m4stg_frac/a1cout[58] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1452), .Q(\i_m4stg_frac/a1c[58] ), 
        .QN(\i_m4stg_frac/n380 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[53]  ( .D(\i_m4stg_frac/a1cout[57] ), 
        .RSTB(\i_m4stg_frac/n854 ), .SETB(1'b1), .CLK(n1481), .Q(
        \i_m4stg_frac/a1c[57] ), .QN(\i_m4stg_frac/n382 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[52]  ( .D(\i_m4stg_frac/a1cout[56] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1460), .Q(\i_m4stg_frac/a1c[56] ), 
        .QN(\i_m4stg_frac/n384 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[51]  ( .D(\i_m4stg_frac/a1cout[55] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1460), .Q(\i_m4stg_frac/a1c[55] ), 
        .QN(\i_m4stg_frac/n386 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[50]  ( .D(\i_m4stg_frac/a1cout[54] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1459), .Q(\i_m4stg_frac/a1c[54] ), 
        .QN(\i_m4stg_frac/n388 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[49]  ( .D(\i_m4stg_frac/a1cout[53] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1459), .Q(\i_m4stg_frac/a1c[53] ), 
        .QN(\i_m4stg_frac/n390 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[48]  ( .D(\i_m4stg_frac/a1cout[52] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1459), .Q(\i_m4stg_frac/a1c[52] ), 
        .QN(\i_m4stg_frac/n392 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[47]  ( .D(\i_m4stg_frac/a1cout[51] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1459), .Q(\i_m4stg_frac/a1c[51] ), 
        .QN(\i_m4stg_frac/n394 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[46]  ( .D(\i_m4stg_frac/a1cout[50] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1459), .Q(\i_m4stg_frac/a1c[50] ), 
        .QN(\i_m4stg_frac/n396 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[45]  ( .D(\i_m4stg_frac/a1cout[49] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1458), .Q(\i_m4stg_frac/a1c[49] ), 
        .QN(\i_m4stg_frac/n398 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[44]  ( .D(\i_m4stg_frac/a1cout[48] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1458), .Q(\i_m4stg_frac/a1c[48] ), 
        .QN(\i_m4stg_frac/n400 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[43]  ( .D(\i_m4stg_frac/a1cout[47] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1458), .Q(\i_m4stg_frac/a1c[47] ), 
        .QN(\i_m4stg_frac/n402 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[42]  ( .D(\i_m4stg_frac/a1cout[46] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1458), .Q(\i_m4stg_frac/a1c[46] ), 
        .QN(\i_m4stg_frac/n404 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[41]  ( .D(\i_m4stg_frac/a1cout[45] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1458), .Q(\i_m4stg_frac/a1c[45] ), 
        .QN(\i_m4stg_frac/n406 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[40]  ( .D(\i_m4stg_frac/a1cout[44] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1458), .Q(\i_m4stg_frac/a1c[44] ), 
        .QN(\i_m4stg_frac/n408 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[39]  ( .D(\i_m4stg_frac/a1cout[43] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1457), .Q(\i_m4stg_frac/a1c[43] ), 
        .QN(\i_m4stg_frac/n410 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[38]  ( .D(\i_m4stg_frac/a1cout[42] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1457), .Q(\i_m4stg_frac/a1c[42] ), 
        .QN(\i_m4stg_frac/n412 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[37]  ( .D(\i_m4stg_frac/a1cout[41] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1457), .Q(\i_m4stg_frac/a1c[41] ), 
        .QN(\i_m4stg_frac/n414 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[36]  ( .D(\i_m4stg_frac/a1cout[40] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1457), .Q(\i_m4stg_frac/a1c[40] ), 
        .QN(\i_m4stg_frac/n416 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[35]  ( .D(\i_m4stg_frac/a1cout[39] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1457), .Q(\i_m4stg_frac/a1c[39] ), 
        .QN(\i_m4stg_frac/n418 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[34]  ( .D(\i_m4stg_frac/a1cout[38] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1457), .Q(\i_m4stg_frac/a1c[38] ), 
        .QN(\i_m4stg_frac/n420 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[33]  ( .D(\i_m4stg_frac/a1cout[37] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1456), .Q(\i_m4stg_frac/a1c[37] ), 
        .QN(\i_m4stg_frac/n422 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[32]  ( .D(\i_m4stg_frac/a1cout[36] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1456), .Q(\i_m4stg_frac/a1c[36] ), 
        .QN(\i_m4stg_frac/n424 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[31]  ( .D(\i_m4stg_frac/a1cout[35] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1456), .Q(\i_m4stg_frac/a1c[35] ), 
        .QN(\i_m4stg_frac/n426 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[30]  ( .D(\i_m4stg_frac/a1cout[34] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1456), .Q(\i_m4stg_frac/a1c[34] ), 
        .QN(\i_m4stg_frac/n428 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[29]  ( .D(\i_m4stg_frac/a1cout[33] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1456), .Q(\i_m4stg_frac/a1c[33] ), 
        .QN(\i_m4stg_frac/n430 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[28]  ( .D(\i_m4stg_frac/a1cout[32] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1456), .Q(\i_m4stg_frac/a1c[32] ), 
        .QN(\i_m4stg_frac/n432 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[27]  ( .D(\i_m4stg_frac/a1cout[31] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1455), .Q(\i_m4stg_frac/a1c[31] ), 
        .QN(\i_m4stg_frac/n434 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[26]  ( .D(\i_m4stg_frac/a1cout[30] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1455), .Q(\i_m4stg_frac/a1c[30] ), 
        .QN(\i_m4stg_frac/n436 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[25]  ( .D(\i_m4stg_frac/a1cout[29] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1455), .Q(\i_m4stg_frac/a1c[29] ), 
        .QN(\i_m4stg_frac/n438 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[24]  ( .D(\i_m4stg_frac/a1cout[28] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1455), .Q(\i_m4stg_frac/a1c[28] ), 
        .QN(\i_m4stg_frac/n440 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[23]  ( .D(\i_m4stg_frac/a1cout[27] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1455), .Q(\i_m4stg_frac/a1c[27] ), 
        .QN(\i_m4stg_frac/n442 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[22]  ( .D(\i_m4stg_frac/a1cout[26] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1455), .Q(\i_m4stg_frac/a1c[26] ), 
        .QN(\i_m4stg_frac/n444 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[21]  ( .D(\i_m4stg_frac/a1cout[25] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1454), .Q(\i_m4stg_frac/a1c[25] ), 
        .QN(\i_m4stg_frac/n446 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[20]  ( .D(\i_m4stg_frac/a1cout[24] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1454), .Q(\i_m4stg_frac/a1c[24] ), 
        .QN(\i_m4stg_frac/n448 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[19]  ( .D(\i_m4stg_frac/a1cout[23] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1454), .Q(\i_m4stg_frac/a1c[23] ), 
        .QN(\i_m4stg_frac/n450 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[18]  ( .D(\i_m4stg_frac/a1cout[22] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1454), .Q(\i_m4stg_frac/a1c[22] ), 
        .QN(\i_m4stg_frac/n452 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[17]  ( .D(\i_m4stg_frac/a1cout[21] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1454), .Q(\i_m4stg_frac/a1c[21] ), 
        .QN(\i_m4stg_frac/n454 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[16]  ( .D(\i_m4stg_frac/a1cout[20] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1453), .Q(\i_m4stg_frac/a1c[20] ), 
        .QN(\i_m4stg_frac/n456 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[15]  ( .D(\i_m4stg_frac/a1cout[19] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1453), .Q(\i_m4stg_frac/a1c[19] ), 
        .QN(\i_m4stg_frac/n458 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[14]  ( .D(\i_m4stg_frac/a1cout[18] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1453), .Q(\i_m4stg_frac/a1c[18] ), 
        .QN(\i_m4stg_frac/n460 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[13]  ( .D(\i_m4stg_frac/a1cout[17] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1453), .Q(\i_m4stg_frac/a1c[17] ), 
        .QN(\i_m4stg_frac/n462 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[12]  ( .D(\i_m4stg_frac/a1cout[16] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1453), .Q(\i_m4stg_frac/a1c[16] ), 
        .QN(\i_m4stg_frac/n464 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[11]  ( .D(\i_m4stg_frac/a1cout[15] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1453), .Q(\i_m4stg_frac/a1c[15] ), 
        .QN(\i_m4stg_frac/n466 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[10]  ( .D(\i_m4stg_frac/a1cout[14] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1452), .Q(\i_m4stg_frac/a1c[14] ), 
        .QN(\i_m4stg_frac/n468 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[9]  ( .D(\i_m4stg_frac/a1cout[13] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1452), .Q(\i_m4stg_frac/a1c[13] ), 
        .QN(\i_m4stg_frac/n470 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[8]  ( .D(\i_m4stg_frac/a1cout[12] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1452), .Q(\i_m4stg_frac/a1c[12] ), 
        .QN(\i_m4stg_frac/n472 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[7]  ( .D(\i_m4stg_frac/a1cout[11] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1452), .Q(\i_m4stg_frac/a1c[11] ), 
        .QN(\i_m4stg_frac/n474 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[6]  ( .D(\i_m4stg_frac/a1cout[10] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1452), .Q(\i_m4stg_frac/a1c[10] ), 
        .QN(\i_m4stg_frac/n476 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[5]  ( .D(\i_m4stg_frac/a1cout[9] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1477), .Q(\i_m4stg_frac/a1c[9] ), 
        .QN(\i_m4stg_frac/n478 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[4]  ( .D(\i_m4stg_frac/a1cout[8] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1472), .Q(\i_m4stg_frac/a1c[8] ), 
        .QN(\i_m4stg_frac/n480 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[3]  ( .D(\i_m4stg_frac/a1cout[7] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1472), .Q(\i_m4stg_frac/a1c[7] ), 
        .QN(\i_m4stg_frac/n482 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[2]  ( .D(\i_m4stg_frac/a1cout[6] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1473), .Q(\i_m4stg_frac/a1c[6] ), 
        .QN(\i_m4stg_frac/n484 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[1]  ( .D(\i_m4stg_frac/a1cout[5] ), 
        .RSTB(\i_m4stg_frac/n854 ), .SETB(1'b1), .CLK(n1474), .Q(
        \i_m4stg_frac/a1c[5] ), .QN(\i_m4stg_frac/n486 ) );
  DFFSSRX1 \i_m4stg_frac/a1cot_dff/q_reg[0]  ( .D(\i_m4stg_frac/a1cout[4] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1459), .Q(\i_m4stg_frac/a1c[4] ), 
        .QN(\i_m4stg_frac/n488 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[81]  ( .D(\i_m4stg_frac/a1sum[81] ), 
        .RSTB(n1522), .SETB(1'b1), .CLK(n1466), .Q(n1339), .QN(
        \i_m4stg_frac/n490 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[79]  ( .D(\i_m4stg_frac/a1sum[79] ), 
        .RSTB(n1525), .SETB(1'b1), .CLK(n1460), .Q(\i_m4stg_frac/a1s[79] ), 
        .QN(\i_m4stg_frac/n494 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[78]  ( .D(\i_m4stg_frac/a1sum[78] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1462), .Q(\i_m4stg_frac/a1s[78] ), 
        .QN(\i_m4stg_frac/n496 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[77]  ( .D(\i_m4stg_frac/a1sum[77] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1462), .Q(\i_m4stg_frac/a1s[77] ), 
        .QN(\i_m4stg_frac/n498 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[76]  ( .D(\i_m4stg_frac/a1sum[76] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1462), .Q(\i_m4stg_frac/a1s[76] ), 
        .QN(\i_m4stg_frac/n500 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[75]  ( .D(\i_m4stg_frac/a1sum[75] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1s[75] ), 
        .QN(\i_m4stg_frac/n502 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[74]  ( .D(\i_m4stg_frac/a1sum[74] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1s[74] ), 
        .QN(\i_m4stg_frac/n504 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[73]  ( .D(\i_m4stg_frac/a1sum[73] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1s[73] ), 
        .QN(\i_m4stg_frac/n506 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[72]  ( .D(\i_m4stg_frac/a1sum[72] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1s[72] ), 
        .QN(\i_m4stg_frac/n508 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[71]  ( .D(\i_m4stg_frac/a1sum[71] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1461), .Q(\i_m4stg_frac/a1s[71] ), 
        .QN(\i_m4stg_frac/n510 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[70]  ( .D(\i_m4stg_frac/a1sum[70] ), 
        .RSTB(n1534), .SETB(1'b1), .CLK(n1483), .Q(\i_m4stg_frac/a1s[70] ), 
        .QN(\i_m4stg_frac/n512 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[69]  ( .D(\i_m4stg_frac/a1sum[69] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1480), .Q(\i_m4stg_frac/a1s[69] ), 
        .QN(\i_m4stg_frac/n514 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[68]  ( .D(\i_m4stg_frac/a1sum[68] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1480), .Q(\i_m4stg_frac/a1s[68] ), 
        .QN(\i_m4stg_frac/n516 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[67]  ( .D(\i_m4stg_frac/a1sum[67] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1477), .Q(\i_m4stg_frac/a1s[67] ), 
        .QN(\i_m4stg_frac/n518 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[66]  ( .D(\i_m4stg_frac/a1sum[66] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1473), .Q(\i_m4stg_frac/a1s[66] ), 
        .QN(\i_m4stg_frac/n520 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[65]  ( .D(\i_m4stg_frac/a1sum[65] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1s[65] ), 
        .QN(\i_m4stg_frac/n522 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[64]  ( .D(\i_m4stg_frac/a1sum[64] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1s[64] ), 
        .QN(\i_m4stg_frac/n524 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[63]  ( .D(\i_m4stg_frac/a1sum[63] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1s[63] ), 
        .QN(\i_m4stg_frac/n526 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[62]  ( .D(\i_m4stg_frac/a1sum[62] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1s[62] ), 
        .QN(\i_m4stg_frac/n528 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[61]  ( .D(\i_m4stg_frac/a1sum[61] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1s[61] ), 
        .QN(\i_m4stg_frac/n530 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[60]  ( .D(\i_m4stg_frac/a1sum[60] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1451), .Q(\i_m4stg_frac/a1s[60] ), 
        .QN(\i_m4stg_frac/n532 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[59]  ( .D(\i_m4stg_frac/a1sum[59] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1450), .Q(\i_m4stg_frac/a1s[59] ), 
        .QN(\i_m4stg_frac/n534 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[58]  ( .D(\i_m4stg_frac/a1sum[58] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1452), .Q(\i_m4stg_frac/a1s[58] ), 
        .QN(\i_m4stg_frac/n536 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[57]  ( .D(\i_m4stg_frac/a1sum[57] ), 
        .RSTB(\i_m4stg_frac/n854 ), .SETB(1'b1), .CLK(n1480), .Q(
        \i_m4stg_frac/a1s[57] ), .QN(\i_m4stg_frac/n538 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[56]  ( .D(\i_m4stg_frac/a1sum[56] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1460), .Q(\i_m4stg_frac/a1s[56] ), 
        .QN(\i_m4stg_frac/n540 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[55]  ( .D(\i_m4stg_frac/a1sum[55] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1460), .Q(\i_m4stg_frac/a1s[55] ), 
        .QN(\i_m4stg_frac/n542 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[54]  ( .D(\i_m4stg_frac/a1sum[54] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1459), .Q(\i_m4stg_frac/a1s[54] ), 
        .QN(\i_m4stg_frac/n544 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[53]  ( .D(\i_m4stg_frac/a1sum[53] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1459), .Q(\i_m4stg_frac/a1s[53] ), 
        .QN(\i_m4stg_frac/n546 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[52]  ( .D(\i_m4stg_frac/a1sum[52] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1459), .Q(\i_m4stg_frac/a1s[52] ), 
        .QN(\i_m4stg_frac/n548 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[51]  ( .D(\i_m4stg_frac/a1sum[51] ), 
        .RSTB(n1552), .SETB(1'b1), .CLK(n1459), .Q(\i_m4stg_frac/a1s[51] ), 
        .QN(\i_m4stg_frac/n550 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[50]  ( .D(\i_m4stg_frac/a1sum[50] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1459), .Q(n1111) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[49]  ( .D(\i_m4stg_frac/a1sum[49] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1458), .Q(n1110) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[48]  ( .D(\i_m4stg_frac/a1sum[48] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1458), .Q(n1109) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[47]  ( .D(\i_m4stg_frac/a1sum[47] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1458), .Q(n1108) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[46]  ( .D(\i_m4stg_frac/a1sum[46] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1458), .Q(n1107) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[45]  ( .D(\i_m4stg_frac/a1sum[45] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1458), .Q(n1106) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[44]  ( .D(\i_m4stg_frac/a1sum[44] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1457), .Q(n1105) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[43]  ( .D(\i_m4stg_frac/a1sum[43] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1457), .Q(n1104) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[42]  ( .D(\i_m4stg_frac/a1sum[42] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1457), .Q(n1103) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[41]  ( .D(\i_m4stg_frac/a1sum[41] ), 
        .RSTB(n1550), .SETB(1'b1), .CLK(n1457), .Q(n1102) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[40]  ( .D(\i_m4stg_frac/a1sum[40] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1457), .Q(n1101) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[39]  ( .D(\i_m4stg_frac/a1sum[39] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1457), .Q(n1100) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[38]  ( .D(\i_m4stg_frac/a1sum[38] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1456), .Q(n1099) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[37]  ( .D(\i_m4stg_frac/a1sum[37] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1456), .Q(n1098) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[36]  ( .D(\i_m4stg_frac/a1sum[36] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1456), .Q(n1097) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[35]  ( .D(\i_m4stg_frac/a1sum[35] ), 
        .RSTB(n1549), .SETB(1'b1), .CLK(n1456), .Q(n1096) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[34]  ( .D(\i_m4stg_frac/a1sum[34] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1456), .Q(n1095) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[33]  ( .D(\i_m4stg_frac/a1sum[33] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1456), .Q(n1094) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[32]  ( .D(\i_m4stg_frac/a1sum[32] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1455), .Q(n1093) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[31]  ( .D(\i_m4stg_frac/a1sum[31] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1455), .Q(n1092) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[30]  ( .D(\i_m4stg_frac/a1sum[30] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1455), .Q(n1091) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[29]  ( .D(\i_m4stg_frac/a1sum[29] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1455), .Q(n1090) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[28]  ( .D(\i_m4stg_frac/a1sum[28] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1455), .Q(n1089) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[27]  ( .D(\i_m4stg_frac/a1sum[27] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1455), .Q(n1088) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[26]  ( .D(\i_m4stg_frac/a1sum[26] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1454), .Q(n1087) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[25]  ( .D(\i_m4stg_frac/a1sum[25] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1454), .Q(n1086) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[24]  ( .D(\i_m4stg_frac/a1sum[24] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1454), .Q(n1085) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[23]  ( .D(\i_m4stg_frac/a1sum[23] ), 
        .RSTB(n1547), .SETB(1'b1), .CLK(n1454), .Q(n1084) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[22]  ( .D(\i_m4stg_frac/a1sum[22] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1454), .Q(n1083) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[21]  ( .D(\i_m4stg_frac/a1sum[21] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1454), .Q(n1082) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[20]  ( .D(\i_m4stg_frac/a1sum[20] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1453), .Q(n1081) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[19]  ( .D(\i_m4stg_frac/a1sum[19] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1453), .Q(n1080) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[18]  ( .D(\i_m4stg_frac/a1sum[18] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1453), .Q(n1079) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[17]  ( .D(\i_m4stg_frac/a1sum[17] ), 
        .RSTB(n1546), .SETB(1'b1), .CLK(n1453), .Q(n1078) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[16]  ( .D(\i_m4stg_frac/a1sum[16] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1453), .Q(n1077) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[15]  ( .D(\i_m4stg_frac/a1sum[15] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1453), .Q(n1076) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[14]  ( .D(\i_m4stg_frac/a1sum[14] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1452), .Q(n1075) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[13]  ( .D(\i_m4stg_frac/a1sum[13] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1452), .Q(n1074) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[12]  ( .D(\i_m4stg_frac/a1sum[12] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1452), .Q(n1067) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[11]  ( .D(\i_m4stg_frac/a1sum[11] ), 
        .RSTB(n1545), .SETB(1'b1), .CLK(n1452), .Q(n1066) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[10]  ( .D(\i_m4stg_frac/a1sum[10] ), 
        .RSTB(n1544), .SETB(1'b1), .CLK(n1452), .Q(n1065) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[9]  ( .D(\i_m4stg_frac/a1sum[9] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1477), .Q(n1064) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[8]  ( .D(\i_m4stg_frac/a1sum[8] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1479), .Q(n1063) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[7]  ( .D(\i_m4stg_frac/a1sum[7] ), 
        .RSTB(n1533), .SETB(1'b1), .CLK(n1472), .Q(n1062) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[6]  ( .D(\i_m4stg_frac/a1sum[6] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1472), .Q(n1061) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[5]  ( .D(\i_m4stg_frac/a1sum[5] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1473), .Q(n1191), .QN(
        \i_m4stg_frac/n642 ) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[4]  ( .D(\i_m4stg_frac/a1sum[4] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1459), .Q(n1126) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[3]  ( .D(\i_m4stg_frac/a1sum[3] ), 
        .RSTB(n1551), .SETB(1'b1), .CLK(n1458), .Q(n1130) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[2]  ( .D(\i_m4stg_frac/a1sum[2] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1450), .Q(n1128) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[1]  ( .D(\i_m4stg_frac/a1sum[1] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1450), .Q(n1129) );
  DFFSSRX1 \i_m4stg_frac/a1sum_dff/q_reg[0]  ( .D(\i_m4stg_frac/a1sum[0] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1450), .Q(n1199), .QN(
        \i_m4stg_frac/n652 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff15/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff15/N5 ), .CLK(n1491), .Q(
        \i_m4stg_frac/b15[2] ), .QN(\i_m4stg_frac/n654 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff15/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff15/N4 ), .CLK(n1490), .Q(n938), .QN(
        \i_m4stg_frac/n655 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff15/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff15/N3 ), .CLK(n1491), .Q(n1123), .QN(
        \i_m4stg_frac/n656 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff14/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff14/N5 ), .CLK(n1491), .Q(n1039), .QN(
        \i_m4stg_frac/n657 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff14/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff14/N4 ), .CLK(n1489), .Q(n1133), .QN(
        \i_m4stg_frac/n658 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff14/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff14/N3 ), .CLK(n1489), .Q(n1313), .QN(
        \i_m4stg_frac/n659 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff13/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff13/N5 ), .CLK(n1489), .Q(n934), .QN(
        \i_m4stg_frac/n660 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff13/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff13/N4 ), .CLK(n1489), .Q(n1143) );
  DFFX1 \i_m4stg_frac/booth/out_dff13/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff13/N3 ), .CLK(n1489), .Q(n949), .QN(
        \i_m4stg_frac/n662 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff12/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff12/N5 ), .CLK(n1489), .Q(
        \i_m4stg_frac/b12[2] ), .QN(\i_m4stg_frac/n663 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff12/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff12/N4 ), .CLK(n1489), .Q(n1116), .QN(
        \i_m4stg_frac/n664 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff12/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff12/N3 ), .CLK(n1489), .Q(n914), .QN(
        \i_m4stg_frac/n665 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff11/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff11/N5 ), .CLK(n1489), .Q(n912), .QN(
        \i_m4stg_frac/n666 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff11/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff11/N4 ), .CLK(n1489), .Q(n1168), .QN(
        \i_m4stg_frac/n667 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff11/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff11/N3 ), .CLK(n1489), .Q(
        \i_m4stg_frac/b11[0] ), .QN(\i_m4stg_frac/n668 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff10/q_reg[2]  ( .D(\i_m4stg_frac/n1283 ), 
        .CLK(n1490), .Q(n937), .QN(\i_m4stg_frac/n669 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff10/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff10/N4 ), .CLK(n1490), .Q(n1142) );
  DFFX1 \i_m4stg_frac/booth/out_dff10/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff10/N3 ), .CLK(n1490), .Q(n948), .QN(
        \i_m4stg_frac/n671 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff9/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff9/N5 ), .CLK(n1490), .Q(
        \i_m4stg_frac/b9[2] ), .QN(\i_m4stg_frac/n672 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff9/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff9/N4 ), .CLK(n1501), .Q(n1117), .QN(
        \i_m4stg_frac/n673 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff9/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff9/N3 ), .CLK(n1501), .Q(n924), .QN(
        \i_m4stg_frac/n674 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff8/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff8/N5 ), .CLK(n1500), .Q(n1040), .QN(
        \i_m4stg_frac/n675 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff8/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff8/N4 ), .CLK(n1500), .Q(n1134), .QN(
        \i_m4stg_frac/n676 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff8/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff8/N3 ), .CLK(n1500), .Q(
        \i_m4stg_frac/b8[0] ), .QN(\i_m4stg_frac/n677 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[75]  ( .D(\i_m4stg_frac/a0cout[79] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1450), .Q(\i_m4stg_frac/a0c[79] ), 
        .QN(\i_m4stg_frac/n683 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[74]  ( .D(\i_m4stg_frac/a0cout[78] ), 
        .RSTB(n1548), .SETB(1'b1), .CLK(n1450), .Q(\i_m4stg_frac/a0c[78] ), 
        .QN(\i_m4stg_frac/n685 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[73]  ( .D(\i_m4stg_frac/a0cout[77] ), 
        .RSTB(n1522), .SETB(1'b1), .CLK(n1450), .Q(\i_m4stg_frac/a0c[77] ), 
        .QN(\i_m4stg_frac/n687 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[72]  ( .D(\i_m4stg_frac/a0cout[76] ), 
        .RSTB(n1522), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0c[76] ), 
        .QN(\i_m4stg_frac/n689 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[71]  ( .D(\i_m4stg_frac/a0cout[75] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0c[75] ), 
        .QN(\i_m4stg_frac/n691 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[70]  ( .D(\i_m4stg_frac/a0cout[74] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0c[74] ), 
        .QN(\i_m4stg_frac/n693 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[69]  ( .D(\i_m4stg_frac/a0cout[73] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0c[73] ), 
        .QN(\i_m4stg_frac/n695 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[68]  ( .D(\i_m4stg_frac/a0cout[72] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0c[72] ), 
        .QN(\i_m4stg_frac/n697 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[67]  ( .D(\i_m4stg_frac/a0cout[71] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0c[71] ), 
        .QN(\i_m4stg_frac/n699 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[66]  ( .D(\i_m4stg_frac/a0cout[70] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0c[70] ), 
        .QN(\i_m4stg_frac/n701 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[65]  ( .D(\i_m4stg_frac/a0cout[69] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1448), .Q(\i_m4stg_frac/a0c[69] ), 
        .QN(\i_m4stg_frac/n703 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[64]  ( .D(\i_m4stg_frac/a0cout[68] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1448), .Q(\i_m4stg_frac/a0c[68] ), 
        .QN(\i_m4stg_frac/n705 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[63]  ( .D(\i_m4stg_frac/a0cout[67] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1448), .Q(\i_m4stg_frac/a0c[67] ), 
        .QN(\i_m4stg_frac/n707 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[62]  ( .D(\i_m4stg_frac/a0cout[66] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1448), .Q(n928) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[61]  ( .D(\i_m4stg_frac/a0cout[65] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1448), .Q(\i_m4stg_frac/a0c[65] ), 
        .QN(\i_m4stg_frac/n711 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[60]  ( .D(\i_m4stg_frac/a0cout[64] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1472), .Q(\i_m4stg_frac/a0c[64] ), 
        .QN(\i_m4stg_frac/n713 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[59]  ( .D(\i_m4stg_frac/a0cout[63] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1472), .Q(\i_m4stg_frac/a0c[63] ), 
        .QN(\i_m4stg_frac/n715 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[58]  ( .D(\i_m4stg_frac/a0cout[62] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1472), .Q(\i_m4stg_frac/a0c[62] ), 
        .QN(\i_m4stg_frac/n717 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[57]  ( .D(\i_m4stg_frac/a0cout[61] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1472), .Q(\i_m4stg_frac/a0c[61] ), 
        .QN(\i_m4stg_frac/n719 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[56]  ( .D(\i_m4stg_frac/a0cout[60] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0c[60] ), 
        .QN(\i_m4stg_frac/n721 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[55]  ( .D(\i_m4stg_frac/a0cout[59] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0c[59] ), 
        .QN(\i_m4stg_frac/n723 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[54]  ( .D(\i_m4stg_frac/a0cout[58] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0c[58] ), 
        .QN(\i_m4stg_frac/n725 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[53]  ( .D(\i_m4stg_frac/a0cout[57] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0c[57] ), 
        .QN(\i_m4stg_frac/n727 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[52]  ( .D(\i_m4stg_frac/a0cout[56] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0c[56] ), 
        .QN(\i_m4stg_frac/n729 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[51]  ( .D(\i_m4stg_frac/a0cout[55] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0c[55] ), 
        .QN(\i_m4stg_frac/n731 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[50]  ( .D(\i_m4stg_frac/a0cout[54] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0c[54] ), 
        .QN(\i_m4stg_frac/n733 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[49]  ( .D(\i_m4stg_frac/a0cout[53] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0c[53] ), 
        .QN(\i_m4stg_frac/n735 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[48]  ( .D(\i_m4stg_frac/a0cout[52] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0c[52] ), 
        .QN(\i_m4stg_frac/n737 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[47]  ( .D(\i_m4stg_frac/a0cout[51] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0c[51] ), 
        .QN(\i_m4stg_frac/n739 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[46]  ( .D(\i_m4stg_frac/a0cout[50] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0c[50] ), 
        .QN(\i_m4stg_frac/n741 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[45]  ( .D(\i_m4stg_frac/a0cout[49] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0c[49] ), 
        .QN(\i_m4stg_frac/n743 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[44]  ( .D(\i_m4stg_frac/a0cout[48] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0c[48] ), 
        .QN(\i_m4stg_frac/n745 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[43]  ( .D(\i_m4stg_frac/a0cout[47] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0c[47] ), 
        .QN(\i_m4stg_frac/n747 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[42]  ( .D(\i_m4stg_frac/a0cout[46] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0c[46] ), 
        .QN(\i_m4stg_frac/n749 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[41]  ( .D(\i_m4stg_frac/a0cout[45] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0c[45] ), 
        .QN(\i_m4stg_frac/n751 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[40]  ( .D(\i_m4stg_frac/a0cout[44] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0c[44] ), 
        .QN(\i_m4stg_frac/n753 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[39]  ( .D(\i_m4stg_frac/a0cout[43] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0c[43] ), 
        .QN(\i_m4stg_frac/n755 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[38]  ( .D(\i_m4stg_frac/a0cout[42] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0c[42] ), 
        .QN(\i_m4stg_frac/n757 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[37]  ( .D(\i_m4stg_frac/a0cout[41] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0c[41] ), 
        .QN(\i_m4stg_frac/n759 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[36]  ( .D(\i_m4stg_frac/a0cout[40] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0c[40] ), 
        .QN(\i_m4stg_frac/n761 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[35]  ( .D(\i_m4stg_frac/a0cout[39] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0c[39] ), 
        .QN(\i_m4stg_frac/n763 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[34]  ( .D(\i_m4stg_frac/a0cout[38] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0c[38] ), 
        .QN(\i_m4stg_frac/n765 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[33]  ( .D(\i_m4stg_frac/a0cout[37] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0c[37] ), 
        .QN(\i_m4stg_frac/n767 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[32]  ( .D(\i_m4stg_frac/a0cout[36] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0c[36] ), 
        .QN(\i_m4stg_frac/n769 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[31]  ( .D(\i_m4stg_frac/a0cout[35] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0c[35] ), 
        .QN(\i_m4stg_frac/n771 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[30]  ( .D(\i_m4stg_frac/a0cout[34] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0c[34] ), 
        .QN(\i_m4stg_frac/n773 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[29]  ( .D(\i_m4stg_frac/a0cout[33] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0c[33] ), 
        .QN(\i_m4stg_frac/n775 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[28]  ( .D(\i_m4stg_frac/a0cout[32] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0c[32] ), 
        .QN(\i_m4stg_frac/n777 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[27]  ( .D(\i_m4stg_frac/a0cout[31] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0c[31] ), 
        .QN(\i_m4stg_frac/n779 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[26]  ( .D(\i_m4stg_frac/a0cout[30] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0c[30] ), 
        .QN(\i_m4stg_frac/n781 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[25]  ( .D(\i_m4stg_frac/a0cout[29] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0c[29] ), 
        .QN(\i_m4stg_frac/n783 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[24]  ( .D(\i_m4stg_frac/a0cout[28] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0c[28] ), 
        .QN(\i_m4stg_frac/n785 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[23]  ( .D(\i_m4stg_frac/a0cout[27] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0c[27] ), 
        .QN(\i_m4stg_frac/n787 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[22]  ( .D(\i_m4stg_frac/a0cout[26] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0c[26] ), 
        .QN(\i_m4stg_frac/n789 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[21]  ( .D(\i_m4stg_frac/a0cout[25] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0c[25] ), 
        .QN(\i_m4stg_frac/n791 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[20]  ( .D(\i_m4stg_frac/a0cout[24] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0c[24] ), 
        .QN(\i_m4stg_frac/n793 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[19]  ( .D(\i_m4stg_frac/a0cout[23] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0c[23] ), 
        .QN(\i_m4stg_frac/n795 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[18]  ( .D(\i_m4stg_frac/a0cout[22] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0c[22] ), 
        .QN(\i_m4stg_frac/n797 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[17]  ( .D(\i_m4stg_frac/a0cout[21] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0c[21] ), 
        .QN(\i_m4stg_frac/n799 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[16]  ( .D(\i_m4stg_frac/a0cout[20] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0c[20] ), 
        .QN(\i_m4stg_frac/n801 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[15]  ( .D(\i_m4stg_frac/a0cout[19] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0c[19] ), 
        .QN(\i_m4stg_frac/n803 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[14]  ( .D(\i_m4stg_frac/a0cout[18] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1464), .Q(\i_m4stg_frac/a0c[18] ), 
        .QN(\i_m4stg_frac/n805 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[13]  ( .D(\i_m4stg_frac/a0cout[17] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1464), .Q(\i_m4stg_frac/a0c[17] ), 
        .QN(\i_m4stg_frac/n807 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[12]  ( .D(\i_m4stg_frac/a0cout[16] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1464), .Q(\i_m4stg_frac/a0c[16] ), 
        .QN(\i_m4stg_frac/n809 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[11]  ( .D(\i_m4stg_frac/a0cout[15] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1464), .Q(\i_m4stg_frac/a0c[15] ), 
        .QN(\i_m4stg_frac/n811 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[10]  ( .D(\i_m4stg_frac/a0cout[14] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1464), .Q(n929) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[9]  ( .D(\i_m4stg_frac/a0cout[13] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1463), .Q(n1331), .QN(
        \i_m4stg_frac/n815 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[8]  ( .D(\i_m4stg_frac/a0cout[12] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1463), .Q(\i_m4stg_frac/a0c[12] ), 
        .QN(\i_m4stg_frac/n817 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[7]  ( .D(\i_m4stg_frac/a0cout[11] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1463), .Q(\i_m4stg_frac/a0c[11] ), 
        .QN(\i_m4stg_frac/n819 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[6]  ( .D(\i_m4stg_frac/a0cout[10] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1463), .Q(\i_m4stg_frac/a0c[10] ), 
        .QN(\i_m4stg_frac/n821 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[5]  ( .D(\i_m4stg_frac/a0cout[9] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1463), .Q(\i_m4stg_frac/a0c[9] ), 
        .QN(\i_m4stg_frac/n823 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[4]  ( .D(\i_m4stg_frac/a0cout[8] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1463), .Q(\i_m4stg_frac/a0c[8] ), 
        .QN(\i_m4stg_frac/n825 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[3]  ( .D(\i_m4stg_frac/a0cout[7] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1462), .Q(\i_m4stg_frac/a0c[7] ), 
        .QN(\i_m4stg_frac/n827 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[2]  ( .D(\i_m4stg_frac/a0cout[6] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1462), .Q(n1188) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[1]  ( .D(\i_m4stg_frac/a0cout[5] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1462), .Q(n1329), .QN(
        \i_m4stg_frac/n831 ) );
  DFFSSRX1 \i_m4stg_frac/a0cot_dff/q_reg[0]  ( .D(\i_m4stg_frac/a0cout[4] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1462), .Q(\i_m4stg_frac/a0c[4] ), 
        .QN(\i_m4stg_frac/n833 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[80]  ( .D(1'b1), .RSTB(n1527), .SETB(
        1'b1), .CLK(n1472), .Q(\i_m4stg_frac/a0s[80] ), .QN(
        \i_m4stg_frac/n837 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[79]  ( .D(\i_m4stg_frac/a0sum[79] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1450), .Q(\i_m4stg_frac/a0s[79] ), 
        .QN(\i_m4stg_frac/n839 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[78]  ( .D(\i_m4stg_frac/a0sum[78] ), 
        .RSTB(n1543), .SETB(1'b1), .CLK(n1450), .Q(\i_m4stg_frac/a0s[78] ), 
        .QN(\i_m4stg_frac/n841 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[77]  ( .D(\i_m4stg_frac/a0sum[77] ), 
        .RSTB(n1522), .SETB(1'b1), .CLK(n1450), .Q(\i_m4stg_frac/a0s[77] ), 
        .QN(\i_m4stg_frac/n843 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[76]  ( .D(\i_m4stg_frac/a0sum[76] ), 
        .RSTB(n1522), .SETB(1'b1), .CLK(n1450), .Q(\i_m4stg_frac/a0s[76] ), 
        .QN(\i_m4stg_frac/n845 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[75]  ( .D(\i_m4stg_frac/a0sum[75] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0s[75] ), 
        .QN(\i_m4stg_frac/n847 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[74]  ( .D(\i_m4stg_frac/a0sum[74] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0s[74] ), 
        .QN(\i_m4stg_frac/n849 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[73]  ( .D(\i_m4stg_frac/a0sum[73] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0s[73] ), 
        .QN(\i_m4stg_frac/n851 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[72]  ( .D(\i_m4stg_frac/a0sum[72] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0s[72] ), 
        .QN(\i_m4stg_frac/n853 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[71]  ( .D(\i_m4stg_frac/a0sum[71] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1448), .Q(\i_m4stg_frac/a0s[71] ), 
        .QN(\i_m4stg_frac/n855 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[70]  ( .D(\i_m4stg_frac/a0sum[70] ), 
        .RSTB(n1521), .SETB(1'b1), .CLK(n1449), .Q(\i_m4stg_frac/a0s[70] ), 
        .QN(\i_m4stg_frac/n857 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[69]  ( .D(\i_m4stg_frac/a0sum[69] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1448), .Q(\i_m4stg_frac/a0s[69] ), 
        .QN(\i_m4stg_frac/n859 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[68]  ( .D(\i_m4stg_frac/a0sum[68] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1448), .Q(\i_m4stg_frac/a0s[68] ), 
        .QN(\i_m4stg_frac/n861 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[67]  ( .D(\i_m4stg_frac/a0sum[67] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1448), .Q(n1330), .QN(
        \i_m4stg_frac/n863 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[66]  ( .D(\i_m4stg_frac/a0sum[66] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1448), .Q(\i_m4stg_frac/a0s[66] ), 
        .QN(\i_m4stg_frac/n865 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[65]  ( .D(\i_m4stg_frac/a0sum[65] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1448), .Q(\i_m4stg_frac/a0s[65] ), 
        .QN(\i_m4stg_frac/n867 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[64]  ( .D(\i_m4stg_frac/a0sum[64] ), 
        .RSTB(n1520), .SETB(1'b1), .CLK(n1454), .Q(\i_m4stg_frac/a0s[64] ), 
        .QN(\i_m4stg_frac/n869 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[63]  ( .D(\i_m4stg_frac/a0sum[63] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1472), .Q(\i_m4stg_frac/a0s[63] ), 
        .QN(\i_m4stg_frac/n871 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[62]  ( .D(\i_m4stg_frac/a0sum[62] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1472), .Q(\i_m4stg_frac/a0s[62] ), 
        .QN(\i_m4stg_frac/n873 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[61]  ( .D(\i_m4stg_frac/a0sum[61] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1472), .Q(\i_m4stg_frac/a0s[61] ), 
        .QN(\i_m4stg_frac/n875 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[60]  ( .D(\i_m4stg_frac/a0sum[60] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0s[60] ), 
        .QN(\i_m4stg_frac/n877 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[59]  ( .D(\i_m4stg_frac/a0sum[59] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0s[59] ), 
        .QN(\i_m4stg_frac/n879 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[58]  ( .D(\i_m4stg_frac/a0sum[58] ), 
        .RSTB(n1519), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0s[58] ), 
        .QN(\i_m4stg_frac/n881 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[57]  ( .D(\i_m4stg_frac/a0sum[57] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0s[57] ), 
        .QN(\i_m4stg_frac/n883 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[56]  ( .D(\i_m4stg_frac/a0sum[56] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0s[56] ), 
        .QN(\i_m4stg_frac/n885 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[55]  ( .D(\i_m4stg_frac/a0sum[55] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1471), .Q(\i_m4stg_frac/a0s[55] ), 
        .QN(\i_m4stg_frac/n887 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[54]  ( .D(\i_m4stg_frac/a0sum[54] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0s[54] ), 
        .QN(\i_m4stg_frac/n889 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[53]  ( .D(\i_m4stg_frac/a0sum[53] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0s[53] ), 
        .QN(\i_m4stg_frac/n891 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[52]  ( .D(\i_m4stg_frac/a0sum[52] ), 
        .RSTB(n1518), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0s[52] ), 
        .QN(\i_m4stg_frac/n893 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[51]  ( .D(\i_m4stg_frac/a0sum[51] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0s[51] ), 
        .QN(\i_m4stg_frac/n895 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[50]  ( .D(\i_m4stg_frac/a0sum[50] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0s[50] ), 
        .QN(\i_m4stg_frac/n897 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[49]  ( .D(\i_m4stg_frac/a0sum[49] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1470), .Q(\i_m4stg_frac/a0s[49] ), 
        .QN(\i_m4stg_frac/n899 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[48]  ( .D(\i_m4stg_frac/a0sum[48] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0s[48] ), 
        .QN(\i_m4stg_frac/n901 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[47]  ( .D(\i_m4stg_frac/a0sum[47] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0s[47] ), 
        .QN(\i_m4stg_frac/n903 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[46]  ( .D(\i_m4stg_frac/a0sum[46] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0s[46] ), 
        .QN(\i_m4stg_frac/n905 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[45]  ( .D(\i_m4stg_frac/a0sum[45] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0s[45] ), 
        .QN(\i_m4stg_frac/n907 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[44]  ( .D(\i_m4stg_frac/a0sum[44] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0s[44] ), 
        .QN(\i_m4stg_frac/n909 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[43]  ( .D(\i_m4stg_frac/a0sum[43] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1469), .Q(\i_m4stg_frac/a0s[43] ), 
        .QN(\i_m4stg_frac/n911 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[42]  ( .D(\i_m4stg_frac/a0sum[42] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0s[42] ), 
        .QN(\i_m4stg_frac/n913 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[41]  ( .D(\i_m4stg_frac/a0sum[41] ), 
        .RSTB(n1516), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0s[41] ), 
        .QN(\i_m4stg_frac/n915 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[40]  ( .D(\i_m4stg_frac/a0sum[40] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0s[40] ), 
        .QN(\i_m4stg_frac/n917 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[39]  ( .D(\i_m4stg_frac/a0sum[39] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0s[39] ), 
        .QN(\i_m4stg_frac/n919 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[38]  ( .D(\i_m4stg_frac/a0sum[38] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0s[38] ), 
        .QN(\i_m4stg_frac/n921 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[37]  ( .D(\i_m4stg_frac/a0sum[37] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1468), .Q(\i_m4stg_frac/a0s[37] ), 
        .QN(\i_m4stg_frac/n923 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[36]  ( .D(\i_m4stg_frac/a0sum[36] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0s[36] ), 
        .QN(\i_m4stg_frac/n925 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[35]  ( .D(\i_m4stg_frac/a0sum[35] ), 
        .RSTB(n1515), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0s[35] ), 
        .QN(\i_m4stg_frac/n927 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[34]  ( .D(\i_m4stg_frac/a0sum[34] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0s[34] ), 
        .QN(\i_m4stg_frac/n929 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[33]  ( .D(\i_m4stg_frac/a0sum[33] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0s[33] ), 
        .QN(\i_m4stg_frac/n931 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[32]  ( .D(\i_m4stg_frac/a0sum[32] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0s[32] ), 
        .QN(\i_m4stg_frac/n933 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[31]  ( .D(\i_m4stg_frac/a0sum[31] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1467), .Q(\i_m4stg_frac/a0s[31] ), 
        .QN(\i_m4stg_frac/n935 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[30]  ( .D(\i_m4stg_frac/a0sum[30] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0s[30] ), 
        .QN(\i_m4stg_frac/n937 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[29]  ( .D(\i_m4stg_frac/a0sum[29] ), 
        .RSTB(n1514), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0s[29] ), 
        .QN(\i_m4stg_frac/n939 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[28]  ( .D(\i_m4stg_frac/a0sum[28] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0s[28] ), 
        .QN(\i_m4stg_frac/n941 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[27]  ( .D(\i_m4stg_frac/a0sum[27] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0s[27] ), 
        .QN(\i_m4stg_frac/n943 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[26]  ( .D(\i_m4stg_frac/a0sum[26] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1466), .Q(\i_m4stg_frac/a0s[26] ), 
        .QN(\i_m4stg_frac/n945 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[25]  ( .D(\i_m4stg_frac/a0sum[25] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0s[25] ), 
        .QN(\i_m4stg_frac/n947 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[24]  ( .D(\i_m4stg_frac/a0sum[24] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0s[24] ), 
        .QN(\i_m4stg_frac/n949 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[23]  ( .D(\i_m4stg_frac/a0sum[23] ), 
        .RSTB(n1513), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0s[23] ), 
        .QN(\i_m4stg_frac/n951 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[22]  ( .D(\i_m4stg_frac/a0sum[22] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0s[22] ), 
        .QN(\i_m4stg_frac/n953 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[21]  ( .D(\i_m4stg_frac/a0sum[21] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0s[21] ), 
        .QN(\i_m4stg_frac/n955 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[20]  ( .D(\i_m4stg_frac/a0sum[20] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1465), .Q(\i_m4stg_frac/a0s[20] ), 
        .QN(\i_m4stg_frac/n957 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[19]  ( .D(\i_m4stg_frac/a0sum[19] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1464), .Q(\i_m4stg_frac/a0s[19] ), 
        .QN(\i_m4stg_frac/n959 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[18]  ( .D(\i_m4stg_frac/a0sum[18] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1464), .Q(\i_m4stg_frac/a0s[18] ), 
        .QN(\i_m4stg_frac/n961 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[17]  ( .D(\i_m4stg_frac/a0sum[17] ), 
        .RSTB(n1512), .SETB(1'b1), .CLK(n1464), .Q(\i_m4stg_frac/a0s[17] ), 
        .QN(\i_m4stg_frac/n963 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[16]  ( .D(\i_m4stg_frac/a0sum[16] ), 
        .RSTB(n1517), .SETB(1'b1), .CLK(n1464), .Q(\i_m4stg_frac/a0s[16] ), 
        .QN(\i_m4stg_frac/n965 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[15]  ( .D(\i_m4stg_frac/a0sum[15] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1464), .Q(n1189) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[14]  ( .D(\i_m4stg_frac/a0sum[14] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1464), .Q(n1192), .QN(
        \i_m4stg_frac/n969 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[13]  ( .D(\i_m4stg_frac/a0sum[13] ), 
        .RSTB(n1532), .SETB(1'b1), .CLK(n1464), .Q(n1112) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[12]  ( .D(\i_m4stg_frac/a0sum[12] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1463), .Q(n1072) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[11]  ( .D(\i_m4stg_frac/a0sum[11] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1463), .Q(n1060) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[10]  ( .D(\i_m4stg_frac/a0sum[10] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1463), .Q(n1069) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[9]  ( .D(\i_m4stg_frac/a0sum[9] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1463), .Q(n1070) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[8]  ( .D(\i_m4stg_frac/a0sum[8] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1463), .Q(n1071) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[7]  ( .D(\i_m4stg_frac/a0sum[7] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1463), .Q(n1068) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[6]  ( .D(\i_m4stg_frac/a0sum[6] ), 
        .RSTB(n1531), .SETB(1'b1), .CLK(n1462), .Q(n1190), .QN(
        \i_m4stg_frac/n985 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[5]  ( .D(\i_m4stg_frac/a0sum[5] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1462), .Q(n1073) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[4]  ( .D(\i_m4stg_frac/a0sum[4] ), 
        .RSTB(n1530), .SETB(1'b1), .CLK(n1462), .Q(n1184), .QN(
        \i_m4stg_frac/n989 ) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[3]  ( .D(\i_m4stg_frac/a0sum[3] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1461), .Q(n1131) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[2]  ( .D(\i_m4stg_frac/a0sum[2] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1460), .Q(n1125) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[1]  ( .D(\i_m4stg_frac/a0sum[1] ), 
        .RSTB(n1528), .SETB(1'b1), .CLK(n1460), .Q(n1120) );
  DFFSSRX1 \i_m4stg_frac/a0sum_dff/q_reg[0]  ( .D(\i_m4stg_frac/a0sum[0] ), 
        .RSTB(n1529), .SETB(1'b1), .CLK(n1460), .Q(n1185), .QN(
        \i_m4stg_frac/n997 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff7/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff7/N5 ), .CLK(n1486), .Q(
        \i_m4stg_frac/b7[2] ), .QN(\i_m4stg_frac/n998 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff7/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff7/N4 ), .CLK(n1486), .Q(n976), .QN(
        \i_m4stg_frac/n999 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff7/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff7/N3 ), .CLK(n1486), .Q(n1196), .QN(
        \i_m4stg_frac/n1000 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff6/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff6/N5 ), .CLK(n1487), .Q(n1038), .QN(
        \i_m4stg_frac/n1001 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff6/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff6/N4 ), .CLK(n1487), .Q(n1229), .QN(
        \i_m4stg_frac/n1002 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff6/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff6/N3 ), .CLK(n1487), .Q(
        \i_m4stg_frac/b6[0] ), .QN(\i_m4stg_frac/n1003 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff5/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff5/N5 ), .CLK(n1487), .Q(n936), .QN(
        \i_m4stg_frac/n1004 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff5/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff5/N4 ), .CLK(n1487), .Q(n1145) );
  DFFX1 \i_m4stg_frac/booth/out_dff5/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff5/N3 ), .CLK(n1487), .Q(n951), .QN(
        \i_m4stg_frac/n1006 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff4/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff4/N5 ), .CLK(n1487), .Q(
        \i_m4stg_frac/b4[2] ), .QN(\i_m4stg_frac/n1007 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff4/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff4/N4 ), .CLK(n1487), .Q(n1118), .QN(
        \i_m4stg_frac/n1008 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff4/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff4/N3 ), .CLK(n1487), .Q(n915), .QN(
        \i_m4stg_frac/n1009 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff3/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff3/N5 ), .CLK(n1487), .Q(n913), .QN(
        \i_m4stg_frac/n1010 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff3/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff3/N4 ), .CLK(n1487), .Q(n1169), .QN(
        \i_m4stg_frac/n1011 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff3/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff3/N3 ), .CLK(n1487), .Q(
        \i_m4stg_frac/b3[0] ), .QN(\i_m4stg_frac/n1012 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff2/q_reg[2]  ( .D(
        \i_m4stg_frac/booth/out_dff2/N5 ), .CLK(n1488), .Q(n935), .QN(
        \i_m4stg_frac/n1013 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff2/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff2/N4 ), .CLK(n1487), .Q(n1144) );
  DFFX1 \i_m4stg_frac/booth/out_dff2/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff2/N3 ), .CLK(n1487), .Q(n950), .QN(
        \i_m4stg_frac/n1015 ) );
  DFFSSRX1 \i_m4stg_frac/booth/out_dff1/q_reg[2]  ( .D(\i_m4stg_frac/n850 ), 
        .RSTB(m2stg_frac2_array_in[3]), .SETB(\i_m4stg_frac/n1684 ), .CLK(
        n1460), .Q(\i_m4stg_frac/b1[2] ), .QN(\i_m4stg_frac/n1016 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff1/q_reg[1]  ( .D(
        \i_m4stg_frac/booth/out_dff1/N4 ), .CLK(n1490), .Q(n933), .QN(
        \i_m4stg_frac/n1017 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff1/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff1/N3 ), .CLK(n1490), .Q(n1135), .QN(
        \i_m4stg_frac/n1018 ) );
  DFFSSRX1 \i_m4stg_frac/booth/out_dff0/q_reg[2]  ( .D(\i_m4stg_frac/n1285 ), 
        .RSTB(\i_m4stg_frac/booth/b0_in1[2] ), .SETB(\i_m4stg_frac/n1692 ), 
        .CLK(n1460), .Q(n1053), .QN(\i_m4stg_frac/n1019 ) );
  DFFSSRX1 \i_m4stg_frac/booth/out_dff0/q_reg[1]  ( .D(\i_m4stg_frac/n850 ), 
        .RSTB(m2stg_frac2_array_in[1]), .SETB(\i_m4stg_frac/n1693 ), .CLK(
        n1460), .Q(n1327), .QN(\i_m4stg_frac/n1020 ) );
  DFFX1 \i_m4stg_frac/booth/out_dff0/q_reg[0]  ( .D(
        \i_m4stg_frac/booth/out_dff0/N3 ), .CLK(n1490), .Q(
        \i_m4stg_frac/b0[0] ), .QN(\i_m4stg_frac/n1021 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[20]  ( .D(
        m2stg_frac2_array_in[52]), .RSTB(n1528), .SETB(1'b1), .CLK(n1355), .Q(
        n1278) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[19]  ( .D(
        m2stg_frac2_array_in[51]), .RSTB(n1525), .SETB(1'b1), .CLK(n1353), .Q(
        n1161), .QN(\i_m4stg_frac/n215 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[18]  ( .D(
        m2stg_frac2_array_in[50]), .RSTB(n1528), .SETB(1'b1), .CLK(n1356), .Q(
        \i_m4stg_frac/booth/b[50] ), .QN(\i_m4stg_frac/n334 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[17]  ( .D(
        m2stg_frac2_array_in[49]), .RSTB(n1525), .SETB(1'b1), .CLK(n1354), .Q(
        \i_m4stg_frac/n201 ), .QN(n1172) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[16]  ( .D(
        m2stg_frac2_array_in[48]), .RSTB(n1528), .SETB(1'b1), .CLK(n1353), .Q(
        \i_m4stg_frac/booth/b[48] ), .QN(\i_m4stg_frac/n343 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[15]  ( .D(
        m2stg_frac2_array_in[47]), .RSTB(n1525), .SETB(1'b1), .CLK(n1355), .Q(
        \i_m4stg_frac/n211 ), .QN(n944) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[14]  ( .D(
        m2stg_frac2_array_in[46]), .RSTB(n1528), .SETB(1'b1), .CLK(n1354), .Q(
        n1323), .QN(\i_m4stg_frac/n341 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[13]  ( .D(
        m2stg_frac2_array_in[45]), .RSTB(n1525), .SETB(1'b1), .CLK(n1356), .Q(
        \i_m4stg_frac/n205 ), .QN(n1173) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[12]  ( .D(
        m2stg_frac2_array_in[44]), .RSTB(n1528), .SETB(1'b1), .CLK(n1355), .Q(
        \i_m4stg_frac/booth/b[44] ), .QN(\i_m4stg_frac/n339 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[11]  ( .D(
        m2stg_frac2_array_in[43]), .RSTB(n1525), .SETB(1'b1), .CLK(n1353), .Q(
        \i_m4stg_frac/n209 ), .QN(n945) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[10]  ( .D(
        m2stg_frac2_array_in[42]), .RSTB(n1523), .SETB(1'b1), .CLK(n1354), .Q(
        n1324), .QN(\i_m4stg_frac/n337 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[9]  ( .D(m2stg_frac2_array_in[41]), .RSTB(n1523), .SETB(1'b1), .CLK(n1355), .Q(\i_m4stg_frac/n203 ), .QN(n946)
         );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[8]  ( .D(m2stg_frac2_array_in[40]), .RSTB(n1523), .SETB(1'b1), .CLK(n1356), .Q(n1325), .QN(\i_m4stg_frac/n336 )
         );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[7]  ( .D(m2stg_frac2_array_in[39]), .RSTB(n1523), .SETB(1'b1), .CLK(n1353), .Q(\i_m4stg_frac/n199 ), .QN(n1174)
         );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[6]  ( .D(m2stg_frac2_array_in[38]), .RSTB(n1522), .SETB(1'b1), .CLK(n1354), .Q(\i_m4stg_frac/booth/b[38] ), .QN(
        \i_m4stg_frac/n335 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[5]  ( .D(m2stg_frac2_array_in[37]), .RSTB(n1522), .SETB(1'b1), .CLK(n1355), .Q(\i_m4stg_frac/n213 ), .QN(n1127)
         );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[4]  ( .D(m2stg_frac2_array_in[36]), .RSTB(n1522), .SETB(1'b1), .CLK(n1356), .Q(\i_m4stg_frac/booth/b[36] ), .QN(
        \i_m4stg_frac/n1277 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[3]  ( .D(m2stg_frac2_array_in[35]), .RSTB(n1522), .SETB(1'b1), .CLK(n1353), .Q(\i_m4stg_frac/n333 ), .QN(n1352)
         );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[2]  ( .D(m2stg_frac2_array_in[34]), .RSTB(n1522), .SETB(1'b1), .CLK(n1354), .Q(\i_m4stg_frac/booth/b[34] ), .QN(
        \i_m4stg_frac/n1281 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[1]  ( .D(m2stg_frac2_array_in[33]), .RSTB(n1522), .SETB(1'b1), .CLK(n1355), .Q(\i_m4stg_frac/booth/b0_in1[2] ), 
        .QN(\i_m4stg_frac/n207 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff/q_reg[0]  ( .D(m2stg_frac2_array_in[32]), .RSTB(n1522), .SETB(1'b1), .CLK(n1356), .Q(\i_m4stg_frac/n300 ), .QN(
        \i_m4stg_frac/n1532 ) );
  DFFSSRX1 \i_m4stg_frac/booth/hld_dff0/q_reg[0]  ( .D(n1538), .RSTB(
        m2stg_frac2_array_in[31]), .SETB(1'b1), .CLK(n1353), .Q(
        \i_m4stg_frac/booth/b[31] ), .QN(\i_m4stg_frac/n345 ) );
  LATCHX1 \i_m4stg_frac/booth/ckbuf_1/clken_reg  ( .CLK(n709), .D(
        \i_m4stg_frac/ckbuf_1/N1 ), .Q(\i_m4stg_frac/booth/ckbuf_1/clken ), 
        .QN(\i_m4stg_frac/n1055 ) );
  LATCHX1 \i_m4stg_frac/booth/ckbuf_0/clken_reg  ( .CLK(n709), .D(
        \i_m4stg_frac/ckbuf_0/N1 ), .Q(\i_m4stg_frac/booth/ckbuf_0/clken ), 
        .QN(\i_m4stg_frac/n1056 ) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[31]  ( .D(m4stg_frac[63]), .RSTB(n1534), 
        .SETB(1'b1), .CLK(n1473), .Q(m4stg_frac[31]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[30]  ( .D(m4stg_frac[62]), .RSTB(n1534), 
        .SETB(1'b1), .CLK(n1473), .Q(m4stg_frac[30]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[29]  ( .D(m4stg_frac[61]), .RSTB(n1534), 
        .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[29]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[28]  ( .D(m4stg_frac[60]), .RSTB(n1534), 
        .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[28]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[27]  ( .D(m4stg_frac[59]), .RSTB(n1534), 
        .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[27]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[26]  ( .D(m4stg_frac[58]), .RSTB(n1512), 
        .SETB(1'b1), .CLK(n1448), .Q(m4stg_frac[26]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[25]  ( .D(m4stg_frac[57]), .RSTB(n1541), 
        .SETB(1'b1), .CLK(n1481), .Q(m4stg_frac[25]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[24]  ( .D(m4stg_frac[56]), .RSTB(n1541), 
        .SETB(1'b1), .CLK(n1480), .Q(m4stg_frac[24]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[23]  ( .D(m4stg_frac[55]), .RSTB(n1540), 
        .SETB(1'b1), .CLK(n1481), .Q(m4stg_frac[23]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[22]  ( .D(m4stg_frac[54]), .RSTB(n1540), 
        .SETB(1'b1), .CLK(n1480), .Q(m4stg_frac[22]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[21]  ( .D(m4stg_frac[53]), .RSTB(n1540), 
        .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[21]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[20]  ( .D(m4stg_frac[52]), .RSTB(n1540), 
        .SETB(1'b1), .CLK(n1480), .Q(m4stg_frac[20]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[19]  ( .D(m4stg_frac[51]), .RSTB(n1540), 
        .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[19]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[18]  ( .D(m4stg_frac[50]), .RSTB(n1540), 
        .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[18]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[17]  ( .D(m4stg_frac[49]), .RSTB(n1539), 
        .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[17]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[16]  ( .D(m4stg_frac[48]), .RSTB(n1539), 
        .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[16]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[15]  ( .D(m4stg_frac[47]), .RSTB(n1539), 
        .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[15]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[14]  ( .D(m4stg_frac[46]), .RSTB(n1539), 
        .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[14]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[13]  ( .D(m4stg_frac[45]), .RSTB(n1539), 
        .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[13]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[12]  ( .D(m4stg_frac[44]), .RSTB(n1539), 
        .SETB(1'b1), .CLK(n1477), .Q(m4stg_frac[12]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[11]  ( .D(m4stg_frac[43]), .RSTB(n1538), 
        .SETB(1'b1), .CLK(n1477), .Q(m4stg_frac[11]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[10]  ( .D(m4stg_frac[42]), .RSTB(n1538), 
        .SETB(1'b1), .CLK(n1477), .Q(m4stg_frac[10]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[9]  ( .D(m4stg_frac[41]), .RSTB(n1541), 
        .SETB(1'b1), .CLK(n1481), .Q(m4stg_frac[9]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[8]  ( .D(m4stg_frac[40]), .RSTB(n1541), 
        .SETB(1'b1), .CLK(n1481), .Q(m4stg_frac[8]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[7]  ( .D(m4stg_frac[39]), .RSTB(n1541), 
        .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[7]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[6]  ( .D(m4stg_frac[38]), .RSTB(n1541), 
        .SETB(1'b1), .CLK(n1481), .Q(m4stg_frac[6]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[5]  ( .D(m4stg_frac[37]), .RSTB(n1542), 
        .SETB(1'b1), .CLK(n1480), .Q(m4stg_frac[5]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[4]  ( .D(m4stg_frac[36]), .RSTB(n1542), 
        .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[4]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[3]  ( .D(m4stg_frac[35]), .RSTB(n1542), 
        .SETB(1'b1), .CLK(n1481), .Q(m4stg_frac[3]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[2]  ( .D(m4stg_frac[34]), .RSTB(n1542), 
        .SETB(1'b1), .CLK(n1483), .Q(m4stg_frac[2]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[1]  ( .D(m4stg_frac[33]), .RSTB(n1542), 
        .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[1]) );
  DFFSSRX1 \i_m4stg_frac/pip_dff/q_reg[0]  ( .D(m4stg_frac[32]), .RSTB(n1542), 
        .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[0]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[73]  ( .D(\i_m4stg_frac/addout[73] ), 
        .RSTB(n1538), .SETB(1'b1), .CLK(n1477), .Q(m4stg_frac_105), .QN(n979)
         );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[72]  ( .D(\i_m4stg_frac/addout[72] ), 
        .RSTB(n1538), .SETB(1'b1), .CLK(n1477), .Q(m4stg_frac[104]), .QN(n1230) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[71]  ( .D(\i_m4stg_frac/addout[71] ), 
        .RSTB(n1538), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[103]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[70]  ( .D(\i_m4stg_frac/addout[70] ), 
        .RSTB(n1538), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[102]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[69]  ( .D(\i_m4stg_frac/addout[69] ), 
        .RSTB(n1538), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[101]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[68]  ( .D(\i_m4stg_frac/addout[68] ), 
        .RSTB(n1538), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[100]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[67]  ( .D(\i_m4stg_frac/addout[67] ), 
        .RSTB(n1538), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[99]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[66]  ( .D(\i_m4stg_frac/addout[66] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[98]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[65]  ( .D(\i_m4stg_frac/addout[65] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[97]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[64]  ( .D(\i_m4stg_frac/addout[64] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[96]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[63]  ( .D(\i_m4stg_frac/addout[63] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[95]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[62]  ( .D(\i_m4stg_frac/addout[62] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[94]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[61]  ( .D(\i_m4stg_frac/addout[61] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[93]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[60]  ( .D(\i_m4stg_frac/addout[60] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1476), .Q(m4stg_frac[92]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[59]  ( .D(\i_m4stg_frac/addout[59] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[91]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[58]  ( .D(\i_m4stg_frac/addout[58] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[90]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[57]  ( .D(\i_m4stg_frac/addout[57] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[89]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[56]  ( .D(\i_m4stg_frac/addout[56] ), 
        .RSTB(n1537), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[88]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[55]  ( .D(\i_m4stg_frac/addout[55] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[87]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[54]  ( .D(\i_m4stg_frac/addout[54] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[86]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[53]  ( .D(\i_m4stg_frac/addout[53] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[85]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[52]  ( .D(\i_m4stg_frac/addout[52] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[84]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[51]  ( .D(\i_m4stg_frac/addout[51] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[83]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[50]  ( .D(\i_m4stg_frac/addout[50] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[82]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[49]  ( .D(\i_m4stg_frac/addout[49] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[81]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[48]  ( .D(\i_m4stg_frac/addout[48] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1475), .Q(m4stg_frac[80]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[47]  ( .D(\i_m4stg_frac/addout[47] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[79]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[46]  ( .D(\i_m4stg_frac/addout[46] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[78]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[45]  ( .D(\i_m4stg_frac/addout[45] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[77]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[44]  ( .D(\i_m4stg_frac/addout[44] ), 
        .RSTB(n1536), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[76]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[43]  ( .D(\i_m4stg_frac/addout[43] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[75]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[42]  ( .D(\i_m4stg_frac/addout[42] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[74]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[41]  ( .D(\i_m4stg_frac/addout[41] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[73]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[40]  ( .D(\i_m4stg_frac/addout[40] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[72]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[39]  ( .D(\i_m4stg_frac/addout[39] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[71]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[38]  ( .D(\i_m4stg_frac/addout[38] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[70]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[37]  ( .D(\i_m4stg_frac/addout[37] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1474), .Q(m4stg_frac[69]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[36]  ( .D(\i_m4stg_frac/addout[36] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1473), .Q(m4stg_frac[68]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[35]  ( .D(\i_m4stg_frac/addout[35] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1473), .Q(m4stg_frac[67]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[34]  ( .D(\i_m4stg_frac/addout[34] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1473), .Q(m4stg_frac[66]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[33]  ( .D(\i_m4stg_frac/addout[33] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1473), .Q(m4stg_frac[65]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[32]  ( .D(\i_m4stg_frac/addout[32] ), 
        .RSTB(n1535), .SETB(1'b1), .CLK(n1473), .Q(m4stg_frac[64]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[31]  ( .D(\i_m4stg_frac/addout[31] ), 
        .RSTB(n1534), .SETB(1'b1), .CLK(n1473), .Q(m4stg_frac[63]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[30]  ( .D(\i_m4stg_frac/addout[30] ), 
        .RSTB(n1534), .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[62]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[29]  ( .D(\i_m4stg_frac/addout[29] ), 
        .RSTB(n1534), .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[61]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[28]  ( .D(\i_m4stg_frac/addout[28] ), 
        .RSTB(n1534), .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[60]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[27]  ( .D(\i_m4stg_frac/addout[27] ), 
        .RSTB(n1534), .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[59]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[26]  ( .D(\i_m4stg_frac/addout[26] ), 
        .RSTB(n1542), .SETB(1'b1), .CLK(n1477), .Q(m4stg_frac[58]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[25]  ( .D(\i_m4stg_frac/addout[25] ), 
        .RSTB(n1541), .SETB(1'b1), .CLK(n1480), .Q(m4stg_frac[57]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[24]  ( .D(\i_m4stg_frac/addout[24] ), 
        .RSTB(n1540), .SETB(1'b1), .CLK(n1481), .Q(m4stg_frac[56]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[23]  ( .D(\i_m4stg_frac/addout[23] ), 
        .RSTB(n1540), .SETB(1'b1), .CLK(n1481), .Q(m4stg_frac[55]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[22]  ( .D(\i_m4stg_frac/addout[22] ), 
        .RSTB(n1540), .SETB(1'b1), .CLK(n1480), .Q(m4stg_frac[54]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[21]  ( .D(\i_m4stg_frac/addout[21] ), 
        .RSTB(n1540), .SETB(1'b1), .CLK(n1480), .Q(m4stg_frac[53]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[20]  ( .D(\i_m4stg_frac/addout[20] ), 
        .RSTB(n1540), .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[52]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[19]  ( .D(\i_m4stg_frac/addout[19] ), 
        .RSTB(n1540), .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[51]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[18]  ( .D(\i_m4stg_frac/addout[18] ), 
        .RSTB(n1539), .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[50]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[17]  ( .D(\i_m4stg_frac/addout[17] ), 
        .RSTB(n1539), .SETB(1'b1), .CLK(n1479), .Q(m4stg_frac[49]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[16]  ( .D(\i_m4stg_frac/addout[16] ), 
        .RSTB(n1539), .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[48]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[15]  ( .D(\i_m4stg_frac/addout[15] ), 
        .RSTB(n1539), .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[47]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[14]  ( .D(\i_m4stg_frac/addout[14] ), 
        .RSTB(n1539), .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[46]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[13]  ( .D(\i_m4stg_frac/addout[13] ), 
        .RSTB(n1539), .SETB(1'b1), .CLK(n1478), .Q(m4stg_frac[45]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[12]  ( .D(\i_m4stg_frac/addout[12] ), 
        .RSTB(n1538), .SETB(1'b1), .CLK(n1477), .Q(m4stg_frac[44]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[11]  ( .D(\i_m4stg_frac/addout[11] ), 
        .RSTB(n1538), .SETB(1'b1), .CLK(n1477), .Q(m4stg_frac[43]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[10]  ( .D(\i_m4stg_frac/addout[10] ), 
        .RSTB(n1538), .SETB(1'b1), .CLK(n1477), .Q(m4stg_frac[42]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[9]  ( .D(\i_m4stg_frac/addout[9] ), 
        .RSTB(n1541), .SETB(1'b1), .CLK(n1481), .Q(m4stg_frac[41]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[8]  ( .D(\i_m4stg_frac/addout[8] ), 
        .RSTB(n1541), .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[40]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[7]  ( .D(\i_m4stg_frac/addout[7] ), 
        .RSTB(n1541), .SETB(1'b1), .CLK(n1481), .Q(m4stg_frac[39]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[6]  ( .D(\i_m4stg_frac/addout[6] ), 
        .RSTB(n1541), .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[38]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[5]  ( .D(\i_m4stg_frac/addout[5] ), 
        .RSTB(n1541), .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[37]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[4]  ( .D(\i_m4stg_frac/addout[4] ), 
        .RSTB(n1542), .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[36]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[3]  ( .D(\i_m4stg_frac/addout[3] ), 
        .RSTB(n1542), .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[35]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[2]  ( .D(\i_m4stg_frac/addout[2] ), 
        .RSTB(n1542), .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[34]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[1]  ( .D(\i_m4stg_frac/addout[1] ), 
        .RSTB(n1542), .SETB(1'b1), .CLK(n1482), .Q(m4stg_frac[33]) );
  DFFSSRX1 \i_m4stg_frac/out_dff/q_reg[0]  ( .D(\i_m4stg_frac/addout[0] ), 
        .RSTB(n1542), .SETB(1'b1), .CLK(n1483), .Q(m4stg_frac[32]) );
  DFFX1 \i_m4stg_frac/co31_dff/q_reg[0]  ( .D(\i_m4stg_frac/co31_dff/N3 ), 
        .CLK(n1486), .Q(\i_m4stg_frac/addin_cin ), .QN(\i_m4stg_frac/n1329 )
         );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[63]  ( .D(1'b1), .RSTB(n1525), .SETB(1'b1), .CLK(n1356), .Q(n907), .QN(\i_m4stg_frac/n1530 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[52]  ( .D(m2stg_frac1_array_in[52]), 
        .RSTB(n1528), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1519 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[51]  ( .D(m2stg_frac1_array_in[51]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1518 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[50]  ( .D(m2stg_frac1_array_in[50]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1517 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[49]  ( .D(m2stg_frac1_array_in[49]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1516 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[48]  ( .D(m2stg_frac1_array_in[48]), 
        .RSTB(n1528), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1515 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[47]  ( .D(m2stg_frac1_array_in[47]), 
        .RSTB(n1528), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1514 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[46]  ( .D(m2stg_frac1_array_in[46]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1513 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[45]  ( .D(m2stg_frac1_array_in[45]), 
        .RSTB(n1528), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1512 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[44]  ( .D(m2stg_frac1_array_in[44]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1511 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[43]  ( .D(m2stg_frac1_array_in[43]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1510 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[42]  ( .D(m2stg_frac1_array_in[42]), 
        .RSTB(n1528), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1509 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[41]  ( .D(m2stg_frac1_array_in[41]), 
        .RSTB(n1528), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1508 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[40]  ( .D(m2stg_frac1_array_in[40]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1507 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[39]  ( .D(m2stg_frac1_array_in[39]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1506 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[38]  ( .D(m2stg_frac1_array_in[38]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1505 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[37]  ( .D(m2stg_frac1_array_in[37]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1504 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[36]  ( .D(m2stg_frac1_array_in[36]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1503 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[35]  ( .D(m2stg_frac1_array_in[35]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1502 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[34]  ( .D(m2stg_frac1_array_in[34]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1501 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[33]  ( .D(m2stg_frac1_array_in[33]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1500 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[32]  ( .D(m2stg_frac1_array_in[32]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1499 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[31]  ( .D(m2stg_frac1_array_in[31]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1498 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[30]  ( .D(m2stg_frac1_array_in[30]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1497 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[29]  ( .D(m2stg_frac1_array_in[29]), 
        .RSTB(n1524), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1496 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[28]  ( .D(m2stg_frac1_array_in[28]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1495 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[27]  ( .D(m2stg_frac1_array_in[27]), 
        .RSTB(n1526), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1494 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[26]  ( .D(m2stg_frac1_array_in[26]), 
        .RSTB(n1526), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1493 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[25]  ( .D(m2stg_frac1_array_in[25]), 
        .RSTB(n1523), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1492 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[24]  ( .D(m2stg_frac1_array_in[24]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1491 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[23]  ( .D(m2stg_frac1_array_in[23]), 
        .RSTB(n1523), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1490 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[22]  ( .D(m2stg_frac1_array_in[22]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1489 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[21]  ( .D(m2stg_frac1_array_in[21]), 
        .RSTB(n1523), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1488 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[20]  ( .D(m2stg_frac1_array_in[20]), 
        .RSTB(n1523), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1487 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[19]  ( .D(m2stg_frac1_array_in[19]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1486 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[18]  ( .D(m2stg_frac1_array_in[18]), 
        .RSTB(n1523), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1485 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[17]  ( .D(m2stg_frac1_array_in[17]), 
        .RSTB(n1527), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1484 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[16]  ( .D(m2stg_frac1_array_in[16]), 
        .RSTB(n1523), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1483 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[15]  ( .D(m2stg_frac1_array_in[15]), 
        .RSTB(n1526), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1482 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[14]  ( .D(m2stg_frac1_array_in[14]), 
        .RSTB(n1523), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1481 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[13]  ( .D(m2stg_frac1_array_in[13]), 
        .RSTB(n1523), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1480 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[12]  ( .D(m2stg_frac1_array_in[12]), 
        .RSTB(n1526), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1479 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[11]  ( .D(m2stg_frac1_array_in[11]), 
        .RSTB(n1526), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1478 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[10]  ( .D(m2stg_frac1_array_in[10]), 
        .RSTB(n1526), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1477 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[9]  ( .D(m2stg_frac1_array_in[9]), .RSTB(
        n1526), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1476 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[8]  ( .D(m2stg_frac1_array_in[8]), .RSTB(
        n1526), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1475 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[7]  ( .D(m2stg_frac1_array_in[7]), .RSTB(
        n1526), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1474 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[6]  ( .D(m2stg_frac1_array_in[6]), .RSTB(
        n1526), .SETB(1'b1), .CLK(n1356), .QN(\i_m4stg_frac/n1473 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[5]  ( .D(m2stg_frac1_array_in[5]), .RSTB(
        n1526), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1472 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[4]  ( .D(m2stg_frac1_array_in[4]), .RSTB(
        n1526), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1471 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[3]  ( .D(m2stg_frac1_array_in[3]), .RSTB(
        n1525), .SETB(1'b1), .CLK(n1355), .QN(\i_m4stg_frac/n1470 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[2]  ( .D(m2stg_frac1_array_in[2]), .RSTB(
        n1525), .SETB(1'b1), .CLK(n1354), .QN(\i_m4stg_frac/n1469 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[1]  ( .D(m2stg_frac1_array_in[1]), .RSTB(
        n1525), .SETB(1'b1), .CLK(n1353), .QN(\i_m4stg_frac/n1468 ) );
  DFFSSRX1 \i_m4stg_frac/ffrs1/q_reg[0]  ( .D(m2stg_frac1_array_in[0]), .RSTB(
        n1525), .SETB(1'b1), .CLK(n1356), .Q(n1034), .QN(\i_m4stg_frac/n1467 )
         );
  DFFX1 \i_m4stg_frac/cyc3_dff/q_reg[0]  ( .D(\i_m4stg_frac/cyc3_dff/N7 ), 
        .CLK(n1490), .Q(\i_m4stg_frac/cyc3 ), .QN(\i_m4stg_frac/n1462 ) );
  DFFX1 \i_m4stg_frac/cyc2_dff/q_reg[0]  ( .D(\i_m4stg_frac/cyc2_dff/N7 ), 
        .CLK(n1490), .Q(\i_m4stg_frac/a1sum[81] ) );
  DFFX1 \i_m4stg_frac/cyc1_dff/q_reg[0]  ( .D(\i_m4stg_frac/cyc1_dff/N7 ), 
        .CLK(n1490), .Q(\i_m4stg_frac/cyc1 ), .QN(\i_m4stg_frac/n1464 ) );
  OR2X1 U669 ( .IN1(\i_m4stg_frac/n1056 ), .IN2(n709), .Q(n911) );
  OR2X1 U670 ( .IN1(n1033), .IN2(\fpu_mul_frac_dp/n833 ), .Q(n1041) );
  OR2X1 U671 ( .IN1(n906), .IN2(\fpu_mul_frac_dp/n765 ), .Q(n1049) );
  OR2X1 U672 ( .IN1(\fpu_mul_frac_dp/n765 ), .IN2(\fpu_mul_frac_dp/n833 ), .Q(
        n1050) );
  AND2X1 U673 ( .IN1(\i_m4stg_frac/n854 ), .IN2(\i_m4stg_frac/a1sum[81] ), .Q(
        n1052) );
  OR2X1 U674 ( .IN1(\i_m4stg_frac/n1055 ), .IN2(n709), .Q(n1057) );
  INVX0 U675 ( .INP(n1057), .ZN(n1353) );
  INVX0 U676 ( .INP(n1057), .ZN(n1354) );
  INVX0 U677 ( .INP(n1057), .ZN(n1355) );
  INVX0 U678 ( .INP(n1057), .ZN(n1356) );
  INVX0 U679 ( .INP(se_mul), .ZN(n1357) );
  INVX0 U680 ( .INP(se_mul), .ZN(n1358) );
  INVX0 U681 ( .INP(se_mul), .ZN(n1359) );
  INVX0 U682 ( .INP(se_mul), .ZN(n1360) );
  INVX0 U683 ( .INP(n1050), .ZN(n1361) );
  INVX0 U684 ( .INP(n1050), .ZN(n1362) );
  INVX0 U685 ( .INP(n1050), .ZN(n1363) );
  INVX0 U686 ( .INP(n1050), .ZN(n1364) );
  INVX0 U687 ( .INP(n1049), .ZN(n1365) );
  INVX0 U688 ( .INP(n1049), .ZN(n1366) );
  INVX0 U689 ( .INP(n1049), .ZN(n1367) );
  INVX0 U690 ( .INP(n1049), .ZN(n1368) );
  INVX0 U691 ( .INP(n1041), .ZN(n1369) );
  INVX0 U692 ( .INP(n1041), .ZN(n1370) );
  INVX0 U693 ( .INP(n1041), .ZN(n1371) );
  INVX0 U694 ( .INP(n1041), .ZN(n1372) );
  INVX0 U695 ( .INP(n1052), .ZN(n1373) );
  INVX0 U696 ( .INP(n1052), .ZN(n1374) );
  INVX0 U697 ( .INP(n1052), .ZN(n1375) );
  INVX0 U698 ( .INP(n1052), .ZN(n1376) );
  INVX0 U699 ( .INP(n9304), .ZN(n1377) );
  INVX0 U700 ( .INP(n9304), .ZN(n1378) );
  INVX0 U701 ( .INP(n9304), .ZN(n1379) );
  INVX0 U702 ( .INP(n9304), .ZN(n1380) );
  NAND3X1 U703 ( .IN1(\i_m4stg_frac/n654 ), .IN2(n938), .IN3(
        \i_m4stg_frac/n656 ), .QN(n3759) );
  NAND2X1 U704 ( .IN1(n3820), .IN2(n1040), .QN(n3587) );
  NAND2X1 U705 ( .IN1(n3614), .IN2(n1039), .QN(n3781) );
  NAND2X1 U706 ( .IN1(n6541), .IN2(n1038), .QN(n6361) );
  NAND2X1 U707 ( .IN1(n3670), .IN2(n912), .QN(n3567) );
  NAND2X1 U708 ( .IN1(n6418), .IN2(n913), .QN(n6312) );
  NAND2X1 U709 ( .IN1(n6569), .IN2(n1053), .QN(n6332) );
  NAND3X1 U710 ( .IN1(\i_m4stg_frac/n657 ), .IN2(n1133), .IN3(
        \i_m4stg_frac/n659 ), .QN(n3818) );
  NAND3X1 U711 ( .IN1(\i_m4stg_frac/n675 ), .IN2(n1134), .IN3(
        \i_m4stg_frac/n677 ), .QN(n3586) );
  NAND3X1 U712 ( .IN1(\i_m4stg_frac/n1016 ), .IN2(n933), .IN3(
        \i_m4stg_frac/n1018 ), .QN(n6337) );
  NAND3X1 U713 ( .IN1(n1196), .IN2(n976), .IN3(\i_m4stg_frac/n998 ), .QN(n6492) );
  NAND3X1 U714 ( .IN1(n938), .IN2(n1123), .IN3(\i_m4stg_frac/n654 ), .QN(n3742) );
  NAND3X1 U715 ( .IN1(n1116), .IN2(n914), .IN3(\i_m4stg_frac/n663 ), .QN(n3891) );
  NAND3X1 U716 ( .IN1(n1118), .IN2(n915), .IN3(\i_m4stg_frac/n1007 ), .QN(
        n6644) );
  NAND3X1 U717 ( .IN1(n1117), .IN2(n924), .IN3(\i_m4stg_frac/n672 ), .QN(n3582) );
  NAND3X1 U718 ( .IN1(\i_m4stg_frac/n669 ), .IN2(n1142), .IN3(
        \i_m4stg_frac/n671 ), .QN(n3594) );
  NAND3X1 U719 ( .IN1(n1144), .IN2(n950), .IN3(\i_m4stg_frac/n1013 ), .QN(
        n6325) );
  NAND3X1 U720 ( .IN1(n1145), .IN2(n951), .IN3(\i_m4stg_frac/n1004 ), .QN(
        n6598) );
  NAND3X1 U721 ( .IN1(n1143), .IN2(n949), .IN3(\i_m4stg_frac/n660 ), .QN(n3845) );
  NAND2X1 U722 ( .IN1(\i_m4stg_frac/n665 ), .IN2(n3630), .QN(n3647) );
  NAND2X1 U723 ( .IN1(\i_m4stg_frac/n1009 ), .IN2(n6377), .QN(n6395) );
  NAND2X1 U724 ( .IN1(n6362), .IN2(\i_m4stg_frac/n1001 ), .QN(n6567) );
  NAND2X1 U725 ( .IN1(\i_m4stg_frac/n674 ), .IN2(n3721), .QN(n3579) );
  NAND2X1 U726 ( .IN1(\i_m4stg_frac/n1010 ), .IN2(n6351), .QN(n6315) );
  NAND2X1 U727 ( .IN1(\i_m4stg_frac/n666 ), .IN2(n3606), .QN(n3570) );
  NAND2X1 U728 ( .IN1(n3506), .IN2(\i_m4stg_frac/n677 ), .QN(n3585) );
  NAND2X1 U729 ( .IN1(\i_m4stg_frac/n659 ), .IN2(n3312), .QN(n3817) );
  NAND2X1 U730 ( .IN1(n6362), .IN2(n1038), .QN(n6566) );
  NAND2X1 U731 ( .IN1(n3602), .IN2(\i_m4stg_frac/n668 ), .QN(n3569) );
  NAND2X1 U732 ( .IN1(n6347), .IN2(\i_m4stg_frac/n1012 ), .QN(n6314) );
  INVX2 U733 ( .INP(n6570), .ZN(n6330) );
  INVX2 U734 ( .INP(n7109), .ZN(n6336) );
  INVX2 U735 ( .INP(n6694), .ZN(n6326) );
  INVX2 U736 ( .INP(n3687), .ZN(n3591) );
  INVX2 U737 ( .INP(n5944), .ZN(n3844) );
  INVX2 U738 ( .INP(n8702), .ZN(n6597) );
  INVX2 U739 ( .INP(n7100), .ZN(n6338) );
  INVX2 U740 ( .INP(n6434), .ZN(n6324) );
  INVX2 U741 ( .INP(n5978), .ZN(n3868) );
  INVX2 U742 ( .INP(n8737), .ZN(n6621) );
  INVX2 U743 ( .INP(n3942), .ZN(n3593) );
  NAND3X1 U744 ( .IN1(\i_m4stg_frac/n663 ), .IN2(n1116), .IN3(
        \i_m4stg_frac/n665 ), .QN(n3550) );
  NAND3X1 U745 ( .IN1(\i_m4stg_frac/n1007 ), .IN2(n1118), .IN3(
        \i_m4stg_frac/n1009 ), .QN(n6294) );
  NAND3X1 U746 ( .IN1(\i_m4stg_frac/n672 ), .IN2(n1117), .IN3(
        \i_m4stg_frac/n674 ), .QN(n3580) );
  NAND3X1 U747 ( .IN1(n1142), .IN2(n948), .IN3(\i_m4stg_frac/n669 ), .QN(n3592) );
  NAND3X1 U748 ( .IN1(\i_m4stg_frac/n660 ), .IN2(n1143), .IN3(
        \i_m4stg_frac/n662 ), .QN(n3869) );
  NAND3X1 U749 ( .IN1(\i_m4stg_frac/n1004 ), .IN2(n1145), .IN3(
        \i_m4stg_frac/n1006 ), .QN(n6622) );
  NAND3X1 U750 ( .IN1(n933), .IN2(n1135), .IN3(\i_m4stg_frac/n1016 ), .QN(
        n6339) );
  NAND3X1 U751 ( .IN1(\i_m4stg_frac/n1013 ), .IN2(n1144), .IN3(
        \i_m4stg_frac/n1015 ), .QN(n6327) );
  INVX2 U752 ( .INP(n9035), .ZN(n8851) );
  NAND2X1 U753 ( .IN1(n3309), .IN2(n1123), .QN(n3741) );
  NOR2X0 U754 ( .IN1(\i_m4stg_frac/n655 ), .IN2(\i_m4stg_frac/n654 ), .QN(
        n3309) );
  NAND2X1 U755 ( .IN1(n6054), .IN2(n1196), .QN(n6491) );
  NAND2X1 U756 ( .IN1(\i_m4stg_frac/n656 ), .IN2(n3309), .QN(n3609) );
  NAND2X1 U757 ( .IN1(n6541), .IN2(\i_m4stg_frac/n1001 ), .QN(n6565) );
  NAND2X1 U758 ( .IN1(n6377), .IN2(n915), .QN(n6643) );
  NAND2X1 U759 ( .IN1(n3721), .IN2(n924), .QN(n3581) );
  NAND2X1 U760 ( .IN1(n3630), .IN2(n914), .QN(n3890) );
  NAND2X1 U761 ( .IN1(\i_m4stg_frac/n675 ), .IN2(n3820), .QN(n3588) );
  NAND2X1 U762 ( .IN1(n3614), .IN2(\i_m4stg_frac/n657 ), .QN(n3782) );
  NAND2X1 U763 ( .IN1(n8619), .IN2(\i_m4stg_frac/n998 ), .QN(n6493) );
  NAND2X1 U764 ( .IN1(n3670), .IN2(\i_m4stg_frac/n666 ), .QN(n3568) );
  NAND2X1 U765 ( .IN1(n6418), .IN2(\i_m4stg_frac/n1010 ), .QN(n6313) );
  NAND2X1 U766 ( .IN1(n6569), .IN2(\i_m4stg_frac/n1019 ), .QN(n6333) );
  INVX0 U767 ( .INP(n1610), .ZN(n1593) );
  INVX0 U768 ( .INP(n1610), .ZN(n1592) );
  INVX0 U769 ( .INP(n1609), .ZN(n1598) );
  INVX0 U770 ( .INP(n1609), .ZN(n1599) );
  INVX0 U771 ( .INP(n1609), .ZN(n1606) );
  INVX0 U772 ( .INP(n1609), .ZN(n1607) );
  INVX0 U773 ( .INP(n1609), .ZN(n1600) );
  INVX0 U774 ( .INP(n1609), .ZN(n1604) );
  INVX0 U775 ( .INP(n1609), .ZN(n1601) );
  INVX0 U776 ( .INP(n1609), .ZN(n1602) );
  INVX0 U777 ( .INP(n1609), .ZN(n1605) );
  INVX0 U778 ( .INP(n1609), .ZN(n1603) );
  INVX0 U779 ( .INP(n1610), .ZN(n1594) );
  INVX0 U780 ( .INP(n1610), .ZN(n1595) );
  INVX0 U781 ( .INP(n1610), .ZN(n1596) );
  INVX0 U782 ( .INP(n1610), .ZN(n1597) );
  INVX0 U783 ( .INP(n1609), .ZN(n1608) );
  INVX0 U784 ( .INP(n1409), .ZN(n1408) );
  INVX0 U785 ( .INP(n1409), .ZN(n1407) );
  INVX0 U786 ( .INP(n1409), .ZN(n1406) );
  INVX0 U787 ( .INP(n1410), .ZN(n1386) );
  INVX0 U788 ( .INP(n1410), .ZN(n1384) );
  INVX0 U789 ( .INP(n1409), .ZN(n1385) );
  INVX0 U790 ( .INP(n1410), .ZN(n1383) );
  INVX0 U791 ( .INP(n1410), .ZN(n1387) );
  INVX0 U792 ( .INP(n1410), .ZN(n1388) );
  INVX0 U793 ( .INP(n1410), .ZN(n1389) );
  INVX0 U794 ( .INP(n1409), .ZN(n1401) );
  INVX0 U795 ( .INP(n1409), .ZN(n1402) );
  INVX0 U796 ( .INP(n1410), .ZN(n1390) );
  INVX0 U797 ( .INP(n1409), .ZN(n1399) );
  INVX0 U798 ( .INP(n1409), .ZN(n1398) );
  INVX0 U799 ( .INP(n1409), .ZN(n1403) );
  INVX0 U800 ( .INP(n1409), .ZN(n1400) );
  INVX0 U801 ( .INP(n1410), .ZN(n1397) );
  INVX0 U802 ( .INP(n1410), .ZN(n1396) );
  INVX0 U803 ( .INP(n1410), .ZN(n1395) );
  INVX0 U804 ( .INP(n1410), .ZN(n1394) );
  INVX0 U805 ( .INP(n1410), .ZN(n1393) );
  INVX0 U806 ( .INP(n1410), .ZN(n1391) );
  INVX0 U807 ( .INP(n1410), .ZN(n1392) );
  INVX0 U808 ( .INP(n1409), .ZN(n1404) );
  INVX0 U809 ( .INP(n1409), .ZN(n1405) );
  INVX0 U810 ( .INP(n1508), .ZN(n1487) );
  INVX0 U811 ( .INP(n1507), .ZN(n1504) );
  INVX0 U812 ( .INP(n1507), .ZN(n1505) );
  INVX0 U813 ( .INP(n1508), .ZN(n1484) );
  INVX0 U814 ( .INP(n1508), .ZN(n1485) );
  INVX0 U815 ( .INP(n1508), .ZN(n1491) );
  INVX0 U816 ( .INP(n1508), .ZN(n1492) );
  INVX0 U817 ( .INP(n1508), .ZN(n1494) );
  INVX0 U818 ( .INP(n1507), .ZN(n1495) );
  INVX0 U819 ( .INP(n1507), .ZN(n1497) );
  INVX0 U820 ( .INP(n1507), .ZN(n1498) );
  INVX0 U821 ( .INP(n1508), .ZN(n1493) );
  INVX0 U822 ( .INP(n1507), .ZN(n1496) );
  INVX0 U823 ( .INP(n1507), .ZN(n1503) );
  INVX0 U824 ( .INP(n1507), .ZN(n1502) );
  INVX0 U825 ( .INP(n1507), .ZN(n1501) );
  INVX0 U826 ( .INP(n1508), .ZN(n1486) );
  INVX0 U827 ( .INP(n1507), .ZN(n1499) );
  INVX0 U828 ( .INP(n1507), .ZN(n1500) );
  INVX0 U829 ( .INP(n1508), .ZN(n1489) );
  INVX0 U830 ( .INP(n1508), .ZN(n1488) );
  INVX0 U831 ( .INP(n1508), .ZN(n1490) );
  INVX0 U832 ( .INP(n1508), .ZN(n1483) );
  INVX0 U833 ( .INP(n1509), .ZN(n1475) );
  INVX0 U834 ( .INP(n1509), .ZN(n1476) );
  INVX0 U835 ( .INP(n1509), .ZN(n1478) );
  INVX0 U836 ( .INP(n1510), .ZN(n1463) );
  INVX0 U837 ( .INP(n1510), .ZN(n1464) );
  INVX0 U838 ( .INP(n1510), .ZN(n1465) );
  INVX0 U839 ( .INP(n1510), .ZN(n1467) );
  INVX0 U840 ( .INP(n1510), .ZN(n1468) );
  INVX0 U841 ( .INP(n1510), .ZN(n1469) );
  INVX0 U842 ( .INP(n1510), .ZN(n1470) );
  INVX0 U843 ( .INP(n1509), .ZN(n1471) );
  INVX0 U844 ( .INP(n1509), .ZN(n1479) );
  INVX0 U845 ( .INP(n1510), .ZN(n1466) );
  INVX0 U846 ( .INP(n1509), .ZN(n1474) );
  INVX0 U847 ( .INP(n1509), .ZN(n1472) );
  INVX0 U848 ( .INP(n1509), .ZN(n1477) );
  INVX0 U849 ( .INP(n1510), .ZN(n1459) );
  INVX0 U850 ( .INP(n1509), .ZN(n1473) );
  INVX0 U851 ( .INP(n1509), .ZN(n1481) );
  INVX0 U852 ( .INP(n1509), .ZN(n1480) );
  INVX0 U853 ( .INP(n1509), .ZN(n1482) );
  INVX0 U854 ( .INP(n1510), .ZN(n1461) );
  INVX0 U855 ( .INP(n1510), .ZN(n1462) );
  INVX0 U856 ( .INP(n1510), .ZN(n1460) );
  INVX0 U857 ( .INP(n1511), .ZN(n1448) );
  INVX0 U858 ( .INP(n1511), .ZN(n1449) );
  INVX0 U859 ( .INP(n1511), .ZN(n1453) );
  INVX0 U860 ( .INP(n1511), .ZN(n1454) );
  INVX0 U861 ( .INP(n1511), .ZN(n1455) );
  INVX0 U862 ( .INP(n1511), .ZN(n1456) );
  INVX0 U863 ( .INP(n1511), .ZN(n1457) );
  INVX0 U864 ( .INP(n1511), .ZN(n1458) );
  INVX0 U865 ( .INP(n1511), .ZN(n1452) );
  INVX0 U866 ( .INP(n1511), .ZN(n1450) );
  INVX0 U867 ( .INP(n1511), .ZN(n1451) );
  INVX0 U868 ( .INP(n1507), .ZN(n1506) );
  INVX0 U869 ( .INP(n1631), .ZN(n1410) );
  INVX0 U870 ( .INP(n1631), .ZN(n1409) );
  INVX0 U871 ( .INP(n604), .ZN(n1609) );
  INVX0 U872 ( .INP(n604), .ZN(n1610) );
  INVX0 U873 ( .INP(n9307), .ZN(n1439) );
  INVX0 U874 ( .INP(n9307), .ZN(n1446) );
  INVX0 U875 ( .INP(n9307), .ZN(n1440) );
  INVX0 U876 ( .INP(n9307), .ZN(n1441) );
  INVX0 U877 ( .INP(n9307), .ZN(n1442) );
  INVX0 U878 ( .INP(n9307), .ZN(n1444) );
  INVX0 U879 ( .INP(n9307), .ZN(n1443) );
  INVX0 U880 ( .INP(n9307), .ZN(n1445) );
  INVX0 U881 ( .INP(n9675), .ZN(n1432) );
  INVX0 U882 ( .INP(n9675), .ZN(n1431) );
  INVX0 U883 ( .INP(n1555), .ZN(n1526) );
  INVX0 U884 ( .INP(n1555), .ZN(n1524) );
  INVX0 U885 ( .INP(n1554), .ZN(n1535) );
  INVX0 U886 ( .INP(n1554), .ZN(n1536) );
  INVX0 U887 ( .INP(n1553), .ZN(n1542) );
  INVX0 U888 ( .INP(n1554), .ZN(n1538) );
  INVX0 U889 ( .INP(n1554), .ZN(n1539) );
  INVX0 U890 ( .INP(n1554), .ZN(n1540) );
  INVX0 U891 ( .INP(n1554), .ZN(n1541) );
  INVX0 U892 ( .INP(n1555), .ZN(n1523) );
  INVX0 U893 ( .INP(n1555), .ZN(n1528) );
  INVX0 U894 ( .INP(n1555), .ZN(n1527) );
  INVX0 U895 ( .INP(n1554), .ZN(n1531) );
  INVX0 U896 ( .INP(n1555), .ZN(n1518) );
  INVX0 U897 ( .INP(n1555), .ZN(n1519) );
  INVX0 U898 ( .INP(n1555), .ZN(n1520) );
  INVX0 U899 ( .INP(n1555), .ZN(n1521) );
  INVX0 U900 ( .INP(n1554), .ZN(n1537) );
  INVX0 U901 ( .INP(n1555), .ZN(n1522) );
  INVX0 U902 ( .INP(n1553), .ZN(n1545) );
  INVX0 U903 ( .INP(n1553), .ZN(n1546) );
  INVX0 U904 ( .INP(n1553), .ZN(n1547) );
  INVX0 U905 ( .INP(n1553), .ZN(n1548) );
  INVX0 U906 ( .INP(n1553), .ZN(n1549) );
  INVX0 U907 ( .INP(n1553), .ZN(n1550) );
  INVX0 U908 ( .INP(n1553), .ZN(n1551) );
  INVX0 U909 ( .INP(n1553), .ZN(n1552) );
  INVX0 U910 ( .INP(n1553), .ZN(n1543) );
  INVX0 U911 ( .INP(n1553), .ZN(n1544) );
  INVX0 U912 ( .INP(n1554), .ZN(n1532) );
  INVX0 U913 ( .INP(n1554), .ZN(n1533) );
  INVX0 U914 ( .INP(n1554), .ZN(n1534) );
  INVX0 U915 ( .INP(n1555), .ZN(n1529) );
  INVX0 U916 ( .INP(n1554), .ZN(n1530) );
  INVX0 U917 ( .INP(n1555), .ZN(n1525) );
  INVX0 U918 ( .INP(n9661), .ZN(n1430) );
  INVX0 U919 ( .INP(n1556), .ZN(n1512) );
  INVX0 U920 ( .INP(n1556), .ZN(n1513) );
  INVX0 U921 ( .INP(n1556), .ZN(n1514) );
  INVX0 U922 ( .INP(n1556), .ZN(n1515) );
  INVX0 U923 ( .INP(n1556), .ZN(n1516) );
  INVX0 U924 ( .INP(n1556), .ZN(n1517) );
  INVX0 U925 ( .INP(n9675), .ZN(n1437) );
  INVX0 U926 ( .INP(n9675), .ZN(n1438) );
  INVX0 U927 ( .INP(n9675), .ZN(n1433) );
  INVX0 U928 ( .INP(n9675), .ZN(n1436) );
  INVX0 U929 ( .INP(n9675), .ZN(n1434) );
  INVX0 U930 ( .INP(n9675), .ZN(n1435) );
  INVX0 U931 ( .INP(n9661), .ZN(n1427) );
  INVX0 U932 ( .INP(n9661), .ZN(n1423) );
  INVX0 U933 ( .INP(n9661), .ZN(n1425) );
  INVX0 U934 ( .INP(n9661), .ZN(n1429) );
  INVX0 U935 ( .INP(n9661), .ZN(n1428) );
  INVX0 U936 ( .INP(n9661), .ZN(n1426) );
  INVX0 U937 ( .INP(n9661), .ZN(n1421) );
  INVX0 U938 ( .INP(n9661), .ZN(n1424) );
  INVX0 U939 ( .INP(n9661), .ZN(n1422) );
  INVX0 U940 ( .INP(n9307), .ZN(n1447) );
  INVX0 U941 ( .INP(n1589), .ZN(n1581) );
  INVX0 U942 ( .INP(n1589), .ZN(n1582) );
  INVX0 U943 ( .INP(n1589), .ZN(n1583) );
  INVX0 U944 ( .INP(n1589), .ZN(n1584) );
  INVX0 U945 ( .INP(n1589), .ZN(n1585) );
  INVX0 U946 ( .INP(n1589), .ZN(n1586) );
  INVX0 U947 ( .INP(n1589), .ZN(n1587) );
  INVX0 U948 ( .INP(n1589), .ZN(n1580) );
  INVX0 U949 ( .INP(n1589), .ZN(n1579) );
  INVX0 U950 ( .INP(n1590), .ZN(n1576) );
  INVX0 U951 ( .INP(n1590), .ZN(n1575) );
  INVX0 U952 ( .INP(n1590), .ZN(n1574) );
  INVX0 U953 ( .INP(n1589), .ZN(n1577) );
  INVX0 U954 ( .INP(n1590), .ZN(n1569) );
  INVX0 U955 ( .INP(n1590), .ZN(n1566) );
  INVX0 U956 ( .INP(n1590), .ZN(n1568) );
  INVX0 U957 ( .INP(n1590), .ZN(n1565) );
  INVX0 U958 ( .INP(n1590), .ZN(n1572) );
  INVX0 U959 ( .INP(n1590), .ZN(n1570) );
  INVX0 U960 ( .INP(n1590), .ZN(n1567) );
  INVX0 U961 ( .INP(n1590), .ZN(n1571) );
  INVX0 U962 ( .INP(n1589), .ZN(n1578) );
  INVX0 U963 ( .INP(n1590), .ZN(n1573) );
  INVX0 U964 ( .INP(n1591), .ZN(n1561) );
  INVX0 U965 ( .INP(n1591), .ZN(n1562) );
  INVX0 U966 ( .INP(n1591), .ZN(n1563) );
  INVX0 U967 ( .INP(n1591), .ZN(n1564) );
  INVX0 U968 ( .INP(n1591), .ZN(n1558) );
  INVX0 U969 ( .INP(n1591), .ZN(n1557) );
  INVX0 U970 ( .INP(n1591), .ZN(n1559) );
  INVX0 U971 ( .INP(n1591), .ZN(n1560) );
  INVX0 U972 ( .INP(n1589), .ZN(n1588) );
  NBUFFX2 U973 ( .INP(n911), .Z(n1507) );
  NBUFFX2 U974 ( .INP(n911), .Z(n1508) );
  NBUFFX2 U975 ( .INP(n911), .Z(n1509) );
  NBUFFX2 U976 ( .INP(n911), .Z(n1510) );
  NBUFFX2 U977 ( .INP(n911), .Z(n1511) );
  INVX0 U978 ( .INP(n1382), .ZN(n1411) );
  INVX0 U979 ( .INP(n1382), .ZN(n1417) );
  INVX0 U980 ( .INP(n1382), .ZN(n1412) );
  INVX0 U981 ( .INP(n1382), .ZN(n1418) );
  INVX0 U982 ( .INP(n1382), .ZN(n1415) );
  INVX0 U983 ( .INP(n1382), .ZN(n1416) );
  INVX0 U984 ( .INP(n1382), .ZN(n1413) );
  INVX0 U985 ( .INP(n1382), .ZN(n1414) );
  INVX0 U986 ( .INP(n1382), .ZN(n1419) );
  INVX0 U987 ( .INP(n1381), .ZN(n1618) );
  INVX0 U988 ( .INP(n1381), .ZN(n1617) );
  INVX0 U989 ( .INP(n1381), .ZN(n1619) );
  INVX0 U990 ( .INP(n1381), .ZN(n1620) );
  INVX0 U991 ( .INP(n1381), .ZN(n1616) );
  INVX0 U992 ( .INP(n1381), .ZN(n1621) );
  INVX0 U993 ( .INP(n1381), .ZN(n1615) );
  INVX0 U994 ( .INP(n1381), .ZN(n1611) );
  INVX0 U995 ( .INP(n1381), .ZN(n1614) );
  INVX0 U996 ( .INP(n1381), .ZN(n1612) );
  INVX0 U997 ( .INP(n1381), .ZN(n1613) );
  INVX0 U998 ( .INP(n1382), .ZN(n1420) );
  INVX0 U999 ( .INP(n1381), .ZN(n1622) );
  INVX0 U1000 ( .INP(\fpu_mul_frac_dp/n832 ), .ZN(n1589) );
  INVX0 U1001 ( .INP(\fpu_mul_frac_dp/n832 ), .ZN(n1590) );
  INVX0 U1002 ( .INP(\i_m4stg_frac/n854 ), .ZN(n1553) );
  INVX0 U1003 ( .INP(\i_m4stg_frac/n854 ), .ZN(n1554) );
  INVX0 U1004 ( .INP(\i_m4stg_frac/n854 ), .ZN(n1555) );
  INVX0 U1005 ( .INP(\fpu_mul_frac_dp/n832 ), .ZN(n1591) );
  INVX0 U1006 ( .INP(\i_m4stg_frac/n854 ), .ZN(n1556) );
  OR2X1 U1007 ( .IN1(n189), .IN2(n709), .Q(n1381) );
  OR2X1 U1008 ( .IN1(\fpu_mul_frac_dp/n831 ), .IN2(\fpu_mul_frac_dp/n834 ), 
        .Q(n1382) );
  OA221X1 U1009 ( .IN1(n1623), .IN2(n1624), .IN3(n449), .IN4(n1625), .IN5(
        n1626), .Q(n94) );
  XOR3X1 U1010 ( .IN1(n1627), .IN2(n1628), .IN3(n1629), .Q(n1623) );
  NOR2X0 U1011 ( .IN1(n443), .IN2(n1630), .QN(n456) );
  AO22X1 U1012 ( .IN1(inq_in2[62]), .IN2(n1602), .IN3(n1395), .IN4(n1194), .Q(
        n371) );
  AO22X1 U1013 ( .IN1(inq_in2[61]), .IN2(n1602), .IN3(n1387), .IN4(n1179), .Q(
        n370) );
  AO22X1 U1014 ( .IN1(inq_in2[60]), .IN2(n1602), .IN3(n1395), .IN4(n1176), .Q(
        n369) );
  AO22X1 U1015 ( .IN1(inq_in2[59]), .IN2(n1602), .IN3(n1395), .IN4(n975), .Q(
        n368) );
  AO22X1 U1016 ( .IN1(inq_in2[58]), .IN2(n1602), .IN3(n1395), .IN4(n902), .Q(
        n367) );
  AO22X1 U1017 ( .IN1(inq_in2[57]), .IN2(n1602), .IN3(n1395), .IN4(n961), .Q(
        n366) );
  AO22X1 U1018 ( .IN1(inq_in2[56]), .IN2(n1602), .IN3(n1395), .IN4(n905), .Q(
        n365) );
  AO22X1 U1019 ( .IN1(inq_in2[55]), .IN2(n1602), .IN3(n1394), .IN4(n964), .Q(
        n364) );
  AO21X1 U1020 ( .IN1(n1386), .IN2(n1231), .IN3(n1632), .Q(n363) );
  AO22X1 U1021 ( .IN1(inq_in2[53]), .IN2(n1602), .IN3(n1394), .IN4(n1228), .Q(
        n362) );
  AO22X1 U1022 ( .IN1(inq_in2[52]), .IN2(n1603), .IN3(n1394), .IN4(n1227), .Q(
        n361) );
  AO22X1 U1023 ( .IN1(inq_in1[62]), .IN2(n1603), .IN3(n1394), .IN4(n1178), .Q(
        n360) );
  AO22X1 U1024 ( .IN1(inq_in1[61]), .IN2(n1603), .IN3(n1394), .IN4(n1175), .Q(
        n359) );
  AO22X1 U1025 ( .IN1(inq_in1[60]), .IN2(n1603), .IN3(n1394), .IN4(n1177), .Q(
        n358) );
  AO22X1 U1026 ( .IN1(inq_in1[59]), .IN2(n1603), .IN3(n1394), .IN4(n965), .Q(
        n357) );
  AO22X1 U1027 ( .IN1(inq_in1[58]), .IN2(n1605), .IN3(n1394), .IN4(n903), .Q(
        n356) );
  AO22X1 U1028 ( .IN1(inq_in1[57]), .IN2(n1603), .IN3(n1394), .IN4(n962), .Q(
        n355) );
  AO22X1 U1029 ( .IN1(inq_in1[56]), .IN2(n1603), .IN3(n1394), .IN4(n904), .Q(
        n354) );
  AO22X1 U1030 ( .IN1(inq_in1[55]), .IN2(n1603), .IN3(n1394), .IN4(n963), .Q(
        n353) );
  AO21X1 U1031 ( .IN1(n1386), .IN2(n1232), .IN3(n1633), .Q(n352) );
  AO22X1 U1032 ( .IN1(inq_in1[53]), .IN2(n1603), .IN3(n1394), .IN4(n1225), .Q(
        n351) );
  AO22X1 U1033 ( .IN1(inq_in1[52]), .IN2(n1603), .IN3(n1394), .IN4(n1226), .Q(
        n350) );
  AO221X1 U1034 ( .IN1(n1634), .IN2(n1635), .IN3(n1385), .IN4(n994), .IN5(
        n1636), .Q(n349) );
  AO21X1 U1035 ( .IN1(n1637), .IN2(n1638), .IN3(n1639), .Q(n1635) );
  AO221X1 U1036 ( .IN1(n1640), .IN2(n1634), .IN3(n1385), .IN4(n989), .IN5(
        n1636), .Q(n348) );
  XOR3X1 U1037 ( .IN1(n1641), .IN2(n1642), .IN3(n1643), .Q(n1640) );
  AO221X1 U1038 ( .IN1(n1644), .IN2(n1634), .IN3(n1385), .IN4(n990), .IN5(
        n1636), .Q(n347) );
  XOR3X1 U1039 ( .IN1(n1645), .IN2(n1646), .IN3(n1647), .Q(n1644) );
  AO221X1 U1040 ( .IN1(n1648), .IN2(n1634), .IN3(n1385), .IN4(n995), .IN5(
        n1636), .Q(n346) );
  XOR3X1 U1041 ( .IN1(n1649), .IN2(n1650), .IN3(n1651), .Q(n1648) );
  AO221X1 U1042 ( .IN1(n1652), .IN2(n1634), .IN3(n1385), .IN4(n991), .IN5(
        n1636), .Q(n345) );
  XOR3X1 U1043 ( .IN1(n1653), .IN2(n1654), .IN3(n1655), .Q(n1652) );
  AO221X1 U1044 ( .IN1(n1656), .IN2(n1634), .IN3(n1385), .IN4(n992), .IN5(
        n1636), .Q(n344) );
  XOR3X1 U1045 ( .IN1(n1657), .IN2(n1658), .IN3(n1659), .Q(n1656) );
  AO221X1 U1046 ( .IN1(n1660), .IN2(n1634), .IN3(n1385), .IN4(n993), .IN5(
        n1636), .Q(n343) );
  NAND2X0 U1047 ( .IN1(n1626), .IN2(n1661), .QN(n1636) );
  XOR3X1 U1048 ( .IN1(n1662), .IN2(n1663), .IN3(n1664), .Q(n1660) );
  AO221X1 U1049 ( .IN1(n1665), .IN2(n1634), .IN3(n1385), .IN4(n1140), .IN5(
        n1666), .Q(n342) );
  NAND2X0 U1050 ( .IN1(n1626), .IN2(n1667), .QN(n1666) );
  XOR3X1 U1051 ( .IN1(n1668), .IN2(n1669), .IN3(n1670), .Q(n1665) );
  AO221X1 U1052 ( .IN1(n1634), .IN2(n1671), .IN3(n1385), .IN4(n1210), .IN5(
        n1672), .Q(n341) );
  INVX0 U1053 ( .INP(n1626), .ZN(n1672) );
  XNOR3X1 U1054 ( .IN1(n1673), .IN2(n1674), .IN3(n1675), .Q(n1671) );
  AO221X1 U1055 ( .IN1(n1634), .IN2(n1676), .IN3(n876), .IN4(n1383), .IN5(
        n1677), .Q(n340) );
  NAND2X0 U1056 ( .IN1(n1678), .IN2(n1667), .QN(n1677) );
  OR2X1 U1057 ( .IN1(n1661), .IN2(\fpu_mul_ctl/n257 ), .Q(n1667) );
  NAND3X0 U1058 ( .IN1(n1592), .IN2(n1679), .IN3(n1680), .QN(n1661) );
  XNOR2X1 U1059 ( .IN1(n1681), .IN2(n1682), .Q(n1676) );
  OA21X1 U1060 ( .IN1(n1683), .IN2(n1684), .IN3(n1685), .Q(n1682) );
  INVX0 U1061 ( .INP(n1624), .ZN(n1634) );
  NAND3X0 U1062 ( .IN1(n1678), .IN2(n1626), .IN3(n1686), .QN(n339) );
  OA22X1 U1063 ( .IN1(n1687), .IN2(n1624), .IN3(n1625), .IN4(n1277), .Q(n1686)
         );
  NAND2X0 U1064 ( .IN1(n1688), .IN2(n1689), .QN(n1624) );
  OA22X1 U1065 ( .IN1(n1690), .IN2(n1681), .IN3(n1683), .IN4(n1684), .Q(n1687)
         );
  NAND2X0 U1066 ( .IN1(m1stg_dblop), .IN2(n1178), .QN(n1681) );
  INVX0 U1067 ( .INP(n1685), .ZN(n1690) );
  NAND2X0 U1068 ( .IN1(n1684), .IN2(n1683), .QN(n1685) );
  AO22X1 U1069 ( .IN1(n1674), .IN2(n1675), .IN3(n1691), .IN4(n1673), .Q(n1683)
         );
  NAND2X0 U1070 ( .IN1(m1stg_dblop), .IN2(n1175), .QN(n1673) );
  OR2X1 U1071 ( .IN1(n1674), .IN2(n1675), .Q(n1691) );
  AO22X1 U1072 ( .IN1(n1629), .IN2(n1628), .IN3(n1692), .IN4(n1627), .Q(n1675)
         );
  NAND2X0 U1073 ( .IN1(m1stg_dblop), .IN2(n1177), .QN(n1627) );
  OR2X1 U1074 ( .IN1(n1629), .IN2(n1628), .Q(n1692) );
  NAND2X0 U1075 ( .IN1(m1stg_dblop), .IN2(n1176), .QN(n1628) );
  AO22X1 U1076 ( .IN1(n1669), .IN2(n1693), .IN3(n1668), .IN4(n1694), .Q(n1629)
         );
  NAND2X0 U1077 ( .IN1(n1695), .IN2(n1670), .QN(n1694) );
  AOI22X1 U1078 ( .IN1(m1stg_sngop), .IN2(n1194), .IN3(m1stg_dblop), .IN4(n975), .QN(n1668) );
  INVX0 U1079 ( .INP(n1670), .ZN(n1693) );
  AO22X1 U1080 ( .IN1(n1664), .IN2(n1663), .IN3(n1696), .IN4(n1662), .Q(n1670)
         );
  AO22X1 U1081 ( .IN1(m1stg_sngop), .IN2(n1179), .IN3(m1stg_dblop), .IN4(n902), 
        .Q(n1662) );
  OR2X1 U1082 ( .IN1(n1663), .IN2(n1664), .Q(n1696) );
  AO22X1 U1083 ( .IN1(m1stg_sngop), .IN2(n1175), .IN3(m1stg_dblop), .IN4(n903), 
        .Q(n1663) );
  AO22X1 U1084 ( .IN1(n1659), .IN2(n1658), .IN3(n1697), .IN4(n1657), .Q(n1664)
         );
  AO22X1 U1085 ( .IN1(m1stg_sngop), .IN2(n1176), .IN3(m1stg_dblop), .IN4(n961), 
        .Q(n1657) );
  OR2X1 U1086 ( .IN1(n1658), .IN2(n1659), .Q(n1697) );
  AO22X1 U1087 ( .IN1(m1stg_sngop), .IN2(n1177), .IN3(m1stg_dblop), .IN4(n962), 
        .Q(n1658) );
  AO22X1 U1088 ( .IN1(n1655), .IN2(n1654), .IN3(n1698), .IN4(n1653), .Q(n1659)
         );
  AO22X1 U1089 ( .IN1(m1stg_sngop), .IN2(n975), .IN3(m1stg_dblop), .IN4(n905), 
        .Q(n1653) );
  OR2X1 U1090 ( .IN1(n1654), .IN2(n1655), .Q(n1698) );
  AO22X1 U1091 ( .IN1(m1stg_sngop), .IN2(n965), .IN3(m1stg_dblop), .IN4(n904), 
        .Q(n1654) );
  AO22X1 U1092 ( .IN1(n1651), .IN2(n1650), .IN3(n1699), .IN4(n1649), .Q(n1655)
         );
  AO22X1 U1093 ( .IN1(m1stg_sngop), .IN2(n902), .IN3(m1stg_dblop), .IN4(n964), 
        .Q(n1649) );
  OR2X1 U1094 ( .IN1(n1650), .IN2(n1651), .Q(n1699) );
  AO22X1 U1095 ( .IN1(m1stg_sngop), .IN2(n903), .IN3(m1stg_dblop), .IN4(n963), 
        .Q(n1650) );
  AO22X1 U1096 ( .IN1(n1647), .IN2(n1646), .IN3(n1700), .IN4(n1645), .Q(n1651)
         );
  AO22X1 U1097 ( .IN1(m1stg_sngop), .IN2(n961), .IN3(m1stg_dblop), .IN4(n1231), 
        .Q(n1645) );
  OR2X1 U1098 ( .IN1(n1646), .IN2(n1647), .Q(n1700) );
  AO22X1 U1099 ( .IN1(m1stg_sngop), .IN2(n962), .IN3(m1stg_dblop), .IN4(n1232), 
        .Q(n1646) );
  AO22X1 U1100 ( .IN1(n1641), .IN2(n1642), .IN3(n1701), .IN4(n1643), .Q(n1647)
         );
  AO22X1 U1101 ( .IN1(m1stg_sngop), .IN2(n904), .IN3(m1stg_dblop), .IN4(n1225), 
        .Q(n1643) );
  OR2X1 U1102 ( .IN1(n1642), .IN2(n1641), .Q(n1701) );
  INVX0 U1103 ( .INP(n1639), .ZN(n1642) );
  NOR2X0 U1104 ( .IN1(n1638), .IN2(n1637), .QN(n1639) );
  AO22X1 U1105 ( .IN1(m1stg_sngop), .IN2(n963), .IN3(m1stg_dblop), .IN4(n1226), 
        .Q(n1637) );
  AO22X1 U1106 ( .IN1(m1stg_sngop), .IN2(n964), .IN3(m1stg_dblop), .IN4(n1227), 
        .Q(n1638) );
  AO22X1 U1107 ( .IN1(m1stg_sngop), .IN2(n905), .IN3(m1stg_dblop), .IN4(n1228), 
        .Q(n1641) );
  INVX0 U1108 ( .INP(n1695), .ZN(n1669) );
  AO22X1 U1109 ( .IN1(m1stg_sngop), .IN2(n1178), .IN3(m1stg_dblop), .IN4(n965), 
        .Q(n1695) );
  NAND2X0 U1110 ( .IN1(m1stg_dblop), .IN2(n1179), .QN(n1674) );
  NAND2X0 U1111 ( .IN1(m1stg_dblop), .IN2(n1194), .QN(n1684) );
  NAND3X0 U1112 ( .IN1(n1592), .IN2(n1679), .IN3(n1702), .QN(n1626) );
  OAI21X1 U1113 ( .IN1(n1625), .IN2(n17), .IN3(n1678), .QN(n338) );
  NAND4X0 U1114 ( .IN1(n1680), .IN2(n1689), .IN3(n1703), .IN4(n1055), .QN(
        n1678) );
  INVX0 U1115 ( .INP(n1688), .ZN(n1703) );
  AO22X1 U1116 ( .IN1(n1597), .IN2(n994), .IN3(n1394), .IN4(n1238), .Q(n337)
         );
  AO22X1 U1117 ( .IN1(n1597), .IN2(n989), .IN3(n1393), .IN4(n1233), .Q(n336)
         );
  AO22X1 U1118 ( .IN1(n1597), .IN2(n990), .IN3(n1393), .IN4(n1234), .Q(n335)
         );
  AO22X1 U1119 ( .IN1(n1597), .IN2(n995), .IN3(n1393), .IN4(n1239), .Q(n334)
         );
  AO22X1 U1120 ( .IN1(n1597), .IN2(n991), .IN3(n1393), .IN4(n1235), .Q(n333)
         );
  AO22X1 U1121 ( .IN1(n1597), .IN2(n992), .IN3(n1393), .IN4(n1236), .Q(n332)
         );
  AO22X1 U1122 ( .IN1(n1597), .IN2(n993), .IN3(n1393), .IN4(n1237), .Q(n331)
         );
  AO22X1 U1123 ( .IN1(n1631), .IN2(n1285), .IN3(n1704), .IN4(n1592), .Q(n330)
         );
  XOR2X1 U1124 ( .IN1(n1140), .IN2(m2stg_fmuls), .Q(n1704) );
  AO22X1 U1125 ( .IN1(n1404), .IN2(n1286), .IN3(n1705), .IN4(n1593), .Q(n329)
         );
  XNOR2X1 U1126 ( .IN1(n449), .IN2(n1706), .Q(n1705) );
  OA21X1 U1127 ( .IN1(n454), .IN2(n1218), .IN3(n1707), .Q(n1706) );
  AO22X1 U1128 ( .IN1(n1631), .IN2(n1348), .IN3(n1708), .IN4(n1593), .Q(n328)
         );
  XOR3X1 U1129 ( .IN1(n441), .IN2(n1709), .IN3(n1710), .Q(n1708) );
  AO22X1 U1130 ( .IN1(n1404), .IN2(n1287), .IN3(n1593), .IN4(n1711), .Q(n327)
         );
  XOR3X1 U1131 ( .IN1(n876), .IN2(n1712), .IN3(n1713), .Q(n1711) );
  AO22X1 U1132 ( .IN1(n1631), .IN2(n1349), .IN3(n1593), .IN4(n1714), .Q(n326)
         );
  XOR3X1 U1133 ( .IN1(n1715), .IN2(n878), .IN3(n1716), .Q(n1714) );
  AO22X1 U1134 ( .IN1(n1404), .IN2(n1288), .IN3(n1717), .IN4(n1593), .Q(n325)
         );
  XOR3X1 U1135 ( .IN1(n1718), .IN2(n17), .IN3(n1715), .Q(n1717) );
  OA22X1 U1136 ( .IN1(n1719), .IN2(n1277), .IN3(n1712), .IN4(n1720), .Q(n1718)
         );
  INVX0 U1137 ( .INP(n1716), .ZN(n1720) );
  NOR2X0 U1138 ( .IN1(n1715), .IN2(n1716), .QN(n1719) );
  AO22X1 U1139 ( .IN1(n1721), .IN2(n1715), .IN3(n876), .IN4(n1722), .Q(n1716)
         );
  NAND2X0 U1140 ( .IN1(n1713), .IN2(n1712), .QN(n1722) );
  INVX0 U1141 ( .INP(n1721), .ZN(n1713) );
  AO21X1 U1142 ( .IN1(n1707), .IN2(n1210), .IN3(n1710), .Q(n1721) );
  OAI22X1 U1143 ( .IN1(n1218), .IN2(n454), .IN3(n1709), .IN4(n449), .QN(n1710)
         );
  INVX0 U1144 ( .INP(n1709), .ZN(n1707) );
  NOR2X0 U1145 ( .IN1(m2stg_fmuls), .IN2(m2stg_fsmuld), .QN(n1709) );
  INVX0 U1146 ( .INP(n1712), .ZN(n1715) );
  NOR2X0 U1147 ( .IN1(m2stg_fmuld), .IN2(m2stg_fmuls), .QN(n1712) );
  AO22X1 U1148 ( .IN1(n1597), .IN2(n1238), .IN3(n1393), .IN4(n968), .Q(n324)
         );
  AO22X1 U1149 ( .IN1(n1597), .IN2(n1233), .IN3(n1393), .IN4(n998), .Q(n323)
         );
  AO22X1 U1150 ( .IN1(n1597), .IN2(n1234), .IN3(n1393), .IN4(n969), .Q(n322)
         );
  AO22X1 U1151 ( .IN1(n1597), .IN2(n1239), .IN3(n1393), .IN4(n1001), .Q(n321)
         );
  AO22X1 U1152 ( .IN1(n1597), .IN2(n1235), .IN3(n1393), .IN4(n970), .Q(n320)
         );
  AO22X1 U1153 ( .IN1(n1597), .IN2(n1236), .IN3(n1393), .IN4(n996), .Q(n319)
         );
  AO22X1 U1154 ( .IN1(n1597), .IN2(n1237), .IN3(n1393), .IN4(n971), .Q(n318)
         );
  AO22X1 U1155 ( .IN1(n1597), .IN2(n1285), .IN3(n1393), .IN4(n972), .Q(n317)
         );
  AO22X1 U1156 ( .IN1(n1597), .IN2(n1286), .IN3(n1392), .IN4(n999), .Q(n316)
         );
  OAI22X1 U1157 ( .IN1(n1723), .IN2(n137), .IN3(n1625), .IN4(n136), .QN(n315)
         );
  AO22X1 U1158 ( .IN1(n1597), .IN2(n1287), .IN3(n1392), .IN4(n997), .Q(n314)
         );
  OAI22X1 U1159 ( .IN1(n1723), .IN2(n145), .IN3(n1625), .IN4(n144), .QN(n313)
         );
  AO22X1 U1160 ( .IN1(n1597), .IN2(n1288), .IN3(n1392), .IN4(n1000), .Q(n312)
         );
  AO22X1 U1161 ( .IN1(n1596), .IN2(n968), .IN3(n1392), .IN4(n1154), .Q(n311)
         );
  OAI22X1 U1162 ( .IN1(n1723), .IN2(n104), .IN3(n1625), .IN4(n103), .QN(n310)
         );
  AO22X1 U1163 ( .IN1(n1596), .IN2(n969), .IN3(n1392), .IN4(n1212), .Q(n309)
         );
  AO22X1 U1164 ( .IN1(n1596), .IN2(n1001), .IN3(n1392), .IN4(n1214), .Q(n308)
         );
  AO22X1 U1165 ( .IN1(n1596), .IN2(n970), .IN3(n1392), .IN4(n1211), .Q(n307)
         );
  AO22X1 U1166 ( .IN1(n1596), .IN2(n996), .IN3(n1392), .IN4(n1213), .Q(n306)
         );
  AO22X1 U1167 ( .IN1(n1596), .IN2(n971), .IN3(n1392), .IN4(n1122), .Q(n305)
         );
  AO22X1 U1168 ( .IN1(n1596), .IN2(n972), .IN3(n1392), .IN4(n1153), .Q(n304)
         );
  OAI22X1 U1169 ( .IN1(n1723), .IN2(n132), .IN3(n1625), .IN4(n453), .QN(n303)
         );
  OAI22X1 U1170 ( .IN1(n1723), .IN2(n136), .IN3(n1625), .IN4(n135), .QN(n302)
         );
  AO22X1 U1171 ( .IN1(n1596), .IN2(n997), .IN3(n1392), .IN4(n1152), .Q(n301)
         );
  OAI22X1 U1172 ( .IN1(n1723), .IN2(n144), .IN3(n1625), .IN4(n143), .QN(n300)
         );
  OAI22X1 U1173 ( .IN1(n1723), .IN2(n148), .IN3(n1625), .IN4(n147), .QN(n299)
         );
  AO22X1 U1174 ( .IN1(n1596), .IN2(n968), .IN3(n1392), .IN4(n895), .Q(n298) );
  AO22X1 U1175 ( .IN1(n1596), .IN2(n998), .IN3(n1392), .IN4(n1115), .Q(n297)
         );
  AO22X1 U1176 ( .IN1(n1596), .IN2(n969), .IN3(n1392), .IN4(n1166), .Q(n296)
         );
  OAI22X1 U1177 ( .IN1(n1723), .IN2(n112), .IN3(n1625), .IN4(n110), .QN(n295)
         );
  AO22X1 U1178 ( .IN1(n1596), .IN2(n970), .IN3(n1391), .IN4(n888), .Q(n294) );
  OAI22X1 U1179 ( .IN1(n1723), .IN2(n120), .IN3(n1625), .IN4(n118), .QN(n293)
         );
  AO22X1 U1180 ( .IN1(n1596), .IN2(n971), .IN3(n1391), .IN4(n1114), .Q(n292)
         );
  AO22X1 U1181 ( .IN1(n1596), .IN2(n972), .IN3(n1391), .IN4(n900), .Q(n291) );
  AO22X1 U1182 ( .IN1(n1596), .IN2(n999), .IN3(n1391), .IN4(n1203), .Q(n290)
         );
  OAI22X1 U1183 ( .IN1(n1723), .IN2(n136), .IN3(n1625), .IN4(n134), .QN(n289)
         );
  OAI22X1 U1184 ( .IN1(n1723), .IN2(n140), .IN3(n1625), .IN4(n138), .QN(n288)
         );
  OAI22X1 U1185 ( .IN1(n1723), .IN2(n144), .IN3(n1625), .IN4(n142), .QN(n287)
         );
  AO22X1 U1186 ( .IN1(n1596), .IN2(n1000), .IN3(n1391), .IN4(n1119), .Q(n286)
         );
  AO22X1 U1187 ( .IN1(n1404), .IN2(m4stg_exp[0]), .IN3(n1724), .IN4(n1725), 
        .Q(n285) );
  AO21X1 U1188 ( .IN1(m3stg_ld0_inv[0]), .IN2(n1154), .IN3(n1726), .Q(n1725)
         );
  AO22X1 U1189 ( .IN1(n1404), .IN2(m4stg_exp[1]), .IN3(n1724), .IN4(n1727), 
        .Q(n284) );
  XOR3X1 U1190 ( .IN1(n103), .IN2(m3stg_ld0_inv[1]), .IN3(n1726), .Q(n1727) );
  AO22X1 U1191 ( .IN1(n1404), .IN2(m4stg_exp[2]), .IN3(n1724), .IN4(n1728), 
        .Q(n283) );
  XOR3X1 U1192 ( .IN1(n1150), .IN2(n107), .IN3(n1729), .Q(n1728) );
  AO22X1 U1193 ( .IN1(n1404), .IN2(m4stg_exp[3]), .IN3(n1724), .IN4(n1730), 
        .Q(n282) );
  XOR3X1 U1194 ( .IN1(n111), .IN2(m3stg_ld0_inv[3]), .IN3(n1731), .Q(n1730) );
  AO22X1 U1195 ( .IN1(n1404), .IN2(m4stg_exp[4]), .IN3(n1724), .IN4(n1732), 
        .Q(n281) );
  XOR3X1 U1196 ( .IN1(n1059), .IN2(n115), .IN3(n1733), .Q(n1732) );
  AO22X1 U1197 ( .IN1(n1404), .IN2(m4stg_exp[5]), .IN3(n1724), .IN4(n1734), 
        .Q(n280) );
  XOR3X1 U1198 ( .IN1(n119), .IN2(m3stg_ld0_inv[5]), .IN3(n1735), .Q(n1734) );
  AO22X1 U1199 ( .IN1(n1405), .IN2(m4stg_exp[6]), .IN3(n1724), .IN4(n1736), 
        .Q(n279) );
  XOR3X1 U1200 ( .IN1(m3stg_ld0_inv[6]), .IN2(n1122), .IN3(n1737), .Q(n1736)
         );
  AO22X1 U1201 ( .IN1(n1405), .IN2(m4stg_exp[7]), .IN3(n1724), .IN4(n1738), 
        .Q(n278) );
  AO21X1 U1202 ( .IN1(n1739), .IN2(n1153), .IN3(n1740), .Q(n1738) );
  AO22X1 U1203 ( .IN1(n1405), .IN2(m4stg_exp[8]), .IN3(n1724), .IN4(n1741), 
        .Q(n277) );
  OAI21X1 U1204 ( .IN1(n1740), .IN2(n453), .IN3(n1742), .QN(n1741) );
  AO22X1 U1205 ( .IN1(n1405), .IN2(m4stg_exp[9]), .IN3(n1724), .IN4(n1743), 
        .Q(n276) );
  OAI21X1 U1206 ( .IN1(n1744), .IN2(n135), .IN3(n1745), .QN(n1743) );
  AO22X1 U1207 ( .IN1(n1405), .IN2(m4stg_exp[10]), .IN3(n1724), .IN4(n1746), 
        .Q(n275) );
  AO21X1 U1208 ( .IN1(n1745), .IN2(n1152), .IN3(n1747), .Q(n1746) );
  AO22X1 U1209 ( .IN1(n1405), .IN2(m4stg_exp[11]), .IN3(n1748), .IN4(n1724), 
        .Q(n274) );
  AND2X1 U1210 ( .IN1(n1594), .IN2(n1749), .Q(n1724) );
  XNOR2X1 U1211 ( .IN1(n143), .IN2(n1747), .Q(n1748) );
  AO221X1 U1212 ( .IN1(n1750), .IN2(n1751), .IN3(n1385), .IN4(mul_exp_out[0]), 
        .IN5(n1752), .Q(n272) );
  INVX0 U1213 ( .INP(n1753), .ZN(n1752) );
  MUX21X1 U1214 ( .IN1(n1754), .IN2(n1755), .S(n1756), .Q(n1753) );
  NAND3X0 U1215 ( .IN1(n1757), .IN2(n1758), .IN3(n1759), .QN(n271) );
  MUX21X1 U1216 ( .IN1(n1760), .IN2(n1761), .S(m5stg_exp[8]), .Q(n1759) );
  OA21X1 U1217 ( .IN1(n1762), .IN2(n1755), .IN3(n1754), .Q(n1761) );
  NAND2X0 U1218 ( .IN1(n1762), .IN2(n1763), .QN(n1760) );
  NAND2X0 U1219 ( .IN1(n1405), .IN2(mul_exp_out[8]), .QN(n1757) );
  NAND3X0 U1220 ( .IN1(n1764), .IN2(n1758), .IN3(n1765), .QN(n270) );
  MUX21X1 U1221 ( .IN1(n1766), .IN2(n1767), .S(m5stg_exp[9]), .Q(n1765) );
  NAND2X0 U1222 ( .IN1(n1405), .IN2(mul_exp_out[9]), .QN(n1764) );
  NAND3X0 U1223 ( .IN1(n1768), .IN2(n1758), .IN3(n1769), .QN(n269) );
  MUX21X1 U1224 ( .IN1(n1770), .IN2(n1771), .S(m5stg_exp[10]), .Q(n1769) );
  OA21X1 U1225 ( .IN1(m5stg_exp[9]), .IN2(n1755), .IN3(n1767), .Q(n1771) );
  AND2X1 U1226 ( .IN1(n1772), .IN2(n1754), .Q(n1767) );
  NAND2X0 U1227 ( .IN1(n594), .IN2(n1773), .QN(n1754) );
  OA21X1 U1228 ( .IN1(n1774), .IN2(n1775), .IN3(n1608), .Q(n594) );
  AO21X1 U1229 ( .IN1(n1762), .IN2(m5stg_exp[8]), .IN3(n1755), .Q(n1772) );
  NAND2X0 U1230 ( .IN1(n1776), .IN2(m5stg_exp[9]), .QN(n1770) );
  INVX0 U1231 ( .INP(n1766), .ZN(n1776) );
  NAND3X0 U1232 ( .IN1(n1763), .IN2(m5stg_exp[8]), .IN3(n1762), .QN(n1766) );
  INVX0 U1233 ( .INP(n1777), .ZN(n1762) );
  NAND2X0 U1234 ( .IN1(n1750), .IN2(m5stg_fmuld), .QN(n1758) );
  INVX0 U1235 ( .INP(n1778), .ZN(n1750) );
  NAND2X0 U1236 ( .IN1(n1405), .IN2(mul_exp_out[10]), .QN(n1768) );
  OA221X1 U1237 ( .IN1(n1779), .IN2(n1755), .IN3(n10), .IN4(n1625), .IN5(n1778), .Q(n196) );
  XOR2X1 U1238 ( .IN1(m5stg_exp[0]), .IN2(n1780), .Q(n1779) );
  OA221X1 U1239 ( .IN1(n1755), .IN2(n1781), .IN3(n9), .IN4(n1625), .IN5(n1778), 
        .Q(n195) );
  NAND2X0 U1240 ( .IN1(n1782), .IN2(n1783), .QN(n1781) );
  AO21X1 U1241 ( .IN1(m5stg_exp[1]), .IN2(m5stg_exp[0]), .IN3(m5stg_exp[2]), 
        .Q(n1782) );
  OA221X1 U1242 ( .IN1(n1755), .IN2(n1784), .IN3(n8), .IN4(n1625), .IN5(n1778), 
        .Q(n194) );
  AO21X1 U1243 ( .IN1(n1783), .IN2(n1785), .IN3(n1786), .Q(n1784) );
  OA221X1 U1244 ( .IN1(n1755), .IN2(n1787), .IN3(n7), .IN4(n1625), .IN5(n1778), 
        .Q(n193) );
  OAI21X1 U1245 ( .IN1(n1786), .IN2(m5stg_exp[4]), .IN3(n1788), .QN(n1787) );
  OA221X1 U1246 ( .IN1(n1755), .IN2(n1789), .IN3(n6), .IN4(n1625), .IN5(n1778), 
        .Q(n192) );
  AO21X1 U1247 ( .IN1(n1788), .IN2(n1790), .IN3(n1791), .Q(n1789) );
  OA221X1 U1248 ( .IN1(n1755), .IN2(n1792), .IN3(n5), .IN4(n1625), .IN5(n1778), 
        .Q(n191) );
  XOR2X1 U1249 ( .IN1(n1793), .IN2(n1791), .Q(n1792) );
  OA221X1 U1250 ( .IN1(n1755), .IN2(n1794), .IN3(n4), .IN4(n1625), .IN5(n1778), 
        .Q(n190) );
  NAND2X0 U1251 ( .IN1(n1795), .IN2(n1777), .QN(n1794) );
  NAND3X0 U1252 ( .IN1(m5stg_exp[6]), .IN2(m5stg_exp[7]), .IN3(n1791), .QN(
        n1777) );
  AO21X1 U1253 ( .IN1(n1791), .IN2(m5stg_exp[6]), .IN3(m5stg_exp[7]), .Q(n1795) );
  INVX0 U1254 ( .INP(n1763), .ZN(n1755) );
  NOR2X0 U1255 ( .IN1(n1796), .IN2(n1774), .QN(n1763) );
  INVX0 U1256 ( .INP(n1797), .ZN(mul_exc_out[3]) );
  NAND2X0 U1257 ( .IN1(\fpu_mul_ctl/n28 ), .IN2(n1797), .QN(mul_exc_out[0]) );
  OA21X1 U1258 ( .IN1(\fpu_mul_ctl/n30 ), .IN2(\fpu_mul_ctl/n32 ), .IN3(
        \fpu_mul_ctl/n31 ), .Q(n1797) );
  MUX21X1 U1259 ( .IN1(n983), .IN2(n1217), .S(n1798), .Q(m6stg_id_in[1]) );
  MUX21X1 U1260 ( .IN1(n984), .IN2(n1216), .S(n1798), .Q(m6stg_id_in[0]) );
  OA21X1 U1261 ( .IN1(n1798), .IN2(\fpu_mul_ctl/m5stg_opdec[4] ), .IN3(n1209), 
        .Q(m6stg_fmul_in) );
  NOR4X0 U1262 ( .IN1(n1799), .IN2(n1800), .IN3(n1801), .IN4(n1802), .QN(
        m4stg_inc_exp_54) );
  NAND3X0 U1263 ( .IN1(n52), .IN2(n447), .IN3(n60), .QN(n1802) );
  NAND3X0 U1264 ( .IN1(n445), .IN2(n444), .IN3(n446), .QN(n1801) );
  NAND3X0 U1265 ( .IN1(n442), .IN2(n44), .IN3(n443), .QN(n1800) );
  NAND4X0 U1266 ( .IN1(n438), .IN2(n37), .IN3(n29), .IN4(m4stg_inc_exp_55), 
        .QN(n1799) );
  NOR3X0 U1267 ( .IN1(n979), .IN2(m4stg_inc_exp_55), .IN3(\fpu_mul_ctl/n1 ), 
        .QN(m4stg_inc_exp_105) );
  NAND4X0 U1268 ( .IN1(n1803), .IN2(n1804), .IN3(n1805), .IN4(n1806), .QN(
        m2stg_frac2_array_in[52]) );
  OA21X1 U1269 ( .IN1(\fpu_mul_frac_dp/n289 ), .IN2(n1807), .IN3(n1808), .Q(
        n1806) );
  NAND2X0 U1270 ( .IN1(n1809), .IN2(n1224), .QN(n1805) );
  AO221X1 U1271 ( .IN1(n1809), .IN2(n1151), .IN3(n1810), .IN4(n916), .IN5(
        n1811), .Q(m2stg_frac2_array_in[51]) );
  AO221X1 U1272 ( .IN1(n1812), .IN2(n1813), .IN3(n1814), .IN4(n1815), .IN5(
        n1816), .Q(n1811) );
  NAND2X0 U1273 ( .IN1(\fpu_mul_frac_dp/n289 ), .IN2(n1817), .QN(n1815) );
  NAND2X0 U1274 ( .IN1(\fpu_mul_frac_dp/n286 ), .IN2(n1818), .QN(n1813) );
  AO221X1 U1275 ( .IN1(n1814), .IN2(n916), .IN3(n1810), .IN4(n891), .IN5(n1819), .Q(m2stg_frac2_array_in[50]) );
  AO221X1 U1276 ( .IN1(n1809), .IN2(n942), .IN3(n1812), .IN4(n1151), .IN5(
        n1816), .Q(n1819) );
  AO221X1 U1277 ( .IN1(n1814), .IN2(n891), .IN3(n1810), .IN4(n1042), .IN5(
        n1820), .Q(m2stg_frac2_array_in[49]) );
  AO221X1 U1278 ( .IN1(n1809), .IN2(n1132), .IN3(n1812), .IN4(n942), .IN5(
        n1816), .Q(n1820) );
  AO221X1 U1279 ( .IN1(n1814), .IN2(n1042), .IN3(n1810), .IN4(n890), .IN5(
        n1821), .Q(m2stg_frac2_array_in[48]) );
  AO221X1 U1280 ( .IN1(n1809), .IN2(n916), .IN3(n1812), .IN4(n1132), .IN5(
        n1816), .Q(n1821) );
  AO221X1 U1281 ( .IN1(n1814), .IN2(n890), .IN3(n1810), .IN4(n918), .IN5(n1822), .Q(m2stg_frac2_array_in[47]) );
  AO221X1 U1282 ( .IN1(n1809), .IN2(n891), .IN3(n1812), .IN4(n916), .IN5(n1816), .Q(n1822) );
  AO221X1 U1283 ( .IN1(n1814), .IN2(n918), .IN3(n1810), .IN4(n1044), .IN5(
        n1823), .Q(m2stg_frac2_array_in[46]) );
  AO221X1 U1284 ( .IN1(n1809), .IN2(n1042), .IN3(n1812), .IN4(n891), .IN5(
        n1816), .Q(n1823) );
  AO221X1 U1285 ( .IN1(n1814), .IN2(n1044), .IN3(n1810), .IN4(n880), .IN5(
        n1824), .Q(m2stg_frac2_array_in[45]) );
  AO221X1 U1286 ( .IN1(n1809), .IN2(n890), .IN3(n1812), .IN4(n1042), .IN5(
        n1816), .Q(n1824) );
  AO221X1 U1287 ( .IN1(n1814), .IN2(n880), .IN3(n1810), .IN4(n917), .IN5(n1825), .Q(m2stg_frac2_array_in[44]) );
  AO221X1 U1288 ( .IN1(n1809), .IN2(n918), .IN3(n1812), .IN4(n890), .IN5(n1816), .Q(n1825) );
  AO221X1 U1289 ( .IN1(n1814), .IN2(n917), .IN3(n1810), .IN4(n1047), .IN5(
        n1826), .Q(m2stg_frac2_array_in[43]) );
  AO221X1 U1290 ( .IN1(n1809), .IN2(n1044), .IN3(n1812), .IN4(n918), .IN5(
        n1816), .Q(n1826) );
  AO221X1 U1291 ( .IN1(n1814), .IN2(n1047), .IN3(n1810), .IN4(n921), .IN5(
        n1827), .Q(m2stg_frac2_array_in[42]) );
  AO221X1 U1292 ( .IN1(n1809), .IN2(n880), .IN3(n1812), .IN4(n1044), .IN5(
        n1816), .Q(n1827) );
  AO221X1 U1293 ( .IN1(n1814), .IN2(n921), .IN3(n1810), .IN4(n1043), .IN5(
        n1828), .Q(m2stg_frac2_array_in[41]) );
  AO221X1 U1294 ( .IN1(n1809), .IN2(n917), .IN3(n1812), .IN4(n880), .IN5(n1816), .Q(n1828) );
  AO221X1 U1295 ( .IN1(n1814), .IN2(n1043), .IN3(n1810), .IN4(n889), .IN5(
        n1829), .Q(m2stg_frac2_array_in[40]) );
  AO221X1 U1296 ( .IN1(n1809), .IN2(n1047), .IN3(n1812), .IN4(n917), .IN5(
        n1816), .Q(n1829) );
  AO221X1 U1297 ( .IN1(n1814), .IN2(n889), .IN3(n1810), .IN4(n920), .IN5(n1830), .Q(m2stg_frac2_array_in[39]) );
  AO221X1 U1298 ( .IN1(n1809), .IN2(n921), .IN3(n1812), .IN4(n1047), .IN5(
        n1816), .Q(n1830) );
  AO221X1 U1299 ( .IN1(n1814), .IN2(n920), .IN3(n1810), .IN4(n1048), .IN5(
        n1831), .Q(m2stg_frac2_array_in[38]) );
  AO221X1 U1300 ( .IN1(n1809), .IN2(n1043), .IN3(n1812), .IN4(n921), .IN5(
        n1816), .Q(n1831) );
  AO221X1 U1301 ( .IN1(n1814), .IN2(n1048), .IN3(n1810), .IN4(n909), .IN5(
        n1832), .Q(m2stg_frac2_array_in[37]) );
  AO221X1 U1302 ( .IN1(n1809), .IN2(n889), .IN3(n1812), .IN4(n1043), .IN5(
        n1816), .Q(n1832) );
  AO221X1 U1303 ( .IN1(n1814), .IN2(n909), .IN3(n1810), .IN4(n1046), .IN5(
        n1833), .Q(m2stg_frac2_array_in[36]) );
  AO221X1 U1304 ( .IN1(n1809), .IN2(n920), .IN3(n1812), .IN4(n889), .IN5(n1816), .Q(n1833) );
  AO221X1 U1305 ( .IN1(n1814), .IN2(n1046), .IN3(n1810), .IN4(n919), .IN5(
        n1834), .Q(m2stg_frac2_array_in[35]) );
  AO221X1 U1306 ( .IN1(n1809), .IN2(n1048), .IN3(n1812), .IN4(n920), .IN5(
        n1816), .Q(n1834) );
  AO221X1 U1307 ( .IN1(n1814), .IN2(n919), .IN3(n1810), .IN4(n1045), .IN5(
        n1835), .Q(m2stg_frac2_array_in[34]) );
  AO221X1 U1308 ( .IN1(n1809), .IN2(n909), .IN3(n1812), .IN4(n1048), .IN5(
        n1816), .Q(n1835) );
  AO221X1 U1309 ( .IN1(n1814), .IN2(n1045), .IN3(n1810), .IN4(n887), .IN5(
        n1836), .Q(m2stg_frac2_array_in[33]) );
  AO221X1 U1310 ( .IN1(n1809), .IN2(n1046), .IN3(n1812), .IN4(n909), .IN5(
        n1816), .Q(n1836) );
  AO221X1 U1311 ( .IN1(n1814), .IN2(n887), .IN3(n1810), .IN4(n958), .IN5(n1837), .Q(m2stg_frac2_array_in[32]) );
  AO221X1 U1312 ( .IN1(n1809), .IN2(n919), .IN3(n1812), .IN4(n1046), .IN5(
        n1816), .Q(n1837) );
  OA22X1 U1313 ( .IN1(\fpu_mul_frac_dp/n752 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n781 ), .IN4(n1839), .Q(m2stg_frac1_array_in[9]) );
  OA22X1 U1314 ( .IN1(\fpu_mul_frac_dp/n781 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n828 ), .IN4(n1839), .Q(m2stg_frac1_array_in[8]) );
  OA22X1 U1315 ( .IN1(\fpu_mul_frac_dp/n787 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n828 ), .IN4(n1838), .Q(m2stg_frac1_array_in[7]) );
  OA22X1 U1316 ( .IN1(\fpu_mul_frac_dp/n756 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n787 ), .IN4(n1838), .Q(m2stg_frac1_array_in[6]) );
  OA22X1 U1317 ( .IN1(\fpu_mul_frac_dp/n756 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n806 ), .IN4(n1839), .Q(m2stg_frac1_array_in[5]) );
  NOR4X0 U1318 ( .IN1(n1840), .IN2(n1841), .IN3(n1842), .IN4(n1843), .QN(
        m2stg_frac1_array_in[52]) );
  NOR2X0 U1319 ( .IN1(\fpu_mul_frac_dp/n335 ), .IN2(n1844), .QN(n1843) );
  INVX0 U1320 ( .INP(n1845), .ZN(n1842) );
  AO22X1 U1321 ( .IN1(n1846), .IN2(n1847), .IN3(n1848), .IN4(n1124), .Q(n1841)
         );
  INVX0 U1322 ( .INP(n1839), .ZN(n1848) );
  NAND4X0 U1323 ( .IN1(n1818), .IN2(n1817), .IN3(n1849), .IN4(n1838), .QN(
        n1840) );
  OA221X1 U1324 ( .IN1(n1850), .IN2(n1838), .IN3(n1851), .IN4(n1849), .IN5(
        n1852), .Q(m2stg_frac1_array_in[51]) );
  OA22X1 U1325 ( .IN1(\fpu_mul_frac_dp/n336 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n339 ), .IN4(n1839), .Q(n1852) );
  NOR2X0 U1326 ( .IN1(n1853), .IN2(n1200), .QN(n1851) );
  NOR2X0 U1327 ( .IN1(n1854), .IN2(n1124), .QN(n1850) );
  OA221X1 U1328 ( .IN1(\fpu_mul_frac_dp/n339 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n337 ), .IN4(n1844), .IN5(n1855), .Q(
        m2stg_frac1_array_in[50]) );
  OA22X1 U1329 ( .IN1(\fpu_mul_frac_dp/n336 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n340 ), .IN4(n1839), .Q(n1855) );
  OA22X1 U1330 ( .IN1(\fpu_mul_frac_dp/n764 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n806 ), .IN4(n1838), .Q(m2stg_frac1_array_in[4]) );
  OA221X1 U1331 ( .IN1(\fpu_mul_frac_dp/n338 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n340 ), .IN4(n1838), .IN5(n1856), .Q(
        m2stg_frac1_array_in[49]) );
  OA22X1 U1332 ( .IN1(\fpu_mul_frac_dp/n337 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n341 ), .IN4(n1839), .Q(n1856) );
  OA221X1 U1333 ( .IN1(\fpu_mul_frac_dp/n341 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n339 ), .IN4(n1844), .IN5(n1857), .Q(
        m2stg_frac1_array_in[48]) );
  OA22X1 U1334 ( .IN1(\fpu_mul_frac_dp/n338 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n342 ), .IN4(n1839), .Q(n1857) );
  OA221X1 U1335 ( .IN1(\fpu_mul_frac_dp/n340 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n342 ), .IN4(n1838), .IN5(n1858), .Q(
        m2stg_frac1_array_in[47]) );
  OA22X1 U1336 ( .IN1(\fpu_mul_frac_dp/n339 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n343 ), .IN4(n1839), .Q(n1858) );
  OA221X1 U1337 ( .IN1(\fpu_mul_frac_dp/n343 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n341 ), .IN4(n1844), .IN5(n1859), .Q(
        m2stg_frac1_array_in[46]) );
  OA22X1 U1338 ( .IN1(\fpu_mul_frac_dp/n340 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n344 ), .IN4(n1839), .Q(n1859) );
  OA221X1 U1339 ( .IN1(\fpu_mul_frac_dp/n344 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n342 ), .IN4(n1844), .IN5(n1860), .Q(
        m2stg_frac1_array_in[45]) );
  OA22X1 U1340 ( .IN1(\fpu_mul_frac_dp/n341 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n345 ), .IN4(n1839), .Q(n1860) );
  OA221X1 U1341 ( .IN1(\fpu_mul_frac_dp/n345 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n342 ), .IN4(n1849), .IN5(n1861), .Q(
        m2stg_frac1_array_in[44]) );
  OA22X1 U1342 ( .IN1(\fpu_mul_frac_dp/n343 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n346 ), .IN4(n1839), .Q(n1861) );
  OA221X1 U1343 ( .IN1(\fpu_mul_frac_dp/n344 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n346 ), .IN4(n1838), .IN5(n1862), .Q(
        m2stg_frac1_array_in[43]) );
  OA22X1 U1344 ( .IN1(\fpu_mul_frac_dp/n343 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n347 ), .IN4(n1839), .Q(n1862) );
  OA221X1 U1345 ( .IN1(\fpu_mul_frac_dp/n347 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n345 ), .IN4(n1844), .IN5(n1863), .Q(
        m2stg_frac1_array_in[42]) );
  OA22X1 U1346 ( .IN1(\fpu_mul_frac_dp/n344 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n348 ), .IN4(n1839), .Q(n1863) );
  OA221X1 U1347 ( .IN1(\fpu_mul_frac_dp/n346 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n348 ), .IN4(n1838), .IN5(n1864), .Q(
        m2stg_frac1_array_in[41]) );
  OA22X1 U1348 ( .IN1(\fpu_mul_frac_dp/n345 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n349 ), .IN4(n1839), .Q(n1864) );
  OA221X1 U1349 ( .IN1(\fpu_mul_frac_dp/n347 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n349 ), .IN4(n1838), .IN5(n1865), .Q(
        m2stg_frac1_array_in[40]) );
  OA22X1 U1350 ( .IN1(\fpu_mul_frac_dp/n346 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n350 ), .IN4(n1839), .Q(n1865) );
  OA22X1 U1351 ( .IN1(\fpu_mul_frac_dp/n764 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n792 ), .IN4(n1839), .Q(m2stg_frac1_array_in[3]) );
  OA221X1 U1352 ( .IN1(\fpu_mul_frac_dp/n348 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n350 ), .IN4(n1838), .IN5(n1866), .Q(
        m2stg_frac1_array_in[39]) );
  OA22X1 U1353 ( .IN1(\fpu_mul_frac_dp/n347 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n351 ), .IN4(n1839), .Q(n1866) );
  OA221X1 U1354 ( .IN1(\fpu_mul_frac_dp/n351 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n348 ), .IN4(n1849), .IN5(n1867), .Q(
        m2stg_frac1_array_in[38]) );
  OA22X1 U1355 ( .IN1(\fpu_mul_frac_dp/n349 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n352 ), .IN4(n1839), .Q(n1867) );
  OA221X1 U1356 ( .IN1(\fpu_mul_frac_dp/n350 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n352 ), .IN4(n1838), .IN5(n1868), .Q(
        m2stg_frac1_array_in[37]) );
  OA22X1 U1357 ( .IN1(\fpu_mul_frac_dp/n349 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n353 ), .IN4(n1839), .Q(n1868) );
  OA221X1 U1358 ( .IN1(\fpu_mul_frac_dp/n351 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n353 ), .IN4(n1838), .IN5(n1869), .Q(
        m2stg_frac1_array_in[36]) );
  OA22X1 U1359 ( .IN1(\fpu_mul_frac_dp/n350 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n354 ), .IN4(n1839), .Q(n1869) );
  OA221X1 U1360 ( .IN1(\fpu_mul_frac_dp/n352 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n354 ), .IN4(n1838), .IN5(n1870), .Q(
        m2stg_frac1_array_in[35]) );
  OA22X1 U1361 ( .IN1(\fpu_mul_frac_dp/n351 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n355 ), .IN4(n1839), .Q(n1870) );
  OA221X1 U1362 ( .IN1(\fpu_mul_frac_dp/n355 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n353 ), .IN4(n1844), .IN5(n1871), .Q(
        m2stg_frac1_array_in[34]) );
  OA22X1 U1363 ( .IN1(\fpu_mul_frac_dp/n352 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n356 ), .IN4(n1839), .Q(n1871) );
  OA221X1 U1364 ( .IN1(\fpu_mul_frac_dp/n356 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n353 ), .IN4(n1849), .IN5(n1872), .Q(
        m2stg_frac1_array_in[33]) );
  OA22X1 U1365 ( .IN1(\fpu_mul_frac_dp/n354 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n357 ), .IN4(n1839), .Q(n1872) );
  OA221X1 U1366 ( .IN1(\fpu_mul_frac_dp/n357 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n354 ), .IN4(n1849), .IN5(n1873), .Q(
        m2stg_frac1_array_in[32]) );
  OA22X1 U1367 ( .IN1(\fpu_mul_frac_dp/n355 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n358 ), .IN4(n1839), .Q(n1873) );
  OA221X1 U1368 ( .IN1(\fpu_mul_frac_dp/n356 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n358 ), .IN4(n1838), .IN5(n1874), .Q(
        m2stg_frac1_array_in[31]) );
  OA22X1 U1369 ( .IN1(\fpu_mul_frac_dp/n355 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n359 ), .IN4(n1839), .Q(n1874) );
  OA221X1 U1370 ( .IN1(\fpu_mul_frac_dp/n357 ), .IN2(n1844), .IN3(
        \fpu_mul_frac_dp/n359 ), .IN4(n1838), .IN5(n1875), .Q(
        m2stg_frac1_array_in[30]) );
  OA22X1 U1371 ( .IN1(\fpu_mul_frac_dp/n356 ), .IN2(n1849), .IN3(
        \fpu_mul_frac_dp/n360 ), .IN4(n1839), .Q(n1875) );
  NAND3X0 U1372 ( .IN1(n1876), .IN2(n910), .IN3(\fpu_mul_ctl/n263 ), .QN(n1844) );
  OA22X1 U1373 ( .IN1(\fpu_mul_frac_dp/n792 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n827 ), .IN4(n1839), .Q(m2stg_frac1_array_in[2]) );
  OA222X1 U1374 ( .IN1(\fpu_mul_frac_dp/n357 ), .IN2(n1849), .IN3(n1839), 
        .IN4(n1207), .IN5(\fpu_mul_frac_dp/n360 ), .IN6(n1838), .Q(
        m2stg_frac1_array_in[29]) );
  NAND3X0 U1375 ( .IN1(n910), .IN2(n1163), .IN3(n1877), .QN(n1849) );
  NAND3X0 U1376 ( .IN1(n1878), .IN2(n1879), .IN3(n1880), .QN(n1877) );
  NAND4X0 U1377 ( .IN1(\fpu_mul_ctl/n256 ), .IN2(n1881), .IN3(n923), .IN4(n894), .QN(n1879) );
  NAND2X0 U1378 ( .IN1(n1853), .IN2(n1818), .QN(n1878) );
  OA22X1 U1379 ( .IN1(\fpu_mul_frac_dp/n785 ), .IN2(n1839), .IN3(n1838), .IN4(
        n1207), .Q(m2stg_frac1_array_in[28]) );
  OA22X1 U1380 ( .IN1(\fpu_mul_frac_dp/n785 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n810 ), .IN4(n1839), .Q(m2stg_frac1_array_in[27]) );
  OA22X1 U1381 ( .IN1(\fpu_mul_frac_dp/n796 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n810 ), .IN4(n1838), .Q(m2stg_frac1_array_in[26]) );
  OA22X1 U1382 ( .IN1(\fpu_mul_frac_dp/n796 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n823 ), .IN4(n1839), .Q(m2stg_frac1_array_in[25]) );
  OA22X1 U1383 ( .IN1(\fpu_mul_frac_dp/n786 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n823 ), .IN4(n1838), .Q(m2stg_frac1_array_in[24]) );
  OA22X1 U1384 ( .IN1(\fpu_mul_frac_dp/n786 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n825 ), .IN4(n1839), .Q(m2stg_frac1_array_in[23]) );
  OA22X1 U1385 ( .IN1(\fpu_mul_frac_dp/n763 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n825 ), .IN4(n1838), .Q(m2stg_frac1_array_in[22]) );
  OA22X1 U1386 ( .IN1(\fpu_mul_frac_dp/n763 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n829 ), .IN4(n1839), .Q(m2stg_frac1_array_in[21]) );
  OA22X1 U1387 ( .IN1(\fpu_mul_frac_dp/n759 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n829 ), .IN4(n1838), .Q(m2stg_frac1_array_in[20]) );
  OA22X1 U1388 ( .IN1(\fpu_mul_frac_dp/n382 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n827 ), .IN4(n1838), .Q(m2stg_frac1_array_in[1]) );
  OA22X1 U1389 ( .IN1(\fpu_mul_frac_dp/n759 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n805 ), .IN4(n1839), .Q(m2stg_frac1_array_in[19]) );
  OA22X1 U1390 ( .IN1(\fpu_mul_frac_dp/n751 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n805 ), .IN4(n1838), .Q(m2stg_frac1_array_in[18]) );
  OA22X1 U1391 ( .IN1(\fpu_mul_frac_dp/n751 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n778 ), .IN4(n1839), .Q(m2stg_frac1_array_in[17]) );
  OA22X1 U1392 ( .IN1(\fpu_mul_frac_dp/n778 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n807 ), .IN4(n1839), .Q(m2stg_frac1_array_in[16]) );
  OA22X1 U1393 ( .IN1(\fpu_mul_frac_dp/n795 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n807 ), .IN4(n1838), .Q(m2stg_frac1_array_in[15]) );
  OA22X1 U1394 ( .IN1(\fpu_mul_frac_dp/n795 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n821 ), .IN4(n1839), .Q(m2stg_frac1_array_in[14]) );
  OA22X1 U1395 ( .IN1(\fpu_mul_frac_dp/n821 ), .IN2(n1838), .IN3(n1839), .IN4(
        n1283), .Q(m2stg_frac1_array_in[13]) );
  OA22X1 U1396 ( .IN1(\fpu_mul_frac_dp/n760 ), .IN2(n1839), .IN3(n1838), .IN4(
        n1283), .Q(m2stg_frac1_array_in[12]) );
  OA22X1 U1397 ( .IN1(\fpu_mul_frac_dp/n760 ), .IN2(n1838), .IN3(
        \fpu_mul_frac_dp/n802 ), .IN4(n1839), .Q(m2stg_frac1_array_in[11]) );
  OA22X1 U1398 ( .IN1(\fpu_mul_frac_dp/n752 ), .IN2(n1839), .IN3(
        \fpu_mul_frac_dp/n802 ), .IN4(n1838), .Q(m2stg_frac1_array_in[10]) );
  NAND3X0 U1399 ( .IN1(n1882), .IN2(n886), .IN3(\fpu_mul_ctl/n263 ), .QN(n1839) );
  OR2X1 U1400 ( .IN1(n1838), .IN2(\fpu_mul_frac_dp/n382 ), .Q(
        m2stg_frac1_array_in[0]) );
  NAND3X0 U1401 ( .IN1(n886), .IN2(n1163), .IN3(n1883), .QN(n1838) );
  NAND3X0 U1402 ( .IN1(n1884), .IN2(n1885), .IN3(n1886), .QN(n1883) );
  NAND4X0 U1403 ( .IN1(\fpu_mul_ctl/n256 ), .IN2(n1887), .IN3(n922), .IN4(n893), .QN(n1885) );
  NAND2X0 U1404 ( .IN1(n1854), .IN2(n1817), .QN(n1884) );
  AND3X1 U1405 ( .IN1(n1680), .IN2(n1679), .IN3(\fpu_mul_ctl/n257 ), .Q(
        m2stg_exp_017f) );
  NOR2X0 U1406 ( .IN1(n1888), .IN2(n1374), .QN(\i_m4stg_frac/psum_dff/N9 ) );
  NOR2X0 U1407 ( .IN1(n1374), .IN2(n1889), .QN(\i_m4stg_frac/psum_dff/N8 ) );
  NOR2X0 U1408 ( .IN1(\i_m4stg_frac/n1462 ), .IN2(n1373), .QN(
        \i_m4stg_frac/psum_dff/N70 ) );
  NOR2X0 U1409 ( .IN1(n1373), .IN2(n1890), .QN(\i_m4stg_frac/psum_dff/N7 ) );
  NOR2X0 U1410 ( .IN1(n1376), .IN2(n1891), .QN(\i_m4stg_frac/psum_dff/N69 ) );
  XOR2X1 U1411 ( .IN1(\i_m4stg_frac/n490 ), .IN2(n1892), .Q(n1891) );
  NOR3X0 U1412 ( .IN1(n1374), .IN2(n1893), .IN3(n1894), .QN(
        \i_m4stg_frac/psum_dff/N68 ) );
  OA21X1 U1413 ( .IN1(n1892), .IN2(n1895), .IN3(n1896), .Q(n1894) );
  AND3X1 U1414 ( .IN1(n1897), .IN2(n1898), .IN3(n1899), .Q(
        \i_m4stg_frac/psum_dff/N67 ) );
  OAI21X1 U1415 ( .IN1(n1900), .IN2(n1901), .IN3(n1902), .QN(n1899) );
  AND2X1 U1416 ( .IN1(\i_m4stg_frac/n340 ), .IN2(\i_m4stg_frac/n494 ), .Q(
        n1901) );
  AND3X1 U1417 ( .IN1(n1897), .IN2(n1903), .IN3(n1904), .Q(
        \i_m4stg_frac/psum_dff/N66 ) );
  OAI21X1 U1418 ( .IN1(n1905), .IN2(n1906), .IN3(n1907), .QN(n1904) );
  AND2X1 U1419 ( .IN1(\i_m4stg_frac/n342 ), .IN2(\i_m4stg_frac/n496 ), .Q(
        n1906) );
  AND3X1 U1420 ( .IN1(n1897), .IN2(n1908), .IN3(n1909), .Q(
        \i_m4stg_frac/psum_dff/N65 ) );
  OAI21X1 U1421 ( .IN1(n1910), .IN2(n1911), .IN3(n1912), .QN(n1909) );
  AND2X1 U1422 ( .IN1(\i_m4stg_frac/n344 ), .IN2(\i_m4stg_frac/n498 ), .Q(
        n1911) );
  AND3X1 U1423 ( .IN1(n1897), .IN2(n1913), .IN3(n1914), .Q(
        \i_m4stg_frac/psum_dff/N64 ) );
  OAI21X1 U1424 ( .IN1(n1915), .IN2(n1916), .IN3(n1917), .QN(n1914) );
  AND2X1 U1425 ( .IN1(\i_m4stg_frac/n346 ), .IN2(\i_m4stg_frac/n500 ), .Q(
        n1916) );
  AND3X1 U1426 ( .IN1(n1897), .IN2(n1918), .IN3(n1919), .Q(
        \i_m4stg_frac/psum_dff/N63 ) );
  OAI21X1 U1427 ( .IN1(n1920), .IN2(n1921), .IN3(n1922), .QN(n1919) );
  AND2X1 U1428 ( .IN1(\i_m4stg_frac/n348 ), .IN2(\i_m4stg_frac/n502 ), .Q(
        n1921) );
  AND3X1 U1429 ( .IN1(n1897), .IN2(n1923), .IN3(n1924), .Q(
        \i_m4stg_frac/psum_dff/N62 ) );
  OAI21X1 U1430 ( .IN1(n1925), .IN2(n1926), .IN3(n1927), .QN(n1924) );
  AND2X1 U1431 ( .IN1(\i_m4stg_frac/n350 ), .IN2(\i_m4stg_frac/n504 ), .Q(
        n1926) );
  AND3X1 U1432 ( .IN1(n1897), .IN2(n1928), .IN3(n1929), .Q(
        \i_m4stg_frac/psum_dff/N61 ) );
  OAI21X1 U1433 ( .IN1(n1930), .IN2(n1931), .IN3(n1932), .QN(n1929) );
  AND2X1 U1434 ( .IN1(\i_m4stg_frac/n352 ), .IN2(\i_m4stg_frac/n506 ), .Q(
        n1931) );
  AND3X1 U1435 ( .IN1(n1897), .IN2(n1933), .IN3(n1934), .Q(
        \i_m4stg_frac/psum_dff/N60 ) );
  OAI21X1 U1436 ( .IN1(n1935), .IN2(n1936), .IN3(n1937), .QN(n1934) );
  AND2X1 U1437 ( .IN1(\i_m4stg_frac/n354 ), .IN2(\i_m4stg_frac/n508 ), .Q(
        n1936) );
  NOR2X0 U1438 ( .IN1(n1375), .IN2(n1938), .QN(\i_m4stg_frac/psum_dff/N6 ) );
  AND3X1 U1439 ( .IN1(n1897), .IN2(n1939), .IN3(n1940), .Q(
        \i_m4stg_frac/psum_dff/N59 ) );
  AO21X1 U1440 ( .IN1(n1937), .IN2(n1941), .IN3(n1942), .Q(n1940) );
  AND3X1 U1441 ( .IN1(n1897), .IN2(n1943), .IN3(n1944), .Q(
        \i_m4stg_frac/psum_dff/N58 ) );
  OAI22X1 U1442 ( .IN1(n1942), .IN2(n1945), .IN3(\i_m4stg_frac/n514 ), .IN4(
        \i_m4stg_frac/n360 ), .QN(n1944) );
  NOR2X0 U1443 ( .IN1(n1946), .IN2(n1376), .QN(\i_m4stg_frac/psum_dff/N57 ) );
  XNOR2X1 U1444 ( .IN1(n1947), .IN2(n1948), .Q(n1946) );
  NOR3X0 U1445 ( .IN1(n1373), .IN2(n1949), .IN3(n1950), .QN(
        \i_m4stg_frac/psum_dff/N56 ) );
  OA21X1 U1446 ( .IN1(n1947), .IN2(n1951), .IN3(n1952), .Q(n1950) );
  NOR2X0 U1447 ( .IN1(n1953), .IN2(n1375), .QN(\i_m4stg_frac/psum_dff/N55 ) );
  XOR2X1 U1448 ( .IN1(n1954), .IN2(n1955), .Q(n1953) );
  AND3X1 U1449 ( .IN1(n1897), .IN2(n1956), .IN3(n1957), .Q(
        \i_m4stg_frac/psum_dff/N54 ) );
  OAI21X1 U1450 ( .IN1(n1958), .IN2(n1959), .IN3(n1960), .QN(n1957) );
  AND2X1 U1451 ( .IN1(n1961), .IN2(n1962), .Q(n1959) );
  AND3X1 U1452 ( .IN1(n1897), .IN2(n1963), .IN3(n1964), .Q(
        \i_m4stg_frac/psum_dff/N53 ) );
  OAI21X1 U1453 ( .IN1(n1965), .IN2(n1966), .IN3(n1967), .QN(n1964) );
  AND2X1 U1454 ( .IN1(n1968), .IN2(n1969), .Q(n1966) );
  AND3X1 U1455 ( .IN1(n1897), .IN2(n1970), .IN3(n1971), .Q(
        \i_m4stg_frac/psum_dff/N52 ) );
  OAI21X1 U1456 ( .IN1(n1972), .IN2(n1973), .IN3(n1974), .QN(n1971) );
  AND2X1 U1457 ( .IN1(n1975), .IN2(n1976), .Q(n1973) );
  AND3X1 U1458 ( .IN1(n1897), .IN2(n1977), .IN3(n1978), .Q(
        \i_m4stg_frac/psum_dff/N51 ) );
  OAI21X1 U1459 ( .IN1(n1979), .IN2(n1980), .IN3(n1981), .QN(n1978) );
  AND2X1 U1460 ( .IN1(n1982), .IN2(n1983), .Q(n1980) );
  AND3X1 U1461 ( .IN1(n1897), .IN2(n1984), .IN3(n1985), .Q(
        \i_m4stg_frac/psum_dff/N50 ) );
  OAI21X1 U1462 ( .IN1(n1986), .IN2(n1987), .IN3(n1988), .QN(n1985) );
  AND2X1 U1463 ( .IN1(n1989), .IN2(n1990), .Q(n1987) );
  NOR2X0 U1464 ( .IN1(n1374), .IN2(n1991), .QN(\i_m4stg_frac/psum_dff/N5 ) );
  AND3X1 U1465 ( .IN1(n1897), .IN2(n1992), .IN3(n1993), .Q(
        \i_m4stg_frac/psum_dff/N49 ) );
  OAI21X1 U1466 ( .IN1(n1994), .IN2(n1995), .IN3(n1996), .QN(n1993) );
  AND2X1 U1467 ( .IN1(n1997), .IN2(n1998), .Q(n1995) );
  AND3X1 U1468 ( .IN1(n1897), .IN2(n1999), .IN3(n2000), .Q(
        \i_m4stg_frac/psum_dff/N48 ) );
  OAI21X1 U1469 ( .IN1(n2001), .IN2(n2002), .IN3(n2003), .QN(n2000) );
  AND2X1 U1470 ( .IN1(n2004), .IN2(n2005), .Q(n2002) );
  AND3X1 U1471 ( .IN1(n1897), .IN2(n2006), .IN3(n2007), .Q(
        \i_m4stg_frac/psum_dff/N47 ) );
  OAI21X1 U1472 ( .IN1(n2008), .IN2(n2009), .IN3(n2010), .QN(n2007) );
  AND2X1 U1473 ( .IN1(n2011), .IN2(n2012), .Q(n2009) );
  AND3X1 U1474 ( .IN1(n1897), .IN2(n2013), .IN3(n2014), .Q(
        \i_m4stg_frac/psum_dff/N46 ) );
  OAI21X1 U1475 ( .IN1(n2015), .IN2(n2016), .IN3(n2017), .QN(n2014) );
  AND2X1 U1476 ( .IN1(n2018), .IN2(n2019), .Q(n2016) );
  NOR2X0 U1477 ( .IN1(n1373), .IN2(n2020), .QN(\i_m4stg_frac/psum_dff/N45 ) );
  NOR2X0 U1478 ( .IN1(n1376), .IN2(n2021), .QN(\i_m4stg_frac/psum_dff/N44 ) );
  NOR2X0 U1479 ( .IN1(n1375), .IN2(n2022), .QN(\i_m4stg_frac/psum_dff/N43 ) );
  NOR2X0 U1480 ( .IN1(n1374), .IN2(n2023), .QN(\i_m4stg_frac/psum_dff/N42 ) );
  NOR2X0 U1481 ( .IN1(n1373), .IN2(n2024), .QN(\i_m4stg_frac/psum_dff/N41 ) );
  NOR2X0 U1482 ( .IN1(n1376), .IN2(n2025), .QN(\i_m4stg_frac/psum_dff/N40 ) );
  NOR2X0 U1483 ( .IN1(n1375), .IN2(n2026), .QN(\i_m4stg_frac/psum_dff/N4 ) );
  NOR2X0 U1484 ( .IN1(n2027), .IN2(n1376), .QN(\i_m4stg_frac/psum_dff/N39 ) );
  NOR2X0 U1485 ( .IN1(n1374), .IN2(n2028), .QN(\i_m4stg_frac/psum_dff/N38 ) );
  NOR2X0 U1486 ( .IN1(n1373), .IN2(n2029), .QN(\i_m4stg_frac/psum_dff/N37 ) );
  NOR2X0 U1487 ( .IN1(n1376), .IN2(n2030), .QN(\i_m4stg_frac/psum_dff/N36 ) );
  NOR2X0 U1488 ( .IN1(n1375), .IN2(n2031), .QN(\i_m4stg_frac/psum_dff/N35 ) );
  NOR2X0 U1489 ( .IN1(n1374), .IN2(n2032), .QN(\i_m4stg_frac/psum_dff/N34 ) );
  NOR2X0 U1490 ( .IN1(n1373), .IN2(n2033), .QN(\i_m4stg_frac/psum_dff/N33 ) );
  NOR2X0 U1491 ( .IN1(n1376), .IN2(n2034), .QN(\i_m4stg_frac/psum_dff/N32 ) );
  NOR2X0 U1492 ( .IN1(n1375), .IN2(n2035), .QN(\i_m4stg_frac/psum_dff/N31 ) );
  NOR2X0 U1493 ( .IN1(n1374), .IN2(n2036), .QN(\i_m4stg_frac/psum_dff/N30 ) );
  NOR2X0 U1494 ( .IN1(n1373), .IN2(n2037), .QN(\i_m4stg_frac/psum_dff/N29 ) );
  NOR2X0 U1495 ( .IN1(n1376), .IN2(n2038), .QN(\i_m4stg_frac/psum_dff/N28 ) );
  NOR2X0 U1496 ( .IN1(n1375), .IN2(n2039), .QN(\i_m4stg_frac/psum_dff/N27 ) );
  NOR2X0 U1497 ( .IN1(n1374), .IN2(n2040), .QN(\i_m4stg_frac/psum_dff/N26 ) );
  NOR2X0 U1498 ( .IN1(n1373), .IN2(n2041), .QN(\i_m4stg_frac/psum_dff/N25 ) );
  NOR2X0 U1499 ( .IN1(n1376), .IN2(n2042), .QN(\i_m4stg_frac/psum_dff/N24 ) );
  NOR2X0 U1500 ( .IN1(n1375), .IN2(n2043), .QN(\i_m4stg_frac/psum_dff/N23 ) );
  NOR2X0 U1501 ( .IN1(n1374), .IN2(n2044), .QN(\i_m4stg_frac/psum_dff/N22 ) );
  NOR2X0 U1502 ( .IN1(n1373), .IN2(n2045), .QN(\i_m4stg_frac/psum_dff/N21 ) );
  NOR2X0 U1503 ( .IN1(n1376), .IN2(n2046), .QN(\i_m4stg_frac/psum_dff/N20 ) );
  NOR2X0 U1504 ( .IN1(n1375), .IN2(n2047), .QN(\i_m4stg_frac/psum_dff/N19 ) );
  NOR2X0 U1505 ( .IN1(n1374), .IN2(n2048), .QN(\i_m4stg_frac/psum_dff/N18 ) );
  NOR2X0 U1506 ( .IN1(n1373), .IN2(n2049), .QN(\i_m4stg_frac/psum_dff/N17 ) );
  NOR2X0 U1507 ( .IN1(n1376), .IN2(n2050), .QN(\i_m4stg_frac/psum_dff/N16 ) );
  NOR2X0 U1508 ( .IN1(n1375), .IN2(n2051), .QN(\i_m4stg_frac/psum_dff/N15 ) );
  NOR2X0 U1509 ( .IN1(n1374), .IN2(n2052), .QN(\i_m4stg_frac/psum_dff/N14 ) );
  NOR2X0 U1510 ( .IN1(n1373), .IN2(n2053), .QN(\i_m4stg_frac/psum_dff/N13 ) );
  NOR2X0 U1511 ( .IN1(n1376), .IN2(n2054), .QN(\i_m4stg_frac/psum_dff/N12 ) );
  NOR2X0 U1512 ( .IN1(n1375), .IN2(n2055), .QN(\i_m4stg_frac/psum_dff/N11 ) );
  NOR2X0 U1513 ( .IN1(n1374), .IN2(n2056), .QN(\i_m4stg_frac/psum_dff/N10 ) );
  NOR3X0 U1514 ( .IN1(n2057), .IN2(n1376), .IN3(n2058), .QN(
        \i_m4stg_frac/pcout_dff/N9 ) );
  NOR3X0 U1515 ( .IN1(n2059), .IN2(n1375), .IN3(n2060), .QN(
        \i_m4stg_frac/pcout_dff/N8 ) );
  AND3X1 U1516 ( .IN1(n1897), .IN2(n1339), .IN3(n1892), .Q(
        \i_m4stg_frac/pcout_dff/N70 ) );
  NOR3X0 U1517 ( .IN1(n2061), .IN2(n1374), .IN3(n2062), .QN(
        \i_m4stg_frac/pcout_dff/N7 ) );
  AND2X1 U1518 ( .IN1(n1897), .IN2(n1893), .Q(\i_m4stg_frac/pcout_dff/N69 ) );
  NOR3X0 U1519 ( .IN1(n1895), .IN2(n1892), .IN3(n1896), .QN(n1893) );
  NOR2X0 U1520 ( .IN1(\i_m4stg_frac/n837 ), .IN2(\i_m4stg_frac/n338 ), .QN(
        n1892) );
  AND2X1 U1521 ( .IN1(\i_m4stg_frac/n837 ), .IN2(\i_m4stg_frac/n338 ), .Q(
        n1895) );
  NOR2X0 U1522 ( .IN1(n1373), .IN2(n1898), .QN(\i_m4stg_frac/pcout_dff/N68 )
         );
  NAND3X0 U1523 ( .IN1(n2063), .IN2(n1896), .IN3(n1905), .QN(n1898) );
  INVX0 U1524 ( .INP(n1900), .ZN(n1896) );
  NOR2X0 U1525 ( .IN1(\i_m4stg_frac/n340 ), .IN2(\i_m4stg_frac/n494 ), .QN(
        n1900) );
  NAND2X0 U1526 ( .IN1(\i_m4stg_frac/n494 ), .IN2(\i_m4stg_frac/n340 ), .QN(
        n2063) );
  NOR2X0 U1527 ( .IN1(n1376), .IN2(n1903), .QN(\i_m4stg_frac/pcout_dff/N67 )
         );
  NAND3X0 U1528 ( .IN1(n2064), .IN2(n1902), .IN3(n1910), .QN(n1903) );
  INVX0 U1529 ( .INP(n1905), .ZN(n1902) );
  NOR2X0 U1530 ( .IN1(\i_m4stg_frac/n342 ), .IN2(\i_m4stg_frac/n496 ), .QN(
        n1905) );
  NAND2X0 U1531 ( .IN1(\i_m4stg_frac/n496 ), .IN2(\i_m4stg_frac/n342 ), .QN(
        n2064) );
  NOR2X0 U1532 ( .IN1(n1375), .IN2(n1908), .QN(\i_m4stg_frac/pcout_dff/N66 )
         );
  NAND3X0 U1533 ( .IN1(n2065), .IN2(n1907), .IN3(n1915), .QN(n1908) );
  INVX0 U1534 ( .INP(n1910), .ZN(n1907) );
  NOR2X0 U1535 ( .IN1(\i_m4stg_frac/n344 ), .IN2(\i_m4stg_frac/n498 ), .QN(
        n1910) );
  NAND2X0 U1536 ( .IN1(\i_m4stg_frac/n498 ), .IN2(\i_m4stg_frac/n344 ), .QN(
        n2065) );
  NOR2X0 U1537 ( .IN1(n1374), .IN2(n1913), .QN(\i_m4stg_frac/pcout_dff/N65 )
         );
  NAND3X0 U1538 ( .IN1(n2066), .IN2(n1912), .IN3(n1920), .QN(n1913) );
  INVX0 U1539 ( .INP(n1915), .ZN(n1912) );
  NOR2X0 U1540 ( .IN1(\i_m4stg_frac/n346 ), .IN2(\i_m4stg_frac/n500 ), .QN(
        n1915) );
  NAND2X0 U1541 ( .IN1(\i_m4stg_frac/n500 ), .IN2(\i_m4stg_frac/n346 ), .QN(
        n2066) );
  NOR2X0 U1542 ( .IN1(n1373), .IN2(n1918), .QN(\i_m4stg_frac/pcout_dff/N64 )
         );
  NAND3X0 U1543 ( .IN1(n2067), .IN2(n1917), .IN3(n1925), .QN(n1918) );
  INVX0 U1544 ( .INP(n1920), .ZN(n1917) );
  NOR2X0 U1545 ( .IN1(\i_m4stg_frac/n348 ), .IN2(\i_m4stg_frac/n502 ), .QN(
        n1920) );
  NAND2X0 U1546 ( .IN1(\i_m4stg_frac/n502 ), .IN2(\i_m4stg_frac/n348 ), .QN(
        n2067) );
  NOR2X0 U1547 ( .IN1(n1376), .IN2(n1923), .QN(\i_m4stg_frac/pcout_dff/N63 )
         );
  NAND3X0 U1548 ( .IN1(n2068), .IN2(n1922), .IN3(n1930), .QN(n1923) );
  INVX0 U1549 ( .INP(n1925), .ZN(n1922) );
  NOR2X0 U1550 ( .IN1(\i_m4stg_frac/n350 ), .IN2(\i_m4stg_frac/n504 ), .QN(
        n1925) );
  NAND2X0 U1551 ( .IN1(\i_m4stg_frac/n504 ), .IN2(\i_m4stg_frac/n350 ), .QN(
        n2068) );
  NOR2X0 U1552 ( .IN1(n1375), .IN2(n1928), .QN(\i_m4stg_frac/pcout_dff/N62 )
         );
  NAND3X0 U1553 ( .IN1(n2069), .IN2(n1927), .IN3(n1935), .QN(n1928) );
  INVX0 U1554 ( .INP(n1930), .ZN(n1927) );
  NOR2X0 U1555 ( .IN1(\i_m4stg_frac/n352 ), .IN2(\i_m4stg_frac/n506 ), .QN(
        n1930) );
  NAND2X0 U1556 ( .IN1(\i_m4stg_frac/n506 ), .IN2(\i_m4stg_frac/n352 ), .QN(
        n2069) );
  NOR2X0 U1557 ( .IN1(n1374), .IN2(n1933), .QN(\i_m4stg_frac/pcout_dff/N61 )
         );
  NAND3X0 U1558 ( .IN1(n2070), .IN2(n1932), .IN3(n2071), .QN(n1933) );
  INVX0 U1559 ( .INP(n1935), .ZN(n1932) );
  NOR2X0 U1560 ( .IN1(\i_m4stg_frac/n354 ), .IN2(\i_m4stg_frac/n508 ), .QN(
        n1935) );
  NAND2X0 U1561 ( .IN1(\i_m4stg_frac/n508 ), .IN2(\i_m4stg_frac/n354 ), .QN(
        n2070) );
  NOR2X0 U1562 ( .IN1(n1373), .IN2(n1939), .QN(\i_m4stg_frac/pcout_dff/N60 )
         );
  NAND3X0 U1563 ( .IN1(n1941), .IN2(n1937), .IN3(n1942), .QN(n1939) );
  INVX0 U1564 ( .INP(n2071), .ZN(n1937) );
  NOR2X0 U1565 ( .IN1(\i_m4stg_frac/n356 ), .IN2(\i_m4stg_frac/n510 ), .QN(
        n2071) );
  NAND2X0 U1566 ( .IN1(\i_m4stg_frac/n356 ), .IN2(\i_m4stg_frac/n510 ), .QN(
        n1941) );
  NOR3X0 U1567 ( .IN1(n2072), .IN2(n1373), .IN3(n2073), .QN(
        \i_m4stg_frac/pcout_dff/N6 ) );
  NOR2X0 U1568 ( .IN1(n1376), .IN2(n1943), .QN(\i_m4stg_frac/pcout_dff/N59 )
         );
  OR4X1 U1569 ( .IN1(n1945), .IN2(n1942), .IN3(\i_m4stg_frac/n360 ), .IN4(
        \i_m4stg_frac/n514 ), .Q(n1943) );
  NOR2X0 U1570 ( .IN1(\i_m4stg_frac/n358 ), .IN2(\i_m4stg_frac/n512 ), .QN(
        n1942) );
  AND2X1 U1571 ( .IN1(\i_m4stg_frac/n358 ), .IN2(\i_m4stg_frac/n512 ), .Q(
        n1945) );
  AND3X1 U1572 ( .IN1(n1897), .IN2(n1948), .IN3(n1947), .Q(
        \i_m4stg_frac/pcout_dff/N58 ) );
  XOR2X1 U1573 ( .IN1(\i_m4stg_frac/n360 ), .IN2(\i_m4stg_frac/n514 ), .Q(
        n1948) );
  AND2X1 U1574 ( .IN1(n1897), .IN2(n1949), .Q(\i_m4stg_frac/pcout_dff/N57 ) );
  NOR3X0 U1575 ( .IN1(n1952), .IN2(n1947), .IN3(n1951), .QN(n1949) );
  AND2X1 U1576 ( .IN1(\i_m4stg_frac/n362 ), .IN2(\i_m4stg_frac/n516 ), .Q(
        n1951) );
  NOR2X0 U1577 ( .IN1(\i_m4stg_frac/n516 ), .IN2(\i_m4stg_frac/n362 ), .QN(
        n1947) );
  OA22X1 U1578 ( .IN1(n2074), .IN2(\i_m4stg_frac/n364 ), .IN3(n2075), .IN4(
        \i_m4stg_frac/n518 ), .Q(n1952) );
  AND2X1 U1579 ( .IN1(\i_m4stg_frac/n364 ), .IN2(n2074), .Q(n2075) );
  AND3X1 U1580 ( .IN1(n1897), .IN2(n1954), .IN3(n1958), .Q(
        \i_m4stg_frac/pcout_dff/N56 ) );
  XNOR3X1 U1581 ( .IN1(\i_m4stg_frac/n518 ), .IN2(\i_m4stg_frac/n364 ), .IN3(
        n2074), .Q(n1954) );
  INVX0 U1582 ( .INP(n2076), .ZN(n2074) );
  NOR2X0 U1583 ( .IN1(n1375), .IN2(n1956), .QN(\i_m4stg_frac/pcout_dff/N55 )
         );
  NAND3X0 U1584 ( .IN1(n2077), .IN2(n1955), .IN3(n1965), .QN(n1956) );
  INVX0 U1585 ( .INP(n1958), .ZN(n1955) );
  NOR2X0 U1586 ( .IN1(n1962), .IN2(n1961), .QN(n1958) );
  NAND2X0 U1587 ( .IN1(n1961), .IN2(n1962), .QN(n2077) );
  AO22X1 U1588 ( .IN1(\i_m4stg_frac/n368 ), .IN2(n2078), .IN3(
        \i_m4stg_frac/n522 ), .IN4(n2079), .Q(n1962) );
  OR2X1 U1589 ( .IN1(\i_m4stg_frac/n368 ), .IN2(n2078), .Q(n2079) );
  AO21X1 U1590 ( .IN1(\i_m4stg_frac/n520 ), .IN2(\i_m4stg_frac/n366 ), .IN3(
        n2076), .Q(n1961) );
  NOR2X0 U1591 ( .IN1(\i_m4stg_frac/n520 ), .IN2(\i_m4stg_frac/n366 ), .QN(
        n2076) );
  NOR2X0 U1592 ( .IN1(n1374), .IN2(n1963), .QN(\i_m4stg_frac/pcout_dff/N54 )
         );
  NAND3X0 U1593 ( .IN1(n2080), .IN2(n1960), .IN3(n1972), .QN(n1963) );
  INVX0 U1594 ( .INP(n1965), .ZN(n1960) );
  NOR2X0 U1595 ( .IN1(n1968), .IN2(n1969), .QN(n1965) );
  NAND2X0 U1596 ( .IN1(n1969), .IN2(n1968), .QN(n2080) );
  AO22X1 U1597 ( .IN1(n2081), .IN2(n2082), .IN3(\i_m4stg_frac/n683 ), .IN4(
        n2083), .Q(n1968) );
  OR2X1 U1598 ( .IN1(n2082), .IN2(n2081), .Q(n2083) );
  XOR3X1 U1599 ( .IN1(\i_m4stg_frac/n522 ), .IN2(\i_m4stg_frac/n368 ), .IN3(
        n2078), .Q(n1969) );
  OA22X1 U1600 ( .IN1(\i_m4stg_frac/n370 ), .IN2(\i_m4stg_frac/n524 ), .IN3(
        n2084), .IN4(\i_m4stg_frac/n837 ), .Q(n2078) );
  AND2X1 U1601 ( .IN1(\i_m4stg_frac/n524 ), .IN2(\i_m4stg_frac/n370 ), .Q(
        n2084) );
  NOR2X0 U1602 ( .IN1(n1373), .IN2(n1970), .QN(\i_m4stg_frac/pcout_dff/N53 )
         );
  NAND3X0 U1603 ( .IN1(n2085), .IN2(n1967), .IN3(n1979), .QN(n1970) );
  INVX0 U1604 ( .INP(n1972), .ZN(n1967) );
  NOR2X0 U1605 ( .IN1(n1975), .IN2(n1976), .QN(n1972) );
  NAND2X0 U1606 ( .IN1(n1976), .IN2(n1975), .QN(n2085) );
  AO22X1 U1607 ( .IN1(n2086), .IN2(n2087), .IN3(\i_m4stg_frac/n685 ), .IN4(
        n2088), .Q(n1975) );
  OR2X1 U1608 ( .IN1(n2087), .IN2(n2086), .Q(n2088) );
  XOR3X1 U1609 ( .IN1(\i_m4stg_frac/n683 ), .IN2(n2081), .IN3(n2082), .Q(n1976) );
  XOR3X1 U1610 ( .IN1(\i_m4stg_frac/n837 ), .IN2(\i_m4stg_frac/n524 ), .IN3(
        \i_m4stg_frac/n370 ), .Q(n2082) );
  OA22X1 U1611 ( .IN1(\i_m4stg_frac/n372 ), .IN2(\i_m4stg_frac/n526 ), .IN3(
        n2089), .IN4(\i_m4stg_frac/n839 ), .Q(n2081) );
  AND2X1 U1612 ( .IN1(\i_m4stg_frac/n526 ), .IN2(\i_m4stg_frac/n372 ), .Q(
        n2089) );
  NOR2X0 U1613 ( .IN1(n1376), .IN2(n1977), .QN(\i_m4stg_frac/pcout_dff/N52 )
         );
  NAND3X0 U1614 ( .IN1(n2090), .IN2(n1974), .IN3(n1986), .QN(n1977) );
  INVX0 U1615 ( .INP(n1979), .ZN(n1974) );
  NOR2X0 U1616 ( .IN1(n1982), .IN2(n1983), .QN(n1979) );
  NAND2X0 U1617 ( .IN1(n1983), .IN2(n1982), .QN(n2090) );
  AO22X1 U1618 ( .IN1(n2091), .IN2(n2092), .IN3(\i_m4stg_frac/n687 ), .IN4(
        n2093), .Q(n1982) );
  OR2X1 U1619 ( .IN1(n2092), .IN2(n2091), .Q(n2093) );
  XOR3X1 U1620 ( .IN1(\i_m4stg_frac/n685 ), .IN2(n2086), .IN3(n2087), .Q(n1983) );
  XOR3X1 U1621 ( .IN1(\i_m4stg_frac/n839 ), .IN2(\i_m4stg_frac/n526 ), .IN3(
        \i_m4stg_frac/n372 ), .Q(n2087) );
  OA22X1 U1622 ( .IN1(\i_m4stg_frac/n374 ), .IN2(\i_m4stg_frac/n528 ), .IN3(
        n2094), .IN4(\i_m4stg_frac/n841 ), .Q(n2086) );
  AND2X1 U1623 ( .IN1(\i_m4stg_frac/n528 ), .IN2(\i_m4stg_frac/n374 ), .Q(
        n2094) );
  NOR2X0 U1624 ( .IN1(n1375), .IN2(n1984), .QN(\i_m4stg_frac/pcout_dff/N51 )
         );
  NAND3X0 U1625 ( .IN1(n2095), .IN2(n1981), .IN3(n1994), .QN(n1984) );
  INVX0 U1626 ( .INP(n1986), .ZN(n1981) );
  NOR2X0 U1627 ( .IN1(n1989), .IN2(n1990), .QN(n1986) );
  NAND2X0 U1628 ( .IN1(n1990), .IN2(n1989), .QN(n2095) );
  AO22X1 U1629 ( .IN1(n2096), .IN2(n2097), .IN3(\i_m4stg_frac/n689 ), .IN4(
        n2098), .Q(n1989) );
  OR2X1 U1630 ( .IN1(n2097), .IN2(n2096), .Q(n2098) );
  XOR3X1 U1631 ( .IN1(\i_m4stg_frac/n687 ), .IN2(n2091), .IN3(n2092), .Q(n1990) );
  XOR3X1 U1632 ( .IN1(\i_m4stg_frac/n841 ), .IN2(\i_m4stg_frac/n528 ), .IN3(
        \i_m4stg_frac/n374 ), .Q(n2092) );
  OA22X1 U1633 ( .IN1(\i_m4stg_frac/n376 ), .IN2(\i_m4stg_frac/n530 ), .IN3(
        n2099), .IN4(\i_m4stg_frac/n843 ), .Q(n2091) );
  AND2X1 U1634 ( .IN1(\i_m4stg_frac/n530 ), .IN2(\i_m4stg_frac/n376 ), .Q(
        n2099) );
  NOR2X0 U1635 ( .IN1(n1374), .IN2(n1992), .QN(\i_m4stg_frac/pcout_dff/N50 )
         );
  NAND3X0 U1636 ( .IN1(n2100), .IN2(n1988), .IN3(n2001), .QN(n1992) );
  INVX0 U1637 ( .INP(n1994), .ZN(n1988) );
  NOR2X0 U1638 ( .IN1(n1997), .IN2(n1998), .QN(n1994) );
  NAND2X0 U1639 ( .IN1(n1998), .IN2(n1997), .QN(n2100) );
  AO22X1 U1640 ( .IN1(n2101), .IN2(n2102), .IN3(\i_m4stg_frac/n691 ), .IN4(
        n2103), .Q(n1997) );
  OR2X1 U1641 ( .IN1(n2102), .IN2(n2101), .Q(n2103) );
  XOR3X1 U1642 ( .IN1(\i_m4stg_frac/n689 ), .IN2(n2096), .IN3(n2097), .Q(n1998) );
  XOR3X1 U1643 ( .IN1(\i_m4stg_frac/n843 ), .IN2(\i_m4stg_frac/n530 ), .IN3(
        \i_m4stg_frac/n376 ), .Q(n2097) );
  OA22X1 U1644 ( .IN1(\i_m4stg_frac/n378 ), .IN2(\i_m4stg_frac/n532 ), .IN3(
        n2104), .IN4(\i_m4stg_frac/n845 ), .Q(n2096) );
  AND2X1 U1645 ( .IN1(\i_m4stg_frac/n532 ), .IN2(\i_m4stg_frac/n378 ), .Q(
        n2104) );
  NOR3X0 U1646 ( .IN1(n2105), .IN2(n1376), .IN3(n2106), .QN(
        \i_m4stg_frac/pcout_dff/N5 ) );
  NOR2X0 U1647 ( .IN1(n1373), .IN2(n1999), .QN(\i_m4stg_frac/pcout_dff/N49 )
         );
  NAND3X0 U1648 ( .IN1(n2107), .IN2(n1996), .IN3(n2008), .QN(n1999) );
  INVX0 U1649 ( .INP(n2001), .ZN(n1996) );
  NOR2X0 U1650 ( .IN1(n2004), .IN2(n2005), .QN(n2001) );
  NAND2X0 U1651 ( .IN1(n2005), .IN2(n2004), .QN(n2107) );
  AO22X1 U1652 ( .IN1(n2108), .IN2(n2109), .IN3(\i_m4stg_frac/n693 ), .IN4(
        n2110), .Q(n2004) );
  OR2X1 U1653 ( .IN1(n2109), .IN2(n2108), .Q(n2110) );
  XOR3X1 U1654 ( .IN1(\i_m4stg_frac/n691 ), .IN2(n2101), .IN3(n2102), .Q(n2005) );
  XOR3X1 U1655 ( .IN1(\i_m4stg_frac/n845 ), .IN2(\i_m4stg_frac/n532 ), .IN3(
        \i_m4stg_frac/n378 ), .Q(n2102) );
  OA22X1 U1656 ( .IN1(\i_m4stg_frac/n380 ), .IN2(\i_m4stg_frac/n534 ), .IN3(
        n2111), .IN4(\i_m4stg_frac/n847 ), .Q(n2101) );
  AND2X1 U1657 ( .IN1(\i_m4stg_frac/n534 ), .IN2(\i_m4stg_frac/n380 ), .Q(
        n2111) );
  NOR2X0 U1658 ( .IN1(n1376), .IN2(n2006), .QN(\i_m4stg_frac/pcout_dff/N48 )
         );
  NAND3X0 U1659 ( .IN1(n2112), .IN2(n2003), .IN3(n2015), .QN(n2006) );
  INVX0 U1660 ( .INP(n2008), .ZN(n2003) );
  NOR2X0 U1661 ( .IN1(n2011), .IN2(n2012), .QN(n2008) );
  NAND2X0 U1662 ( .IN1(n2012), .IN2(n2011), .QN(n2112) );
  AO22X1 U1663 ( .IN1(n2113), .IN2(n2114), .IN3(\i_m4stg_frac/n695 ), .IN4(
        n2115), .Q(n2011) );
  OR2X1 U1664 ( .IN1(n2114), .IN2(n2113), .Q(n2115) );
  XOR3X1 U1665 ( .IN1(\i_m4stg_frac/n693 ), .IN2(n2108), .IN3(n2109), .Q(n2012) );
  XOR3X1 U1666 ( .IN1(\i_m4stg_frac/n847 ), .IN2(\i_m4stg_frac/n534 ), .IN3(
        \i_m4stg_frac/n380 ), .Q(n2109) );
  OA22X1 U1667 ( .IN1(\i_m4stg_frac/n382 ), .IN2(\i_m4stg_frac/n536 ), .IN3(
        n2116), .IN4(\i_m4stg_frac/n849 ), .Q(n2108) );
  AND2X1 U1668 ( .IN1(\i_m4stg_frac/n536 ), .IN2(\i_m4stg_frac/n382 ), .Q(
        n2116) );
  NOR2X0 U1669 ( .IN1(n1375), .IN2(n2013), .QN(\i_m4stg_frac/pcout_dff/N47 )
         );
  NAND3X0 U1670 ( .IN1(n2117), .IN2(n2010), .IN3(n2118), .QN(n2013) );
  INVX0 U1671 ( .INP(n2015), .ZN(n2010) );
  NOR2X0 U1672 ( .IN1(n2018), .IN2(n2019), .QN(n2015) );
  NAND2X0 U1673 ( .IN1(n2019), .IN2(n2018), .QN(n2117) );
  AO22X1 U1674 ( .IN1(n2119), .IN2(n2120), .IN3(\i_m4stg_frac/n697 ), .IN4(
        n2121), .Q(n2018) );
  OR2X1 U1675 ( .IN1(n2120), .IN2(n2119), .Q(n2121) );
  XOR3X1 U1676 ( .IN1(\i_m4stg_frac/n695 ), .IN2(n2113), .IN3(n2114), .Q(n2019) );
  XOR3X1 U1677 ( .IN1(\i_m4stg_frac/n849 ), .IN2(\i_m4stg_frac/n536 ), .IN3(
        \i_m4stg_frac/n382 ), .Q(n2114) );
  OA22X1 U1678 ( .IN1(\i_m4stg_frac/n384 ), .IN2(\i_m4stg_frac/n538 ), .IN3(
        n2122), .IN4(\i_m4stg_frac/n851 ), .Q(n2113) );
  AND2X1 U1679 ( .IN1(\i_m4stg_frac/n538 ), .IN2(\i_m4stg_frac/n384 ), .Q(
        n2122) );
  NOR2X0 U1680 ( .IN1(n1374), .IN2(n2123), .QN(\i_m4stg_frac/pcout_dff/N46 )
         );
  NOR2X0 U1681 ( .IN1(n1373), .IN2(n2124), .QN(\i_m4stg_frac/pcout_dff/N45 )
         );
  NOR2X0 U1682 ( .IN1(n1376), .IN2(n2125), .QN(\i_m4stg_frac/pcout_dff/N44 )
         );
  NOR3X0 U1683 ( .IN1(n2126), .IN2(n1375), .IN3(n2127), .QN(
        \i_m4stg_frac/pcout_dff/N43 ) );
  NOR2X0 U1684 ( .IN1(n1375), .IN2(n2128), .QN(\i_m4stg_frac/pcout_dff/N42 )
         );
  AND3X1 U1685 ( .IN1(n2129), .IN2(n1897), .IN3(n2130), .Q(
        \i_m4stg_frac/pcout_dff/N41 ) );
  NOR3X0 U1686 ( .IN1(n1373), .IN2(n2131), .IN3(n2132), .QN(
        \i_m4stg_frac/pcout_dff/N40 ) );
  NOR3X0 U1687 ( .IN1(n2133), .IN2(n1374), .IN3(n2134), .QN(
        \i_m4stg_frac/pcout_dff/N4 ) );
  NOR3X0 U1688 ( .IN1(n2135), .IN2(n1373), .IN3(n2136), .QN(
        \i_m4stg_frac/pcout_dff/N39 ) );
  NOR3X0 U1689 ( .IN1(n2137), .IN2(n1376), .IN3(n2138), .QN(
        \i_m4stg_frac/pcout_dff/N38 ) );
  NOR3X0 U1690 ( .IN1(n2139), .IN2(n1375), .IN3(n2140), .QN(
        \i_m4stg_frac/pcout_dff/N37 ) );
  NOR3X0 U1691 ( .IN1(n2141), .IN2(n1374), .IN3(n2142), .QN(
        \i_m4stg_frac/pcout_dff/N36 ) );
  NOR3X0 U1692 ( .IN1(n2143), .IN2(n1373), .IN3(n2144), .QN(
        \i_m4stg_frac/pcout_dff/N35 ) );
  NOR3X0 U1693 ( .IN1(n2145), .IN2(n1376), .IN3(n2146), .QN(
        \i_m4stg_frac/pcout_dff/N34 ) );
  NOR3X0 U1694 ( .IN1(n2147), .IN2(n1375), .IN3(n2148), .QN(
        \i_m4stg_frac/pcout_dff/N33 ) );
  NOR3X0 U1695 ( .IN1(n2149), .IN2(n1374), .IN3(n2150), .QN(
        \i_m4stg_frac/pcout_dff/N32 ) );
  NOR3X0 U1696 ( .IN1(n2151), .IN2(n1373), .IN3(n2152), .QN(
        \i_m4stg_frac/pcout_dff/N31 ) );
  NOR3X0 U1697 ( .IN1(n2153), .IN2(n1376), .IN3(n2154), .QN(
        \i_m4stg_frac/pcout_dff/N30 ) );
  NOR3X0 U1698 ( .IN1(n2155), .IN2(n1375), .IN3(n2156), .QN(
        \i_m4stg_frac/pcout_dff/N29 ) );
  NOR3X0 U1699 ( .IN1(n2157), .IN2(n1374), .IN3(n2158), .QN(
        \i_m4stg_frac/pcout_dff/N28 ) );
  NOR3X0 U1700 ( .IN1(n2159), .IN2(n1373), .IN3(n2160), .QN(
        \i_m4stg_frac/pcout_dff/N27 ) );
  NOR3X0 U1701 ( .IN1(n2161), .IN2(n1376), .IN3(n2162), .QN(
        \i_m4stg_frac/pcout_dff/N26 ) );
  NOR3X0 U1702 ( .IN1(n2163), .IN2(n1375), .IN3(n2164), .QN(
        \i_m4stg_frac/pcout_dff/N25 ) );
  NOR3X0 U1703 ( .IN1(n2165), .IN2(n1374), .IN3(n2166), .QN(
        \i_m4stg_frac/pcout_dff/N24 ) );
  NOR3X0 U1704 ( .IN1(n2167), .IN2(n1373), .IN3(n2168), .QN(
        \i_m4stg_frac/pcout_dff/N23 ) );
  NOR3X0 U1705 ( .IN1(n2169), .IN2(n1376), .IN3(n2170), .QN(
        \i_m4stg_frac/pcout_dff/N22 ) );
  NOR3X0 U1706 ( .IN1(n2171), .IN2(n1375), .IN3(n2172), .QN(
        \i_m4stg_frac/pcout_dff/N21 ) );
  NOR3X0 U1707 ( .IN1(n2173), .IN2(n1374), .IN3(n2174), .QN(
        \i_m4stg_frac/pcout_dff/N20 ) );
  NOR3X0 U1708 ( .IN1(n2175), .IN2(n1373), .IN3(n2176), .QN(
        \i_m4stg_frac/pcout_dff/N19 ) );
  NOR3X0 U1709 ( .IN1(n2177), .IN2(n1376), .IN3(n2178), .QN(
        \i_m4stg_frac/pcout_dff/N18 ) );
  NOR3X0 U1710 ( .IN1(n2179), .IN2(n1375), .IN3(n2180), .QN(
        \i_m4stg_frac/pcout_dff/N17 ) );
  NOR3X0 U1711 ( .IN1(n2181), .IN2(n1374), .IN3(n2182), .QN(
        \i_m4stg_frac/pcout_dff/N16 ) );
  NOR3X0 U1712 ( .IN1(n2183), .IN2(n1373), .IN3(n2184), .QN(
        \i_m4stg_frac/pcout_dff/N15 ) );
  NOR3X0 U1713 ( .IN1(n2185), .IN2(n1376), .IN3(n2186), .QN(
        \i_m4stg_frac/pcout_dff/N14 ) );
  NOR3X0 U1714 ( .IN1(n2187), .IN2(n1375), .IN3(n2188), .QN(
        \i_m4stg_frac/pcout_dff/N13 ) );
  NOR3X0 U1715 ( .IN1(n2189), .IN2(n1374), .IN3(n2190), .QN(
        \i_m4stg_frac/pcout_dff/N12 ) );
  AND3X1 U1716 ( .IN1(n2191), .IN2(n1897), .IN3(n2192), .Q(
        \i_m4stg_frac/pcout_dff/N11 ) );
  INVX0 U1717 ( .INP(n2193), .ZN(n2191) );
  AND3X1 U1718 ( .IN1(n2194), .IN2(n2195), .IN3(n1897), .Q(
        \i_m4stg_frac/pcout_dff/N10 ) );
  INVX0 U1719 ( .INP(n1375), .ZN(n1897) );
  INVX0 U1720 ( .INP(n2196), .ZN(n2194) );
  AND3X1 U1721 ( .IN1(n2197), .IN2(n1536), .IN3(n2198), .Q(\i_m4stg_frac/n637 ) );
  NOR3X0 U1722 ( .IN1(n2199), .IN2(se_mul64), .IN3(n2200), .QN(
        \i_m4stg_frac/n635 ) );
  AND3X1 U1723 ( .IN1(n2201), .IN2(\i_m4stg_frac/n854 ), .IN3(n2202), .Q(
        \i_m4stg_frac/n633 ) );
  OAI21X1 U1724 ( .IN1(n2203), .IN2(n2204), .IN3(n2205), .QN(n2201) );
  AND2X1 U1725 ( .IN1(n2206), .IN2(n2207), .Q(n2204) );
  NOR2X0 U1726 ( .IN1(se_mul64), .IN2(n2208), .QN(\i_m4stg_frac/n631 ) );
  XOR2X1 U1727 ( .IN1(n2203), .IN2(n2209), .Q(n2208) );
  NOR2X0 U1728 ( .IN1(se_mul64), .IN2(n2023), .QN(\i_m4stg_frac/n629 ) );
  XNOR2X1 U1729 ( .IN1(n2127), .IN2(n2126), .Q(n2023) );
  NOR2X0 U1730 ( .IN1(se_mul64), .IN2(n2022), .QN(\i_m4stg_frac/n627 ) );
  NAND2X0 U1731 ( .IN1(n2210), .IN2(n2125), .QN(n2022) );
  AO22X1 U1732 ( .IN1(n2211), .IN2(n2212), .IN3(n2213), .IN4(n2214), .Q(n2210)
         );
  NOR2X0 U1733 ( .IN1(se_mul64), .IN2(n2021), .QN(\i_m4stg_frac/n625 ) );
  AO21X1 U1734 ( .IN1(n2214), .IN2(n2215), .IN3(n2216), .Q(n2021) );
  INVX0 U1735 ( .INP(n2124), .ZN(n2216) );
  AO21X1 U1736 ( .IN1(n2217), .IN2(n2218), .IN3(n2219), .Q(n2215) );
  NOR2X0 U1737 ( .IN1(se_mul64), .IN2(n2020), .QN(\i_m4stg_frac/n623 ) );
  AO21X1 U1738 ( .IN1(n2220), .IN2(n2221), .IN3(n2222), .Q(n2020) );
  INVX0 U1739 ( .INP(n2123), .ZN(n2222) );
  NAND3X0 U1740 ( .IN1(n2223), .IN2(n2017), .IN3(n2219), .QN(n2123) );
  INVX0 U1741 ( .INP(n2118), .ZN(n2017) );
  NAND2X0 U1742 ( .IN1(n2224), .IN2(n2225), .QN(n2223) );
  AO21X1 U1743 ( .IN1(n2224), .IN2(n2225), .IN3(n2118), .Q(n2221) );
  NOR2X0 U1744 ( .IN1(n2225), .IN2(n2224), .QN(n2118) );
  AO22X1 U1745 ( .IN1(n2226), .IN2(n2227), .IN3(\i_m4stg_frac/n699 ), .IN4(
        n2228), .Q(n2225) );
  OR2X1 U1746 ( .IN1(n2227), .IN2(n2226), .Q(n2228) );
  XOR3X1 U1747 ( .IN1(\i_m4stg_frac/n697 ), .IN2(n2119), .IN3(n2120), .Q(n2224) );
  XOR3X1 U1748 ( .IN1(\i_m4stg_frac/n851 ), .IN2(\i_m4stg_frac/n538 ), .IN3(
        \i_m4stg_frac/n384 ), .Q(n2120) );
  OA22X1 U1749 ( .IN1(\i_m4stg_frac/n386 ), .IN2(\i_m4stg_frac/n540 ), .IN3(
        n2229), .IN4(\i_m4stg_frac/n853 ), .Q(n2119) );
  AND2X1 U1750 ( .IN1(\i_m4stg_frac/n540 ), .IN2(\i_m4stg_frac/n386 ), .Q(
        n2229) );
  AND3X1 U1751 ( .IN1(n2230), .IN2(n1535), .IN3(n2231), .Q(\i_m4stg_frac/n621 ) );
  NOR2X0 U1752 ( .IN1(se_mul64), .IN2(n2232), .QN(\i_m4stg_frac/n619 ) );
  XOR3X1 U1753 ( .IN1(\i_m4stg_frac/ps[32] ), .IN2(\i_m4stg_frac/pc[31] ), 
        .IN3(\i_m4stg_frac/n997 ), .Q(n2232) );
  AND3X1 U1754 ( .IN1(n2233), .IN2(\i_m4stg_frac/n854 ), .IN3(n2234), .Q(
        \i_m4stg_frac/n617 ) );
  OR2X1 U1755 ( .IN1(n2235), .IN2(n2236), .Q(n2233) );
  NOR2X0 U1756 ( .IN1(se_mul64), .IN2(n2237), .QN(\i_m4stg_frac/n615 ) );
  XNOR2X1 U1757 ( .IN1(n2234), .IN2(n2238), .Q(n2237) );
  AND3X1 U1758 ( .IN1(n2239), .IN2(\i_m4stg_frac/n854 ), .IN3(n2240), .Q(
        \i_m4stg_frac/n613 ) );
  AO22X1 U1759 ( .IN1(n2205), .IN2(n2241), .IN3(n2242), .IN4(n2243), .Q(n2239)
         );
  NOR2X0 U1760 ( .IN1(se_mul64), .IN2(n2244), .QN(\i_m4stg_frac/n611 ) );
  XNOR3X1 U1761 ( .IN1(n2245), .IN2(n2246), .IN3(n2247), .Q(n2244) );
  NOR2X0 U1762 ( .IN1(se_mul64), .IN2(n2248), .QN(\i_m4stg_frac/n609 ) );
  XNOR2X1 U1763 ( .IN1(n2249), .IN2(n2250), .Q(n2248) );
  NOR3X0 U1764 ( .IN1(n2251), .IN2(se_mul64), .IN3(n2252), .QN(
        \i_m4stg_frac/n607 ) );
  NOR3X0 U1765 ( .IN1(n2253), .IN2(se_mul64), .IN3(n2254), .QN(
        \i_m4stg_frac/n605 ) );
  NOR3X0 U1766 ( .IN1(n2255), .IN2(se_mul64), .IN3(n2256), .QN(
        \i_m4stg_frac/n603 ) );
  NOR3X0 U1767 ( .IN1(n2257), .IN2(se_mul64), .IN3(n2258), .QN(
        \i_m4stg_frac/n601 ) );
  NOR3X0 U1768 ( .IN1(n2259), .IN2(se_mul64), .IN3(n2260), .QN(
        \i_m4stg_frac/n599 ) );
  NOR3X0 U1769 ( .IN1(n2261), .IN2(se_mul64), .IN3(n2262), .QN(
        \i_m4stg_frac/n597 ) );
  NOR3X0 U1770 ( .IN1(n2263), .IN2(se_mul64), .IN3(n2264), .QN(
        \i_m4stg_frac/n595 ) );
  NOR3X0 U1771 ( .IN1(n2265), .IN2(se_mul64), .IN3(n2266), .QN(
        \i_m4stg_frac/n593 ) );
  NOR3X0 U1772 ( .IN1(n2267), .IN2(se_mul64), .IN3(n2268), .QN(
        \i_m4stg_frac/n591 ) );
  NOR3X0 U1773 ( .IN1(n2269), .IN2(se_mul64), .IN3(n2270), .QN(
        \i_m4stg_frac/n589 ) );
  NOR3X0 U1774 ( .IN1(n2271), .IN2(se_mul64), .IN3(n2272), .QN(
        \i_m4stg_frac/n587 ) );
  NOR3X0 U1775 ( .IN1(n2273), .IN2(se_mul64), .IN3(n2274), .QN(
        \i_m4stg_frac/n585 ) );
  NOR3X0 U1776 ( .IN1(n2275), .IN2(se_mul64), .IN3(n2276), .QN(
        \i_m4stg_frac/n583 ) );
  NOR3X0 U1777 ( .IN1(n2277), .IN2(se_mul64), .IN3(n2278), .QN(
        \i_m4stg_frac/n581 ) );
  NOR3X0 U1778 ( .IN1(n2279), .IN2(se_mul64), .IN3(n2280), .QN(
        \i_m4stg_frac/n579 ) );
  NOR3X0 U1779 ( .IN1(n2281), .IN2(se_mul64), .IN3(n2282), .QN(
        \i_m4stg_frac/n577 ) );
  NOR3X0 U1780 ( .IN1(n2283), .IN2(se_mul64), .IN3(n2284), .QN(
        \i_m4stg_frac/n575 ) );
  NOR3X0 U1781 ( .IN1(n2285), .IN2(se_mul64), .IN3(n2286), .QN(
        \i_m4stg_frac/n573 ) );
  NOR3X0 U1782 ( .IN1(n2134), .IN2(se_mul64), .IN3(n2133), .QN(
        \i_m4stg_frac/n571 ) );
  NOR3X0 U1783 ( .IN1(n2106), .IN2(se_mul64), .IN3(n2105), .QN(
        \i_m4stg_frac/n569 ) );
  NOR3X0 U1784 ( .IN1(n2073), .IN2(se_mul64), .IN3(n2072), .QN(
        \i_m4stg_frac/n567 ) );
  NOR3X0 U1785 ( .IN1(n2062), .IN2(se_mul64), .IN3(n2061), .QN(
        \i_m4stg_frac/n565 ) );
  NOR3X0 U1786 ( .IN1(n2060), .IN2(se_mul64), .IN3(n2059), .QN(
        \i_m4stg_frac/n563 ) );
  NOR3X0 U1787 ( .IN1(n2058), .IN2(se_mul64), .IN3(n2057), .QN(
        \i_m4stg_frac/n561 ) );
  NOR3X0 U1788 ( .IN1(n2287), .IN2(se_mul64), .IN3(n2196), .QN(
        \i_m4stg_frac/n559 ) );
  NOR3X0 U1789 ( .IN1(n2288), .IN2(se_mul64), .IN3(n2193), .QN(
        \i_m4stg_frac/n557 ) );
  NOR3X0 U1790 ( .IN1(n2190), .IN2(se_mul64), .IN3(n2189), .QN(
        \i_m4stg_frac/n555 ) );
  NOR3X0 U1791 ( .IN1(n2188), .IN2(se_mul64), .IN3(n2187), .QN(
        \i_m4stg_frac/n553 ) );
  NOR3X0 U1792 ( .IN1(n2186), .IN2(se_mul64), .IN3(n2185), .QN(
        \i_m4stg_frac/n551 ) );
  NOR3X0 U1793 ( .IN1(n2184), .IN2(se_mul64), .IN3(n2183), .QN(
        \i_m4stg_frac/n549 ) );
  NOR3X0 U1794 ( .IN1(n2182), .IN2(se_mul64), .IN3(n2181), .QN(
        \i_m4stg_frac/n547 ) );
  NOR3X0 U1795 ( .IN1(n2180), .IN2(se_mul64), .IN3(n2179), .QN(
        \i_m4stg_frac/n545 ) );
  NOR3X0 U1796 ( .IN1(n2178), .IN2(se_mul64), .IN3(n2177), .QN(
        \i_m4stg_frac/n543 ) );
  NOR3X0 U1797 ( .IN1(n2176), .IN2(se_mul64), .IN3(n2175), .QN(
        \i_m4stg_frac/n541 ) );
  NOR3X0 U1798 ( .IN1(n2174), .IN2(se_mul64), .IN3(n2173), .QN(
        \i_m4stg_frac/n539 ) );
  NOR3X0 U1799 ( .IN1(n2172), .IN2(se_mul64), .IN3(n2171), .QN(
        \i_m4stg_frac/n537 ) );
  NOR3X0 U1800 ( .IN1(n2170), .IN2(se_mul64), .IN3(n2169), .QN(
        \i_m4stg_frac/n535 ) );
  NOR3X0 U1801 ( .IN1(n2168), .IN2(se_mul64), .IN3(n2167), .QN(
        \i_m4stg_frac/n533 ) );
  NOR3X0 U1802 ( .IN1(n2166), .IN2(se_mul64), .IN3(n2165), .QN(
        \i_m4stg_frac/n531 ) );
  NOR3X0 U1803 ( .IN1(n2164), .IN2(se_mul64), .IN3(n2163), .QN(
        \i_m4stg_frac/n529 ) );
  NOR3X0 U1804 ( .IN1(n2162), .IN2(se_mul64), .IN3(n2161), .QN(
        \i_m4stg_frac/n527 ) );
  NOR3X0 U1805 ( .IN1(n2160), .IN2(se_mul64), .IN3(n2159), .QN(
        \i_m4stg_frac/n525 ) );
  NOR3X0 U1806 ( .IN1(n2158), .IN2(se_mul64), .IN3(n2157), .QN(
        \i_m4stg_frac/n523 ) );
  NOR3X0 U1807 ( .IN1(n2156), .IN2(se_mul64), .IN3(n2155), .QN(
        \i_m4stg_frac/n521 ) );
  NOR3X0 U1808 ( .IN1(n2154), .IN2(se_mul64), .IN3(n2153), .QN(
        \i_m4stg_frac/n519 ) );
  NOR3X0 U1809 ( .IN1(n2152), .IN2(se_mul64), .IN3(n2151), .QN(
        \i_m4stg_frac/n517 ) );
  NOR3X0 U1810 ( .IN1(n2150), .IN2(se_mul64), .IN3(n2149), .QN(
        \i_m4stg_frac/n515 ) );
  NOR3X0 U1811 ( .IN1(n2148), .IN2(se_mul64), .IN3(n2147), .QN(
        \i_m4stg_frac/n513 ) );
  NOR3X0 U1812 ( .IN1(n2146), .IN2(se_mul64), .IN3(n2145), .QN(
        \i_m4stg_frac/n511 ) );
  NOR3X0 U1813 ( .IN1(n2144), .IN2(se_mul64), .IN3(n2143), .QN(
        \i_m4stg_frac/n509 ) );
  NOR3X0 U1814 ( .IN1(n2142), .IN2(se_mul64), .IN3(n2141), .QN(
        \i_m4stg_frac/n507 ) );
  NOR3X0 U1815 ( .IN1(n2140), .IN2(se_mul64), .IN3(n2139), .QN(
        \i_m4stg_frac/n505 ) );
  NOR3X0 U1816 ( .IN1(n2138), .IN2(se_mul64), .IN3(n2137), .QN(
        \i_m4stg_frac/n503 ) );
  NOR3X0 U1817 ( .IN1(n2136), .IN2(se_mul64), .IN3(n2135), .QN(
        \i_m4stg_frac/n501 ) );
  NOR3X0 U1818 ( .IN1(n2132), .IN2(se_mul64), .IN3(n2131), .QN(
        \i_m4stg_frac/n499 ) );
  NOR3X0 U1819 ( .IN1(n2289), .IN2(se_mul64), .IN3(n2290), .QN(
        \i_m4stg_frac/n497 ) );
  NOR2X0 U1820 ( .IN1(se_mul64), .IN2(n2128), .QN(\i_m4stg_frac/n495 ) );
  NOR3X0 U1821 ( .IN1(n2291), .IN2(se_mul64), .IN3(n2292), .QN(
        \i_m4stg_frac/n493 ) );
  NOR2X0 U1822 ( .IN1(se_mul64), .IN2(n2293), .QN(\i_m4stg_frac/n492 ) );
  XNOR2X1 U1823 ( .IN1(n2268), .IN2(n2267), .Q(n2293) );
  AO21X1 U1824 ( .IN1(n2294), .IN2(n2295), .IN3(n2250), .Q(n2267) );
  AO22X1 U1825 ( .IN1(n2296), .IN2(n2297), .IN3(n2298), .IN4(n2299), .Q(n2268)
         );
  OR2X1 U1826 ( .IN1(n2297), .IN2(n2296), .Q(n2299) );
  NOR2X0 U1827 ( .IN1(se_mul64), .IN2(n2300), .QN(\i_m4stg_frac/n491 ) );
  XNOR2X1 U1828 ( .IN1(n2291), .IN2(n2292), .Q(n2300) );
  XOR3X1 U1829 ( .IN1(\i_m4stg_frac/n831 ), .IN2(n2301), .IN3(n2302), .Q(n2292) );
  AO22X1 U1830 ( .IN1(n2303), .IN2(n2304), .IN3(\i_m4stg_frac/n833 ), .IN4(
        n2305), .Q(n2291) );
  NAND2X0 U1831 ( .IN1(n2306), .IN2(n2307), .QN(n2305) );
  INVX0 U1832 ( .INP(n2306), .ZN(n2304) );
  NOR2X0 U1833 ( .IN1(se_mul64), .IN2(n2308), .QN(\i_m4stg_frac/n489 ) );
  XNOR2X1 U1834 ( .IN1(n2230), .IN2(n2231), .Q(n2308) );
  XOR3X1 U1835 ( .IN1(n1188), .IN2(n2309), .IN3(n2310), .Q(n2231) );
  OA22X1 U1836 ( .IN1(n2301), .IN2(n2302), .IN3(n1329), .IN4(n2311), .Q(n2230)
         );
  AND2X1 U1837 ( .IN1(n2302), .IN2(n2301), .Q(n2311) );
  XNOR3X1 U1838 ( .IN1(\i_m4stg_frac/ps[38] ), .IN2(\i_m4stg_frac/pc[37] ), 
        .IN3(\i_m4stg_frac/n985 ), .Q(n2302) );
  AO22X1 U1839 ( .IN1(\i_m4stg_frac/pc[36] ), .IN2(n1073), .IN3(
        \i_m4stg_frac/ps[37] ), .IN4(n2312), .Q(n2301) );
  OR2X1 U1840 ( .IN1(n1073), .IN2(\i_m4stg_frac/pc[36] ), .Q(n2312) );
  NOR2X0 U1841 ( .IN1(se_mul64), .IN2(n2313), .QN(\i_m4stg_frac/n487 ) );
  XNOR2X1 U1842 ( .IN1(n2197), .IN2(n2198), .Q(n2313) );
  XNOR3X1 U1843 ( .IN1(\i_m4stg_frac/n827 ), .IN2(n2314), .IN3(n2315), .Q(
        n2198) );
  OA22X1 U1844 ( .IN1(n2309), .IN2(n2310), .IN3(n1188), .IN4(n2316), .Q(n2197)
         );
  AND2X1 U1845 ( .IN1(n2310), .IN2(n2309), .Q(n2316) );
  XOR3X1 U1846 ( .IN1(\i_m4stg_frac/ps[39] ), .IN2(\i_m4stg_frac/pc[38] ), 
        .IN3(n1068), .Q(n2310) );
  AO22X1 U1847 ( .IN1(\i_m4stg_frac/pc[37] ), .IN2(n1190), .IN3(
        \i_m4stg_frac/ps[38] ), .IN4(n2317), .Q(n2309) );
  OR2X1 U1848 ( .IN1(n1190), .IN2(\i_m4stg_frac/pc[37] ), .Q(n2317) );
  NOR2X0 U1849 ( .IN1(se_mul64), .IN2(n2318), .QN(\i_m4stg_frac/n485 ) );
  XNOR2X1 U1850 ( .IN1(n2253), .IN2(n2254), .Q(n2318) );
  XNOR3X1 U1851 ( .IN1(\i_m4stg_frac/n821 ), .IN2(n2319), .IN3(n2320), .Q(
        n2254) );
  AO22X1 U1852 ( .IN1(n2321), .IN2(n2322), .IN3(\i_m4stg_frac/n823 ), .IN4(
        n2323), .Q(n2253) );
  NAND2X0 U1853 ( .IN1(n2324), .IN2(n2325), .QN(n2323) );
  INVX0 U1854 ( .INP(n2324), .ZN(n2322) );
  NOR2X0 U1855 ( .IN1(se_mul64), .IN2(n2326), .QN(\i_m4stg_frac/n483 ) );
  XNOR2X1 U1856 ( .IN1(n2255), .IN2(n2256), .Q(n2326) );
  XNOR3X1 U1857 ( .IN1(\i_m4stg_frac/n819 ), .IN2(n2327), .IN3(n2328), .Q(
        n2256) );
  AO22X1 U1858 ( .IN1(n2319), .IN2(n2329), .IN3(\i_m4stg_frac/n821 ), .IN4(
        n2330), .Q(n2255) );
  NAND2X0 U1859 ( .IN1(n2320), .IN2(n2331), .QN(n2330) );
  INVX0 U1860 ( .INP(n2320), .ZN(n2329) );
  XOR3X1 U1861 ( .IN1(\i_m4stg_frac/ps[43] ), .IN2(\i_m4stg_frac/pc[42] ), 
        .IN3(n1060), .Q(n2320) );
  INVX0 U1862 ( .INP(n2331), .ZN(n2319) );
  AO22X1 U1863 ( .IN1(\i_m4stg_frac/pc[41] ), .IN2(n1069), .IN3(
        \i_m4stg_frac/ps[42] ), .IN4(n2332), .Q(n2331) );
  OR2X1 U1864 ( .IN1(n1069), .IN2(\i_m4stg_frac/pc[41] ), .Q(n2332) );
  NOR2X0 U1865 ( .IN1(se_mul64), .IN2(n2333), .QN(\i_m4stg_frac/n481 ) );
  XNOR2X1 U1866 ( .IN1(n2257), .IN2(n2258), .Q(n2333) );
  XNOR3X1 U1867 ( .IN1(\i_m4stg_frac/n817 ), .IN2(n2334), .IN3(n2335), .Q(
        n2258) );
  AO22X1 U1868 ( .IN1(n2327), .IN2(n2336), .IN3(\i_m4stg_frac/n819 ), .IN4(
        n2337), .Q(n2257) );
  NAND2X0 U1869 ( .IN1(n2328), .IN2(n2338), .QN(n2337) );
  INVX0 U1870 ( .INP(n2328), .ZN(n2336) );
  XOR3X1 U1871 ( .IN1(\i_m4stg_frac/ps[44] ), .IN2(\i_m4stg_frac/pc[43] ), 
        .IN3(n1072), .Q(n2328) );
  INVX0 U1872 ( .INP(n2338), .ZN(n2327) );
  AO22X1 U1873 ( .IN1(\i_m4stg_frac/pc[42] ), .IN2(n1060), .IN3(
        \i_m4stg_frac/ps[43] ), .IN4(n2339), .Q(n2338) );
  OR2X1 U1874 ( .IN1(n1060), .IN2(\i_m4stg_frac/pc[42] ), .Q(n2339) );
  NOR2X0 U1875 ( .IN1(se_mul64), .IN2(n2340), .QN(\i_m4stg_frac/n479 ) );
  XNOR2X1 U1876 ( .IN1(n2341), .IN2(n2342), .Q(n2340) );
  NOR2X0 U1877 ( .IN1(se_mul64), .IN2(n2343), .QN(\i_m4stg_frac/n477 ) );
  XNOR2X1 U1878 ( .IN1(n2261), .IN2(n2262), .Q(n2343) );
  XOR3X1 U1879 ( .IN1(n2344), .IN2(n2345), .IN3(n2346), .Q(n2262) );
  AO22X1 U1880 ( .IN1(n2347), .IN2(n2348), .IN3(n2349), .IN4(n2350), .Q(n2261)
         );
  NAND2X0 U1881 ( .IN1(n2351), .IN2(n2352), .QN(n2349) );
  INVX0 U1882 ( .INP(n2351), .ZN(n2348) );
  INVX0 U1883 ( .INP(n2352), .ZN(n2347) );
  NOR2X0 U1884 ( .IN1(se_mul64), .IN2(n2353), .QN(\i_m4stg_frac/n475 ) );
  XNOR2X1 U1885 ( .IN1(n2263), .IN2(n2264), .Q(n2353) );
  XOR3X1 U1886 ( .IN1(n2354), .IN2(n2355), .IN3(n2356), .Q(n2264) );
  AO22X1 U1887 ( .IN1(n2345), .IN2(n2346), .IN3(n2344), .IN4(n2357), .Q(n2263)
         );
  OR2X1 U1888 ( .IN1(n2346), .IN2(n2345), .Q(n2357) );
  XOR3X1 U1889 ( .IN1(\i_m4stg_frac/n963 ), .IN2(\i_m4stg_frac/n809 ), .IN3(
        n2358), .Q(n2344) );
  OA22X1 U1890 ( .IN1(n2359), .IN2(\i_m4stg_frac/n811 ), .IN3(n2360), .IN4(
        \i_m4stg_frac/n965 ), .Q(n2346) );
  AND2X1 U1891 ( .IN1(\i_m4stg_frac/n811 ), .IN2(n2359), .Q(n2360) );
  AOI22X1 U1892 ( .IN1(\i_m4stg_frac/pc[47] ), .IN2(n1199), .IN3(
        \i_m4stg_frac/ps[48] ), .IN4(n2361), .QN(n2345) );
  OR2X1 U1893 ( .IN1(n1199), .IN2(\i_m4stg_frac/pc[47] ), .Q(n2361) );
  NOR2X0 U1894 ( .IN1(se_mul64), .IN2(n2362), .QN(\i_m4stg_frac/n473 ) );
  XNOR2X1 U1895 ( .IN1(n2265), .IN2(n2266), .Q(n2362) );
  XOR3X1 U1896 ( .IN1(n2298), .IN2(n2297), .IN3(n2296), .Q(n2266) );
  OA22X1 U1897 ( .IN1(n2363), .IN2(\i_m4stg_frac/n807 ), .IN3(n2364), .IN4(
        \i_m4stg_frac/n961 ), .Q(n2296) );
  AND2X1 U1898 ( .IN1(\i_m4stg_frac/n807 ), .IN2(n2363), .Q(n2364) );
  AOI22X1 U1899 ( .IN1(\i_m4stg_frac/pc[49] ), .IN2(n1128), .IN3(
        \i_m4stg_frac/ps[50] ), .IN4(n2365), .QN(n2297) );
  OR2X1 U1900 ( .IN1(n1128), .IN2(\i_m4stg_frac/pc[49] ), .Q(n2365) );
  XOR3X1 U1901 ( .IN1(\i_m4stg_frac/n959 ), .IN2(\i_m4stg_frac/n805 ), .IN3(
        n2366), .Q(n2298) );
  AO22X1 U1902 ( .IN1(n2355), .IN2(n2356), .IN3(n2354), .IN4(n2367), .Q(n2265)
         );
  OR2X1 U1903 ( .IN1(n2356), .IN2(n2355), .Q(n2367) );
  XOR3X1 U1904 ( .IN1(\i_m4stg_frac/n961 ), .IN2(\i_m4stg_frac/n807 ), .IN3(
        n2363), .Q(n2354) );
  XNOR3X1 U1905 ( .IN1(\i_m4stg_frac/ps[50] ), .IN2(\i_m4stg_frac/pc[49] ), 
        .IN3(n1128), .Q(n2363) );
  OA22X1 U1906 ( .IN1(n2358), .IN2(\i_m4stg_frac/n809 ), .IN3(n2368), .IN4(
        \i_m4stg_frac/n963 ), .Q(n2356) );
  AND2X1 U1907 ( .IN1(\i_m4stg_frac/n809 ), .IN2(n2358), .Q(n2368) );
  XNOR3X1 U1908 ( .IN1(\i_m4stg_frac/ps[49] ), .IN2(\i_m4stg_frac/pc[48] ), 
        .IN3(n1129), .Q(n2358) );
  AOI22X1 U1909 ( .IN1(\i_m4stg_frac/pc[48] ), .IN2(n1129), .IN3(
        \i_m4stg_frac/ps[49] ), .IN4(n2369), .QN(n2355) );
  OR2X1 U1910 ( .IN1(n1129), .IN2(\i_m4stg_frac/pc[48] ), .Q(n2369) );
  NOR2X0 U1911 ( .IN1(se_mul64), .IN2(n2370), .QN(\i_m4stg_frac/n471 ) );
  XNOR2X1 U1912 ( .IN1(n2269), .IN2(n2270), .Q(n2370) );
  XOR3X1 U1913 ( .IN1(n2371), .IN2(n2372), .IN3(n2373), .Q(n2270) );
  AO22X1 U1914 ( .IN1(n2374), .IN2(n2375), .IN3(n2376), .IN4(n2377), .Q(n2269)
         );
  OR2X1 U1915 ( .IN1(n2374), .IN2(n2375), .Q(n2377) );
  NOR2X0 U1916 ( .IN1(se_mul64), .IN2(n2378), .QN(\i_m4stg_frac/n469 ) );
  XNOR2X1 U1917 ( .IN1(n2271), .IN2(n2272), .Q(n2378) );
  XOR3X1 U1918 ( .IN1(n2379), .IN2(n2380), .IN3(n2381), .Q(n2272) );
  AO22X1 U1919 ( .IN1(n2372), .IN2(n2373), .IN3(n2371), .IN4(n2382), .Q(n2271)
         );
  OR2X1 U1920 ( .IN1(n2373), .IN2(n2372), .Q(n2382) );
  XOR3X1 U1921 ( .IN1(\i_m4stg_frac/n953 ), .IN2(\i_m4stg_frac/n799 ), .IN3(
        \i_m4stg_frac/n486 ), .Q(n2371) );
  XNOR3X1 U1922 ( .IN1(n2383), .IN2(n2384), .IN3(n2385), .Q(n2373) );
  AOI22X1 U1923 ( .IN1(n2386), .IN2(n2387), .IN3(n2388), .IN4(n2389), .QN(
        n2372) );
  OR2X1 U1924 ( .IN1(n2387), .IN2(n2386), .Q(n2389) );
  NOR2X0 U1925 ( .IN1(se_mul64), .IN2(n2390), .QN(\i_m4stg_frac/n467 ) );
  XNOR2X1 U1926 ( .IN1(n2273), .IN2(n2274), .Q(n2390) );
  XOR3X1 U1927 ( .IN1(n2391), .IN2(n2392), .IN3(n2393), .Q(n2274) );
  AO22X1 U1928 ( .IN1(n2380), .IN2(n2381), .IN3(n2379), .IN4(n2394), .Q(n2273)
         );
  OR2X1 U1929 ( .IN1(n2381), .IN2(n2380), .Q(n2394) );
  XOR3X1 U1930 ( .IN1(\i_m4stg_frac/n951 ), .IN2(\i_m4stg_frac/n797 ), .IN3(
        \i_m4stg_frac/n484 ), .Q(n2379) );
  XNOR3X1 U1931 ( .IN1(n2395), .IN2(n2396), .IN3(n2397), .Q(n2381) );
  AOI22X1 U1932 ( .IN1(n2384), .IN2(n2383), .IN3(n2385), .IN4(n2398), .QN(
        n2380) );
  OR2X1 U1933 ( .IN1(n2384), .IN2(n2383), .Q(n2398) );
  XOR3X1 U1934 ( .IN1(\i_m4stg_frac/ps[54] ), .IN2(\i_m4stg_frac/pc[53] ), 
        .IN3(n1061), .Q(n2385) );
  AO22X1 U1935 ( .IN1(\i_m4stg_frac/pc[52] ), .IN2(n1191), .IN3(
        \i_m4stg_frac/ps[53] ), .IN4(n2399), .Q(n2383) );
  OR2X1 U1936 ( .IN1(n1191), .IN2(\i_m4stg_frac/pc[52] ), .Q(n2399) );
  OAI22X1 U1937 ( .IN1(\i_m4stg_frac/n488 ), .IN2(\i_m4stg_frac/n801 ), .IN3(
        n2400), .IN4(\i_m4stg_frac/n955 ), .QN(n2384) );
  AND2X1 U1938 ( .IN1(\i_m4stg_frac/n488 ), .IN2(\i_m4stg_frac/n801 ), .Q(
        n2400) );
  NOR2X0 U1939 ( .IN1(se_mul64), .IN2(n2401), .QN(\i_m4stg_frac/n465 ) );
  XNOR2X1 U1940 ( .IN1(n2275), .IN2(n2276), .Q(n2401) );
  XOR3X1 U1941 ( .IN1(n2402), .IN2(n2403), .IN3(n2404), .Q(n2276) );
  AO22X1 U1942 ( .IN1(n2392), .IN2(n2393), .IN3(n2391), .IN4(n2405), .Q(n2275)
         );
  OR2X1 U1943 ( .IN1(n2393), .IN2(n2392), .Q(n2405) );
  XOR3X1 U1944 ( .IN1(\i_m4stg_frac/n949 ), .IN2(\i_m4stg_frac/n795 ), .IN3(
        \i_m4stg_frac/n482 ), .Q(n2391) );
  XNOR3X1 U1945 ( .IN1(n2406), .IN2(n2407), .IN3(n2408), .Q(n2393) );
  AOI22X1 U1946 ( .IN1(n2396), .IN2(n2395), .IN3(n2397), .IN4(n2409), .QN(
        n2392) );
  OR2X1 U1947 ( .IN1(n2396), .IN2(n2395), .Q(n2409) );
  XOR3X1 U1948 ( .IN1(\i_m4stg_frac/ps[55] ), .IN2(\i_m4stg_frac/pc[54] ), 
        .IN3(n1062), .Q(n2397) );
  AO22X1 U1949 ( .IN1(\i_m4stg_frac/pc[53] ), .IN2(n1061), .IN3(
        \i_m4stg_frac/ps[54] ), .IN4(n2410), .Q(n2395) );
  OR2X1 U1950 ( .IN1(n1061), .IN2(\i_m4stg_frac/pc[53] ), .Q(n2410) );
  OAI22X1 U1951 ( .IN1(\i_m4stg_frac/n486 ), .IN2(\i_m4stg_frac/n799 ), .IN3(
        n2411), .IN4(\i_m4stg_frac/n953 ), .QN(n2396) );
  AND2X1 U1952 ( .IN1(\i_m4stg_frac/n486 ), .IN2(\i_m4stg_frac/n799 ), .Q(
        n2411) );
  NOR2X0 U1953 ( .IN1(se_mul64), .IN2(n2412), .QN(\i_m4stg_frac/n463 ) );
  XNOR2X1 U1954 ( .IN1(n2277), .IN2(n2278), .Q(n2412) );
  XOR3X1 U1955 ( .IN1(n2413), .IN2(n2414), .IN3(n2415), .Q(n2278) );
  AO22X1 U1956 ( .IN1(n2403), .IN2(n2404), .IN3(n2402), .IN4(n2416), .Q(n2277)
         );
  OR2X1 U1957 ( .IN1(n2404), .IN2(n2403), .Q(n2416) );
  XOR3X1 U1958 ( .IN1(\i_m4stg_frac/n947 ), .IN2(\i_m4stg_frac/n793 ), .IN3(
        \i_m4stg_frac/n480 ), .Q(n2402) );
  XNOR3X1 U1959 ( .IN1(n2417), .IN2(n2418), .IN3(n2419), .Q(n2404) );
  AOI22X1 U1960 ( .IN1(n2407), .IN2(n2406), .IN3(n2408), .IN4(n2420), .QN(
        n2403) );
  OR2X1 U1961 ( .IN1(n2407), .IN2(n2406), .Q(n2420) );
  XOR3X1 U1962 ( .IN1(\i_m4stg_frac/ps[56] ), .IN2(\i_m4stg_frac/pc[55] ), 
        .IN3(n1063), .Q(n2408) );
  AO22X1 U1963 ( .IN1(\i_m4stg_frac/pc[54] ), .IN2(n1062), .IN3(
        \i_m4stg_frac/ps[55] ), .IN4(n2421), .Q(n2406) );
  OR2X1 U1964 ( .IN1(n1062), .IN2(\i_m4stg_frac/pc[54] ), .Q(n2421) );
  OAI22X1 U1965 ( .IN1(\i_m4stg_frac/n484 ), .IN2(\i_m4stg_frac/n797 ), .IN3(
        n2422), .IN4(\i_m4stg_frac/n951 ), .QN(n2407) );
  AND2X1 U1966 ( .IN1(\i_m4stg_frac/n484 ), .IN2(\i_m4stg_frac/n797 ), .Q(
        n2422) );
  NOR2X0 U1967 ( .IN1(se_mul64), .IN2(n2423), .QN(\i_m4stg_frac/n461 ) );
  XNOR2X1 U1968 ( .IN1(n2279), .IN2(n2280), .Q(n2423) );
  XOR3X1 U1969 ( .IN1(n2424), .IN2(n2425), .IN3(n2426), .Q(n2280) );
  AO22X1 U1970 ( .IN1(n2414), .IN2(n2415), .IN3(n2413), .IN4(n2427), .Q(n2279)
         );
  OR2X1 U1971 ( .IN1(n2415), .IN2(n2414), .Q(n2427) );
  XOR3X1 U1972 ( .IN1(\i_m4stg_frac/n945 ), .IN2(\i_m4stg_frac/n791 ), .IN3(
        \i_m4stg_frac/n478 ), .Q(n2413) );
  XNOR3X1 U1973 ( .IN1(n2428), .IN2(n2429), .IN3(n2430), .Q(n2415) );
  AOI22X1 U1974 ( .IN1(n2418), .IN2(n2417), .IN3(n2419), .IN4(n2431), .QN(
        n2414) );
  OR2X1 U1975 ( .IN1(n2418), .IN2(n2417), .Q(n2431) );
  XOR3X1 U1976 ( .IN1(\i_m4stg_frac/ps[57] ), .IN2(\i_m4stg_frac/pc[56] ), 
        .IN3(n1064), .Q(n2419) );
  AO22X1 U1977 ( .IN1(\i_m4stg_frac/pc[55] ), .IN2(n1063), .IN3(
        \i_m4stg_frac/ps[56] ), .IN4(n2432), .Q(n2417) );
  OR2X1 U1978 ( .IN1(n1063), .IN2(\i_m4stg_frac/pc[55] ), .Q(n2432) );
  OAI22X1 U1979 ( .IN1(\i_m4stg_frac/n482 ), .IN2(\i_m4stg_frac/n795 ), .IN3(
        n2433), .IN4(\i_m4stg_frac/n949 ), .QN(n2418) );
  AND2X1 U1980 ( .IN1(\i_m4stg_frac/n482 ), .IN2(\i_m4stg_frac/n795 ), .Q(
        n2433) );
  NOR2X0 U1981 ( .IN1(se_mul64), .IN2(n2434), .QN(\i_m4stg_frac/n459 ) );
  XNOR2X1 U1982 ( .IN1(n2281), .IN2(n2282), .Q(n2434) );
  XOR3X1 U1983 ( .IN1(n2435), .IN2(n2436), .IN3(n2437), .Q(n2282) );
  AO22X1 U1984 ( .IN1(n2425), .IN2(n2426), .IN3(n2424), .IN4(n2438), .Q(n2281)
         );
  OR2X1 U1985 ( .IN1(n2426), .IN2(n2425), .Q(n2438) );
  XOR3X1 U1986 ( .IN1(\i_m4stg_frac/n943 ), .IN2(\i_m4stg_frac/n789 ), .IN3(
        \i_m4stg_frac/n476 ), .Q(n2424) );
  XNOR3X1 U1987 ( .IN1(n2439), .IN2(n2440), .IN3(n2441), .Q(n2426) );
  AOI22X1 U1988 ( .IN1(n2429), .IN2(n2428), .IN3(n2430), .IN4(n2442), .QN(
        n2425) );
  OR2X1 U1989 ( .IN1(n2429), .IN2(n2428), .Q(n2442) );
  XOR3X1 U1990 ( .IN1(\i_m4stg_frac/ps[58] ), .IN2(\i_m4stg_frac/pc[57] ), 
        .IN3(n1065), .Q(n2430) );
  AO22X1 U1991 ( .IN1(\i_m4stg_frac/pc[56] ), .IN2(n1064), .IN3(
        \i_m4stg_frac/ps[57] ), .IN4(n2443), .Q(n2428) );
  OR2X1 U1992 ( .IN1(n1064), .IN2(\i_m4stg_frac/pc[56] ), .Q(n2443) );
  OAI22X1 U1993 ( .IN1(\i_m4stg_frac/n480 ), .IN2(\i_m4stg_frac/n793 ), .IN3(
        n2444), .IN4(\i_m4stg_frac/n947 ), .QN(n2429) );
  AND2X1 U1994 ( .IN1(\i_m4stg_frac/n480 ), .IN2(\i_m4stg_frac/n793 ), .Q(
        n2444) );
  NOR2X0 U1995 ( .IN1(se_mul64), .IN2(n2445), .QN(\i_m4stg_frac/n457 ) );
  XNOR2X1 U1996 ( .IN1(n2283), .IN2(n2284), .Q(n2445) );
  XOR3X1 U1997 ( .IN1(n2446), .IN2(n2447), .IN3(n2448), .Q(n2284) );
  AO22X1 U1998 ( .IN1(n2436), .IN2(n2437), .IN3(n2435), .IN4(n2449), .Q(n2283)
         );
  OR2X1 U1999 ( .IN1(n2437), .IN2(n2436), .Q(n2449) );
  XOR3X1 U2000 ( .IN1(\i_m4stg_frac/n941 ), .IN2(\i_m4stg_frac/n787 ), .IN3(
        \i_m4stg_frac/n474 ), .Q(n2435) );
  XNOR3X1 U2001 ( .IN1(n2450), .IN2(n2451), .IN3(n2452), .Q(n2437) );
  AOI22X1 U2002 ( .IN1(n2440), .IN2(n2439), .IN3(n2441), .IN4(n2453), .QN(
        n2436) );
  OR2X1 U2003 ( .IN1(n2440), .IN2(n2439), .Q(n2453) );
  XOR3X1 U2004 ( .IN1(\i_m4stg_frac/ps[59] ), .IN2(\i_m4stg_frac/pc[58] ), 
        .IN3(n1066), .Q(n2441) );
  AO22X1 U2005 ( .IN1(\i_m4stg_frac/pc[57] ), .IN2(n1065), .IN3(
        \i_m4stg_frac/ps[58] ), .IN4(n2454), .Q(n2439) );
  OR2X1 U2006 ( .IN1(n1065), .IN2(\i_m4stg_frac/pc[57] ), .Q(n2454) );
  OAI22X1 U2007 ( .IN1(\i_m4stg_frac/n478 ), .IN2(\i_m4stg_frac/n791 ), .IN3(
        n2455), .IN4(\i_m4stg_frac/n945 ), .QN(n2440) );
  AND2X1 U2008 ( .IN1(\i_m4stg_frac/n478 ), .IN2(\i_m4stg_frac/n791 ), .Q(
        n2455) );
  NOR2X0 U2009 ( .IN1(se_mul64), .IN2(n2456), .QN(\i_m4stg_frac/n455 ) );
  XNOR2X1 U2010 ( .IN1(n2285), .IN2(n2286), .Q(n2456) );
  XOR3X1 U2011 ( .IN1(n2457), .IN2(n2458), .IN3(n2459), .Q(n2286) );
  AO22X1 U2012 ( .IN1(n2447), .IN2(n2448), .IN3(n2446), .IN4(n2460), .Q(n2285)
         );
  OR2X1 U2013 ( .IN1(n2448), .IN2(n2447), .Q(n2460) );
  XOR3X1 U2014 ( .IN1(\i_m4stg_frac/n939 ), .IN2(\i_m4stg_frac/n785 ), .IN3(
        \i_m4stg_frac/n472 ), .Q(n2446) );
  XNOR3X1 U2015 ( .IN1(n2461), .IN2(n2462), .IN3(n2463), .Q(n2448) );
  AOI22X1 U2016 ( .IN1(n2451), .IN2(n2450), .IN3(n2452), .IN4(n2464), .QN(
        n2447) );
  OR2X1 U2017 ( .IN1(n2451), .IN2(n2450), .Q(n2464) );
  XOR3X1 U2018 ( .IN1(\i_m4stg_frac/ps[60] ), .IN2(\i_m4stg_frac/pc[59] ), 
        .IN3(n1067), .Q(n2452) );
  AO22X1 U2019 ( .IN1(\i_m4stg_frac/pc[58] ), .IN2(n1066), .IN3(
        \i_m4stg_frac/ps[59] ), .IN4(n2465), .Q(n2450) );
  OR2X1 U2020 ( .IN1(n1066), .IN2(\i_m4stg_frac/pc[58] ), .Q(n2465) );
  OAI22X1 U2021 ( .IN1(\i_m4stg_frac/n476 ), .IN2(\i_m4stg_frac/n789 ), .IN3(
        n2466), .IN4(\i_m4stg_frac/n943 ), .QN(n2451) );
  AND2X1 U2022 ( .IN1(\i_m4stg_frac/n476 ), .IN2(\i_m4stg_frac/n789 ), .Q(
        n2466) );
  NOR2X0 U2023 ( .IN1(se_mul64), .IN2(n2467), .QN(\i_m4stg_frac/n453 ) );
  XNOR2X1 U2024 ( .IN1(n2134), .IN2(n2133), .Q(n2467) );
  XOR3X1 U2025 ( .IN1(n2468), .IN2(n2469), .IN3(n2470), .Q(n2133) );
  AO22X1 U2026 ( .IN1(n2471), .IN2(n2472), .IN3(n2457), .IN4(n2473), .Q(n2134)
         );
  NAND2X0 U2027 ( .IN1(n2459), .IN2(n2458), .QN(n2473) );
  XOR3X1 U2028 ( .IN1(\i_m4stg_frac/n937 ), .IN2(\i_m4stg_frac/n783 ), .IN3(
        \i_m4stg_frac/n470 ), .Q(n2457) );
  INVX0 U2029 ( .INP(n2459), .ZN(n2472) );
  XOR3X1 U2030 ( .IN1(n2474), .IN2(n2475), .IN3(n2476), .Q(n2459) );
  INVX0 U2031 ( .INP(n2458), .ZN(n2471) );
  AO22X1 U2032 ( .IN1(n2462), .IN2(n2461), .IN3(n2463), .IN4(n2477), .Q(n2458)
         );
  OR2X1 U2033 ( .IN1(n2461), .IN2(n2462), .Q(n2477) );
  XOR3X1 U2034 ( .IN1(\i_m4stg_frac/ps[61] ), .IN2(\i_m4stg_frac/pc[60] ), 
        .IN3(n1074), .Q(n2463) );
  AO22X1 U2035 ( .IN1(\i_m4stg_frac/pc[59] ), .IN2(n1067), .IN3(
        \i_m4stg_frac/ps[60] ), .IN4(n2478), .Q(n2461) );
  OR2X1 U2036 ( .IN1(n1067), .IN2(\i_m4stg_frac/pc[59] ), .Q(n2478) );
  OAI22X1 U2037 ( .IN1(\i_m4stg_frac/n474 ), .IN2(\i_m4stg_frac/n787 ), .IN3(
        n2479), .IN4(\i_m4stg_frac/n941 ), .QN(n2462) );
  AND2X1 U2038 ( .IN1(\i_m4stg_frac/n787 ), .IN2(\i_m4stg_frac/n474 ), .Q(
        n2479) );
  NOR2X0 U2039 ( .IN1(se_mul64), .IN2(n2480), .QN(\i_m4stg_frac/n451 ) );
  XNOR2X1 U2040 ( .IN1(n2199), .IN2(n2200), .Q(n2480) );
  XNOR3X1 U2041 ( .IN1(\i_m4stg_frac/n825 ), .IN2(n2481), .IN3(n2482), .Q(
        n2200) );
  AO22X1 U2042 ( .IN1(n2483), .IN2(n2484), .IN3(\i_m4stg_frac/n827 ), .IN4(
        n2485), .Q(n2199) );
  NAND2X0 U2043 ( .IN1(n2315), .IN2(n2314), .QN(n2485) );
  INVX0 U2044 ( .INP(n2315), .ZN(n2484) );
  XOR3X1 U2045 ( .IN1(\i_m4stg_frac/ps[40] ), .IN2(\i_m4stg_frac/pc[39] ), 
        .IN3(n1071), .Q(n2315) );
  INVX0 U2046 ( .INP(n2314), .ZN(n2483) );
  AO22X1 U2047 ( .IN1(\i_m4stg_frac/pc[38] ), .IN2(n1068), .IN3(
        \i_m4stg_frac/ps[39] ), .IN4(n2486), .Q(n2314) );
  OR2X1 U2048 ( .IN1(n1068), .IN2(\i_m4stg_frac/pc[38] ), .Q(n2486) );
  NOR2X0 U2049 ( .IN1(se_mul64), .IN2(n2487), .QN(\i_m4stg_frac/n449 ) );
  XNOR2X1 U2050 ( .IN1(n2251), .IN2(n2252), .Q(n2487) );
  XNOR3X1 U2051 ( .IN1(\i_m4stg_frac/n823 ), .IN2(n2321), .IN3(n2324), .Q(
        n2252) );
  XOR3X1 U2052 ( .IN1(\i_m4stg_frac/ps[42] ), .IN2(\i_m4stg_frac/pc[41] ), 
        .IN3(n1069), .Q(n2324) );
  INVX0 U2053 ( .INP(n2325), .ZN(n2321) );
  AO22X1 U2054 ( .IN1(\i_m4stg_frac/pc[40] ), .IN2(n1070), .IN3(
        \i_m4stg_frac/ps[41] ), .IN4(n2488), .Q(n2325) );
  OR2X1 U2055 ( .IN1(n1070), .IN2(\i_m4stg_frac/pc[40] ), .Q(n2488) );
  AO22X1 U2056 ( .IN1(n2481), .IN2(n2489), .IN3(\i_m4stg_frac/n825 ), .IN4(
        n2490), .Q(n2251) );
  NAND2X0 U2057 ( .IN1(n2482), .IN2(n2491), .QN(n2490) );
  INVX0 U2058 ( .INP(n2482), .ZN(n2489) );
  XOR3X1 U2059 ( .IN1(\i_m4stg_frac/ps[41] ), .IN2(\i_m4stg_frac/pc[40] ), 
        .IN3(n1070), .Q(n2482) );
  INVX0 U2060 ( .INP(n2491), .ZN(n2481) );
  AO22X1 U2061 ( .IN1(\i_m4stg_frac/pc[39] ), .IN2(n1071), .IN3(
        \i_m4stg_frac/ps[40] ), .IN4(n2492), .Q(n2491) );
  OR2X1 U2062 ( .IN1(n1071), .IN2(\i_m4stg_frac/pc[39] ), .Q(n2492) );
  NOR2X0 U2063 ( .IN1(se_mul64), .IN2(n2493), .QN(\i_m4stg_frac/n447 ) );
  XNOR2X1 U2064 ( .IN1(n2259), .IN2(n2260), .Q(n2493) );
  XOR3X1 U2065 ( .IN1(\i_m4stg_frac/n815 ), .IN2(n2494), .IN3(n2495), .Q(n2260) );
  AO22X1 U2066 ( .IN1(n2334), .IN2(n2496), .IN3(\i_m4stg_frac/n817 ), .IN4(
        n2497), .Q(n2259) );
  NAND2X0 U2067 ( .IN1(n2335), .IN2(n2498), .QN(n2497) );
  INVX0 U2068 ( .INP(n2335), .ZN(n2496) );
  XOR3X1 U2069 ( .IN1(\i_m4stg_frac/ps[45] ), .IN2(\i_m4stg_frac/pc[44] ), 
        .IN3(n1112), .Q(n2335) );
  INVX0 U2070 ( .INP(n2498), .ZN(n2334) );
  AO22X1 U2071 ( .IN1(\i_m4stg_frac/pc[43] ), .IN2(n1072), .IN3(
        \i_m4stg_frac/ps[44] ), .IN4(n2499), .Q(n2498) );
  OR2X1 U2072 ( .IN1(n1072), .IN2(\i_m4stg_frac/pc[43] ), .Q(n2499) );
  NOR3X0 U2073 ( .IN1(n2500), .IN2(se_mul64), .IN3(n2209), .QN(
        \i_m4stg_frac/n445 ) );
  XNOR3X1 U2074 ( .IN1(\i_m4stg_frac/n833 ), .IN2(n2303), .IN3(n2306), .Q(
        n2209) );
  XOR3X1 U2075 ( .IN1(\i_m4stg_frac/ps[37] ), .IN2(\i_m4stg_frac/pc[36] ), 
        .IN3(n1073), .Q(n2306) );
  INVX0 U2076 ( .INP(n2307), .ZN(n2303) );
  AO22X1 U2077 ( .IN1(\i_m4stg_frac/pc[35] ), .IN2(n1184), .IN3(
        \i_m4stg_frac/ps[36] ), .IN4(n2501), .Q(n2307) );
  OR2X1 U2078 ( .IN1(n1184), .IN2(\i_m4stg_frac/pc[35] ), .Q(n2501) );
  AND3X1 U2079 ( .IN1(n2250), .IN2(\i_m4stg_frac/n854 ), .IN3(n2249), .Q(
        \i_m4stg_frac/n443 ) );
  XNOR3X1 U2080 ( .IN1(n2376), .IN2(n2374), .IN3(n2375), .Q(n2249) );
  OA22X1 U2081 ( .IN1(n2502), .IN2(n2503), .IN3(n2504), .IN4(n2505), .Q(n2375)
         );
  AND2X1 U2082 ( .IN1(n2502), .IN2(n2503), .Q(n2505) );
  XNOR3X1 U2083 ( .IN1(n2388), .IN2(n2387), .IN3(n2386), .Q(n2374) );
  XNOR3X1 U2084 ( .IN1(\i_m4stg_frac/ps[53] ), .IN2(\i_m4stg_frac/pc[52] ), 
        .IN3(\i_m4stg_frac/n642 ), .Q(n2386) );
  AO22X1 U2085 ( .IN1(\i_m4stg_frac/pc[51] ), .IN2(n1126), .IN3(
        \i_m4stg_frac/ps[52] ), .IN4(n2506), .Q(n2387) );
  OR2X1 U2086 ( .IN1(n1126), .IN2(\i_m4stg_frac/pc[51] ), .Q(n2506) );
  XOR3X1 U2087 ( .IN1(\i_m4stg_frac/n955 ), .IN2(\i_m4stg_frac/n801 ), .IN3(
        \i_m4stg_frac/n488 ), .Q(n2376) );
  NOR2X0 U2088 ( .IN1(n2295), .IN2(n2294), .QN(n2250) );
  XOR3X1 U2089 ( .IN1(n2504), .IN2(n2502), .IN3(n2503), .Q(n2294) );
  OA22X1 U2090 ( .IN1(n2366), .IN2(\i_m4stg_frac/n805 ), .IN3(n2507), .IN4(
        \i_m4stg_frac/n959 ), .Q(n2503) );
  AND2X1 U2091 ( .IN1(\i_m4stg_frac/n805 ), .IN2(n2366), .Q(n2507) );
  XNOR3X1 U2092 ( .IN1(\i_m4stg_frac/ps[51] ), .IN2(\i_m4stg_frac/pc[50] ), 
        .IN3(n1130), .Q(n2366) );
  AOI22X1 U2093 ( .IN1(\i_m4stg_frac/pc[50] ), .IN2(n1130), .IN3(
        \i_m4stg_frac/ps[51] ), .IN4(n2508), .QN(n2502) );
  OR2X1 U2094 ( .IN1(n1130), .IN2(\i_m4stg_frac/pc[50] ), .Q(n2508) );
  XNOR3X1 U2095 ( .IN1(\i_m4stg_frac/ps[52] ), .IN2(\i_m4stg_frac/pc[51] ), 
        .IN3(n1126), .Q(n2504) );
  AO21X1 U2096 ( .IN1(\i_m4stg_frac/n957 ), .IN2(\i_m4stg_frac/n803 ), .IN3(
        n2388), .Q(n2295) );
  NOR2X0 U2097 ( .IN1(\i_m4stg_frac/n957 ), .IN2(\i_m4stg_frac/n803 ), .QN(
        n2388) );
  NOR2X0 U2098 ( .IN1(se_mul64), .IN2(n2024), .QN(\i_m4stg_frac/n441 ) );
  NAND2X0 U2099 ( .IN1(n2509), .IN2(n2128), .QN(n2024) );
  NAND3X0 U2100 ( .IN1(n2510), .IN2(n2127), .IN3(n2511), .QN(n2128) );
  AO21X1 U2101 ( .IN1(n2510), .IN2(n2127), .IN3(n2511), .Q(n2509) );
  AO22X1 U2102 ( .IN1(n2512), .IN2(n2513), .IN3(n2514), .IN4(n2515), .Q(n2511)
         );
  OR2X1 U2103 ( .IN1(n2513), .IN2(n2512), .Q(n2515) );
  OAI221X1 U2104 ( .IN1(n2516), .IN2(\i_m4stg_frac/n707 ), .IN3(n2517), .IN4(
        n2518), .IN5(n2519), .QN(n2510) );
  NOR2X0 U2105 ( .IN1(n2520), .IN2(n2521), .QN(n2516) );
  NOR2X0 U2106 ( .IN1(se_mul64), .IN2(n2026), .QN(\i_m4stg_frac/n439 ) );
  XNOR2X1 U2107 ( .IN1(n2106), .IN2(n2105), .Q(n2026) );
  XOR3X1 U2108 ( .IN1(n2522), .IN2(n2523), .IN3(n2524), .Q(n2105) );
  AO22X1 U2109 ( .IN1(n2469), .IN2(n2470), .IN3(n2468), .IN4(n2525), .Q(n2106)
         );
  OR2X1 U2110 ( .IN1(n2470), .IN2(n2469), .Q(n2525) );
  XOR3X1 U2111 ( .IN1(\i_m4stg_frac/n935 ), .IN2(\i_m4stg_frac/n781 ), .IN3(
        \i_m4stg_frac/n468 ), .Q(n2468) );
  XNOR3X1 U2112 ( .IN1(n2526), .IN2(n2527), .IN3(n2528), .Q(n2470) );
  AOI22X1 U2113 ( .IN1(n2475), .IN2(n2474), .IN3(n2476), .IN4(n2529), .QN(
        n2469) );
  OR2X1 U2114 ( .IN1(n2474), .IN2(n2475), .Q(n2529) );
  XOR3X1 U2115 ( .IN1(\i_m4stg_frac/ps[62] ), .IN2(\i_m4stg_frac/pc[61] ), 
        .IN3(n1075), .Q(n2476) );
  AO22X1 U2116 ( .IN1(\i_m4stg_frac/pc[60] ), .IN2(n1074), .IN3(
        \i_m4stg_frac/ps[61] ), .IN4(n2530), .Q(n2474) );
  OR2X1 U2117 ( .IN1(n1074), .IN2(\i_m4stg_frac/pc[60] ), .Q(n2530) );
  OAI22X1 U2118 ( .IN1(\i_m4stg_frac/n472 ), .IN2(\i_m4stg_frac/n785 ), .IN3(
        n2531), .IN4(\i_m4stg_frac/n939 ), .QN(n2475) );
  AND2X1 U2119 ( .IN1(\i_m4stg_frac/n785 ), .IN2(\i_m4stg_frac/n472 ), .Q(
        n2531) );
  NOR2X0 U2120 ( .IN1(se_mul64), .IN2(n1991), .QN(\i_m4stg_frac/n437 ) );
  XNOR2X1 U2121 ( .IN1(n2073), .IN2(n2072), .Q(n1991) );
  XOR3X1 U2122 ( .IN1(n2532), .IN2(n2533), .IN3(n2534), .Q(n2072) );
  AO22X1 U2123 ( .IN1(n2523), .IN2(n2524), .IN3(n2522), .IN4(n2535), .Q(n2073)
         );
  OR2X1 U2124 ( .IN1(n2524), .IN2(n2523), .Q(n2535) );
  XOR3X1 U2125 ( .IN1(\i_m4stg_frac/n933 ), .IN2(\i_m4stg_frac/n779 ), .IN3(
        \i_m4stg_frac/n466 ), .Q(n2522) );
  XNOR3X1 U2126 ( .IN1(n2536), .IN2(n2537), .IN3(n2538), .Q(n2524) );
  AOI22X1 U2127 ( .IN1(n2527), .IN2(n2526), .IN3(n2528), .IN4(n2539), .QN(
        n2523) );
  OR2X1 U2128 ( .IN1(n2526), .IN2(n2527), .Q(n2539) );
  XOR3X1 U2129 ( .IN1(\i_m4stg_frac/ps[63] ), .IN2(\i_m4stg_frac/pc[62] ), 
        .IN3(n1076), .Q(n2528) );
  AO22X1 U2130 ( .IN1(\i_m4stg_frac/pc[61] ), .IN2(n1075), .IN3(
        \i_m4stg_frac/ps[62] ), .IN4(n2540), .Q(n2526) );
  OR2X1 U2131 ( .IN1(n1075), .IN2(\i_m4stg_frac/pc[61] ), .Q(n2540) );
  OAI22X1 U2132 ( .IN1(\i_m4stg_frac/n470 ), .IN2(\i_m4stg_frac/n783 ), .IN3(
        n2541), .IN4(\i_m4stg_frac/n937 ), .QN(n2527) );
  AND2X1 U2133 ( .IN1(\i_m4stg_frac/n783 ), .IN2(\i_m4stg_frac/n470 ), .Q(
        n2541) );
  NOR2X0 U2134 ( .IN1(se_mul64), .IN2(n1938), .QN(\i_m4stg_frac/n435 ) );
  XNOR2X1 U2135 ( .IN1(n2062), .IN2(n2061), .Q(n1938) );
  XOR3X1 U2136 ( .IN1(n2542), .IN2(n2543), .IN3(n2544), .Q(n2061) );
  AO22X1 U2137 ( .IN1(n2533), .IN2(n2534), .IN3(n2532), .IN4(n2545), .Q(n2062)
         );
  OR2X1 U2138 ( .IN1(n2534), .IN2(n2533), .Q(n2545) );
  XOR3X1 U2139 ( .IN1(\i_m4stg_frac/n931 ), .IN2(\i_m4stg_frac/n777 ), .IN3(
        \i_m4stg_frac/n464 ), .Q(n2532) );
  XNOR3X1 U2140 ( .IN1(n2546), .IN2(n2547), .IN3(n2548), .Q(n2534) );
  AOI22X1 U2141 ( .IN1(n2537), .IN2(n2536), .IN3(n2538), .IN4(n2549), .QN(
        n2533) );
  OR2X1 U2142 ( .IN1(n2536), .IN2(n2537), .Q(n2549) );
  XOR3X1 U2143 ( .IN1(\i_m4stg_frac/ps[64] ), .IN2(\i_m4stg_frac/pc[63] ), 
        .IN3(n1077), .Q(n2538) );
  AO22X1 U2144 ( .IN1(\i_m4stg_frac/pc[62] ), .IN2(n1076), .IN3(
        \i_m4stg_frac/ps[63] ), .IN4(n2550), .Q(n2536) );
  OR2X1 U2145 ( .IN1(n1076), .IN2(\i_m4stg_frac/pc[62] ), .Q(n2550) );
  OAI22X1 U2146 ( .IN1(\i_m4stg_frac/n468 ), .IN2(\i_m4stg_frac/n781 ), .IN3(
        n2551), .IN4(\i_m4stg_frac/n935 ), .QN(n2537) );
  AND2X1 U2147 ( .IN1(\i_m4stg_frac/n781 ), .IN2(\i_m4stg_frac/n468 ), .Q(
        n2551) );
  NOR2X0 U2148 ( .IN1(se_mul64), .IN2(n1890), .QN(\i_m4stg_frac/n433 ) );
  XNOR2X1 U2149 ( .IN1(n2060), .IN2(n2059), .Q(n1890) );
  XOR3X1 U2150 ( .IN1(n2552), .IN2(n2553), .IN3(n2554), .Q(n2059) );
  AO22X1 U2151 ( .IN1(n2543), .IN2(n2544), .IN3(n2542), .IN4(n2555), .Q(n2060)
         );
  OR2X1 U2152 ( .IN1(n2544), .IN2(n2543), .Q(n2555) );
  XOR3X1 U2153 ( .IN1(\i_m4stg_frac/n929 ), .IN2(\i_m4stg_frac/n775 ), .IN3(
        \i_m4stg_frac/n462 ), .Q(n2542) );
  XNOR3X1 U2154 ( .IN1(n2556), .IN2(n2557), .IN3(n2558), .Q(n2544) );
  AOI22X1 U2155 ( .IN1(n2547), .IN2(n2546), .IN3(n2548), .IN4(n2559), .QN(
        n2543) );
  OR2X1 U2156 ( .IN1(n2546), .IN2(n2547), .Q(n2559) );
  XOR3X1 U2157 ( .IN1(\i_m4stg_frac/ps[65] ), .IN2(\i_m4stg_frac/pc[64] ), 
        .IN3(n1078), .Q(n2548) );
  AO22X1 U2158 ( .IN1(\i_m4stg_frac/pc[63] ), .IN2(n1077), .IN3(
        \i_m4stg_frac/ps[64] ), .IN4(n2560), .Q(n2546) );
  OR2X1 U2159 ( .IN1(n1077), .IN2(\i_m4stg_frac/pc[63] ), .Q(n2560) );
  OAI22X1 U2160 ( .IN1(\i_m4stg_frac/n466 ), .IN2(\i_m4stg_frac/n779 ), .IN3(
        n2561), .IN4(\i_m4stg_frac/n933 ), .QN(n2547) );
  AND2X1 U2161 ( .IN1(\i_m4stg_frac/n779 ), .IN2(\i_m4stg_frac/n466 ), .Q(
        n2561) );
  NOR2X0 U2162 ( .IN1(se_mul64), .IN2(n1889), .QN(\i_m4stg_frac/n431 ) );
  XNOR2X1 U2163 ( .IN1(n2058), .IN2(n2057), .Q(n1889) );
  XOR3X1 U2164 ( .IN1(n2562), .IN2(n2563), .IN3(n2564), .Q(n2057) );
  AO22X1 U2165 ( .IN1(n2553), .IN2(n2554), .IN3(n2552), .IN4(n2565), .Q(n2058)
         );
  OR2X1 U2166 ( .IN1(n2554), .IN2(n2553), .Q(n2565) );
  XOR3X1 U2167 ( .IN1(\i_m4stg_frac/n927 ), .IN2(\i_m4stg_frac/n773 ), .IN3(
        \i_m4stg_frac/n460 ), .Q(n2552) );
  XNOR3X1 U2168 ( .IN1(n2566), .IN2(n2567), .IN3(n2568), .Q(n2554) );
  AOI22X1 U2169 ( .IN1(n2557), .IN2(n2556), .IN3(n2558), .IN4(n2569), .QN(
        n2553) );
  OR2X1 U2170 ( .IN1(n2556), .IN2(n2557), .Q(n2569) );
  XOR3X1 U2171 ( .IN1(\i_m4stg_frac/ps[66] ), .IN2(\i_m4stg_frac/pc[65] ), 
        .IN3(n1079), .Q(n2558) );
  AO22X1 U2172 ( .IN1(\i_m4stg_frac/pc[64] ), .IN2(n1078), .IN3(
        \i_m4stg_frac/ps[65] ), .IN4(n2570), .Q(n2556) );
  OR2X1 U2173 ( .IN1(n1078), .IN2(\i_m4stg_frac/pc[64] ), .Q(n2570) );
  OAI22X1 U2174 ( .IN1(\i_m4stg_frac/n464 ), .IN2(\i_m4stg_frac/n777 ), .IN3(
        n2571), .IN4(\i_m4stg_frac/n931 ), .QN(n2557) );
  AND2X1 U2175 ( .IN1(\i_m4stg_frac/n777 ), .IN2(\i_m4stg_frac/n464 ), .Q(
        n2571) );
  NOR2X0 U2176 ( .IN1(se_mul64), .IN2(n1888), .QN(\i_m4stg_frac/n429 ) );
  XOR2X1 U2177 ( .IN1(n2196), .IN2(n2195), .Q(n1888) );
  INVX0 U2178 ( .INP(n2287), .ZN(n2195) );
  AO22X1 U2179 ( .IN1(n2563), .IN2(n2564), .IN3(n2562), .IN4(n2572), .Q(n2287)
         );
  OR2X1 U2180 ( .IN1(n2564), .IN2(n2563), .Q(n2572) );
  XOR3X1 U2181 ( .IN1(\i_m4stg_frac/n925 ), .IN2(\i_m4stg_frac/n771 ), .IN3(
        \i_m4stg_frac/n458 ), .Q(n2562) );
  XNOR3X1 U2182 ( .IN1(n2573), .IN2(n2574), .IN3(n2575), .Q(n2564) );
  AOI22X1 U2183 ( .IN1(n2567), .IN2(n2566), .IN3(n2568), .IN4(n2576), .QN(
        n2563) );
  OR2X1 U2184 ( .IN1(n2566), .IN2(n2567), .Q(n2576) );
  XOR3X1 U2185 ( .IN1(\i_m4stg_frac/ps[67] ), .IN2(\i_m4stg_frac/pc[66] ), 
        .IN3(n1080), .Q(n2568) );
  AO22X1 U2186 ( .IN1(\i_m4stg_frac/pc[65] ), .IN2(n1079), .IN3(
        \i_m4stg_frac/ps[66] ), .IN4(n2577), .Q(n2566) );
  OR2X1 U2187 ( .IN1(n1079), .IN2(\i_m4stg_frac/pc[65] ), .Q(n2577) );
  OAI22X1 U2188 ( .IN1(\i_m4stg_frac/n462 ), .IN2(\i_m4stg_frac/n775 ), .IN3(
        n2578), .IN4(\i_m4stg_frac/n929 ), .QN(n2567) );
  AND2X1 U2189 ( .IN1(\i_m4stg_frac/n775 ), .IN2(\i_m4stg_frac/n462 ), .Q(
        n2578) );
  XOR3X1 U2190 ( .IN1(n2579), .IN2(n2580), .IN3(n2581), .Q(n2196) );
  NOR2X0 U2191 ( .IN1(se_mul64), .IN2(n2056), .QN(\i_m4stg_frac/n427 ) );
  XOR2X1 U2192 ( .IN1(n2193), .IN2(n2192), .Q(n2056) );
  INVX0 U2193 ( .INP(n2288), .ZN(n2192) );
  AO22X1 U2194 ( .IN1(n2580), .IN2(n2581), .IN3(n2579), .IN4(n2582), .Q(n2288)
         );
  OR2X1 U2195 ( .IN1(n2581), .IN2(n2580), .Q(n2582) );
  XOR3X1 U2196 ( .IN1(\i_m4stg_frac/n923 ), .IN2(\i_m4stg_frac/n769 ), .IN3(
        \i_m4stg_frac/n456 ), .Q(n2579) );
  XNOR3X1 U2197 ( .IN1(n2583), .IN2(n2584), .IN3(n2585), .Q(n2581) );
  AOI22X1 U2198 ( .IN1(n2574), .IN2(n2573), .IN3(n2575), .IN4(n2586), .QN(
        n2580) );
  OR2X1 U2199 ( .IN1(n2574), .IN2(n2573), .Q(n2586) );
  XOR3X1 U2200 ( .IN1(\i_m4stg_frac/ps[68] ), .IN2(\i_m4stg_frac/pc[67] ), 
        .IN3(n1081), .Q(n2575) );
  AO22X1 U2201 ( .IN1(\i_m4stg_frac/pc[66] ), .IN2(n1080), .IN3(
        \i_m4stg_frac/ps[67] ), .IN4(n2587), .Q(n2573) );
  OR2X1 U2202 ( .IN1(n1080), .IN2(\i_m4stg_frac/pc[66] ), .Q(n2587) );
  OAI22X1 U2203 ( .IN1(\i_m4stg_frac/n460 ), .IN2(\i_m4stg_frac/n773 ), .IN3(
        n2588), .IN4(\i_m4stg_frac/n927 ), .QN(n2574) );
  AND2X1 U2204 ( .IN1(\i_m4stg_frac/n773 ), .IN2(\i_m4stg_frac/n460 ), .Q(
        n2588) );
  XNOR3X1 U2205 ( .IN1(n2589), .IN2(n2590), .IN3(n2591), .Q(n2193) );
  NOR2X0 U2206 ( .IN1(se_mul64), .IN2(n2055), .QN(\i_m4stg_frac/n425 ) );
  XNOR2X1 U2207 ( .IN1(n2190), .IN2(n2189), .Q(n2055) );
  XOR3X1 U2208 ( .IN1(n2592), .IN2(n2593), .IN3(n2594), .Q(n2189) );
  AO22X1 U2209 ( .IN1(n2590), .IN2(n2595), .IN3(n2589), .IN4(n2596), .Q(n2190)
         );
  NAND2X0 U2210 ( .IN1(n2591), .IN2(n2597), .QN(n2596) );
  XOR3X1 U2211 ( .IN1(\i_m4stg_frac/n921 ), .IN2(\i_m4stg_frac/n767 ), .IN3(
        \i_m4stg_frac/n454 ), .Q(n2589) );
  INVX0 U2212 ( .INP(n2591), .ZN(n2595) );
  XOR3X1 U2213 ( .IN1(n2598), .IN2(n2599), .IN3(n2600), .Q(n2591) );
  INVX0 U2214 ( .INP(n2597), .ZN(n2590) );
  AO22X1 U2215 ( .IN1(n2584), .IN2(n2583), .IN3(n2585), .IN4(n2601), .Q(n2597)
         );
  OR2X1 U2216 ( .IN1(n2584), .IN2(n2583), .Q(n2601) );
  XOR3X1 U2217 ( .IN1(\i_m4stg_frac/ps[69] ), .IN2(\i_m4stg_frac/pc[68] ), 
        .IN3(n1082), .Q(n2585) );
  AO22X1 U2218 ( .IN1(\i_m4stg_frac/pc[67] ), .IN2(n1081), .IN3(
        \i_m4stg_frac/ps[68] ), .IN4(n2602), .Q(n2583) );
  OR2X1 U2219 ( .IN1(n1081), .IN2(\i_m4stg_frac/pc[67] ), .Q(n2602) );
  OAI22X1 U2220 ( .IN1(\i_m4stg_frac/n458 ), .IN2(\i_m4stg_frac/n771 ), .IN3(
        n2603), .IN4(\i_m4stg_frac/n925 ), .QN(n2584) );
  AND2X1 U2221 ( .IN1(\i_m4stg_frac/n458 ), .IN2(\i_m4stg_frac/n771 ), .Q(
        n2603) );
  NOR2X0 U2222 ( .IN1(se_mul64), .IN2(n2054), .QN(\i_m4stg_frac/n423 ) );
  XNOR2X1 U2223 ( .IN1(n2188), .IN2(n2187), .Q(n2054) );
  XOR3X1 U2224 ( .IN1(n2604), .IN2(n2605), .IN3(n2606), .Q(n2187) );
  AO22X1 U2225 ( .IN1(n2593), .IN2(n2594), .IN3(n2592), .IN4(n2607), .Q(n2188)
         );
  OR2X1 U2226 ( .IN1(n2594), .IN2(n2593), .Q(n2607) );
  XOR3X1 U2227 ( .IN1(\i_m4stg_frac/n919 ), .IN2(\i_m4stg_frac/n765 ), .IN3(
        \i_m4stg_frac/n452 ), .Q(n2592) );
  XNOR3X1 U2228 ( .IN1(n2608), .IN2(n2609), .IN3(n2610), .Q(n2594) );
  AOI22X1 U2229 ( .IN1(n2599), .IN2(n2598), .IN3(n2600), .IN4(n2611), .QN(
        n2593) );
  OR2X1 U2230 ( .IN1(n2598), .IN2(n2599), .Q(n2611) );
  XOR3X1 U2231 ( .IN1(\i_m4stg_frac/ps[70] ), .IN2(\i_m4stg_frac/pc[69] ), 
        .IN3(n1083), .Q(n2600) );
  AO22X1 U2232 ( .IN1(\i_m4stg_frac/pc[68] ), .IN2(n1082), .IN3(
        \i_m4stg_frac/ps[69] ), .IN4(n2612), .Q(n2598) );
  OR2X1 U2233 ( .IN1(n1082), .IN2(\i_m4stg_frac/pc[68] ), .Q(n2612) );
  OAI22X1 U2234 ( .IN1(\i_m4stg_frac/n456 ), .IN2(\i_m4stg_frac/n769 ), .IN3(
        n2613), .IN4(\i_m4stg_frac/n923 ), .QN(n2599) );
  AND2X1 U2235 ( .IN1(\i_m4stg_frac/n456 ), .IN2(\i_m4stg_frac/n769 ), .Q(
        n2613) );
  NOR2X0 U2236 ( .IN1(se_mul64), .IN2(n2053), .QN(\i_m4stg_frac/n421 ) );
  XNOR2X1 U2237 ( .IN1(n2186), .IN2(n2185), .Q(n2053) );
  XOR3X1 U2238 ( .IN1(n2614), .IN2(n2615), .IN3(n2616), .Q(n2185) );
  AO22X1 U2239 ( .IN1(n2605), .IN2(n2606), .IN3(n2604), .IN4(n2617), .Q(n2186)
         );
  OR2X1 U2240 ( .IN1(n2606), .IN2(n2605), .Q(n2617) );
  XOR3X1 U2241 ( .IN1(\i_m4stg_frac/n917 ), .IN2(\i_m4stg_frac/n763 ), .IN3(
        \i_m4stg_frac/n450 ), .Q(n2604) );
  XNOR3X1 U2242 ( .IN1(n2618), .IN2(n2619), .IN3(n2620), .Q(n2606) );
  AOI22X1 U2243 ( .IN1(n2609), .IN2(n2608), .IN3(n2610), .IN4(n2621), .QN(
        n2605) );
  OR2X1 U2244 ( .IN1(n2608), .IN2(n2609), .Q(n2621) );
  XOR3X1 U2245 ( .IN1(\i_m4stg_frac/ps[71] ), .IN2(\i_m4stg_frac/pc[70] ), 
        .IN3(n1084), .Q(n2610) );
  AO22X1 U2246 ( .IN1(\i_m4stg_frac/pc[69] ), .IN2(n1083), .IN3(
        \i_m4stg_frac/ps[70] ), .IN4(n2622), .Q(n2608) );
  OR2X1 U2247 ( .IN1(n1083), .IN2(\i_m4stg_frac/pc[69] ), .Q(n2622) );
  OAI22X1 U2248 ( .IN1(\i_m4stg_frac/n454 ), .IN2(\i_m4stg_frac/n767 ), .IN3(
        n2623), .IN4(\i_m4stg_frac/n921 ), .QN(n2609) );
  AND2X1 U2249 ( .IN1(\i_m4stg_frac/n767 ), .IN2(\i_m4stg_frac/n454 ), .Q(
        n2623) );
  NOR2X0 U2250 ( .IN1(se_mul64), .IN2(n2052), .QN(\i_m4stg_frac/n419 ) );
  XNOR2X1 U2251 ( .IN1(n2184), .IN2(n2183), .Q(n2052) );
  XOR3X1 U2252 ( .IN1(n2624), .IN2(n2625), .IN3(n2626), .Q(n2183) );
  AO22X1 U2253 ( .IN1(n2615), .IN2(n2616), .IN3(n2614), .IN4(n2627), .Q(n2184)
         );
  OR2X1 U2254 ( .IN1(n2616), .IN2(n2615), .Q(n2627) );
  XOR3X1 U2255 ( .IN1(\i_m4stg_frac/n915 ), .IN2(\i_m4stg_frac/n761 ), .IN3(
        \i_m4stg_frac/n448 ), .Q(n2614) );
  XNOR3X1 U2256 ( .IN1(n2628), .IN2(n2629), .IN3(n2630), .Q(n2616) );
  AOI22X1 U2257 ( .IN1(n2619), .IN2(n2618), .IN3(n2620), .IN4(n2631), .QN(
        n2615) );
  OR2X1 U2258 ( .IN1(n2618), .IN2(n2619), .Q(n2631) );
  XOR3X1 U2259 ( .IN1(\i_m4stg_frac/ps[72] ), .IN2(\i_m4stg_frac/pc[71] ), 
        .IN3(n1085), .Q(n2620) );
  AO22X1 U2260 ( .IN1(\i_m4stg_frac/pc[70] ), .IN2(n1084), .IN3(
        \i_m4stg_frac/ps[71] ), .IN4(n2632), .Q(n2618) );
  OR2X1 U2261 ( .IN1(n1084), .IN2(\i_m4stg_frac/pc[70] ), .Q(n2632) );
  OAI22X1 U2262 ( .IN1(\i_m4stg_frac/n452 ), .IN2(\i_m4stg_frac/n765 ), .IN3(
        n2633), .IN4(\i_m4stg_frac/n919 ), .QN(n2619) );
  AND2X1 U2263 ( .IN1(\i_m4stg_frac/n765 ), .IN2(\i_m4stg_frac/n452 ), .Q(
        n2633) );
  NOR2X0 U2264 ( .IN1(se_mul64), .IN2(n2051), .QN(\i_m4stg_frac/n417 ) );
  XNOR2X1 U2265 ( .IN1(n2182), .IN2(n2181), .Q(n2051) );
  XOR3X1 U2266 ( .IN1(n2634), .IN2(n2635), .IN3(n2636), .Q(n2181) );
  AO22X1 U2267 ( .IN1(n2625), .IN2(n2626), .IN3(n2624), .IN4(n2637), .Q(n2182)
         );
  OR2X1 U2268 ( .IN1(n2626), .IN2(n2625), .Q(n2637) );
  XOR3X1 U2269 ( .IN1(\i_m4stg_frac/n913 ), .IN2(\i_m4stg_frac/n759 ), .IN3(
        \i_m4stg_frac/n446 ), .Q(n2624) );
  XNOR3X1 U2270 ( .IN1(n2638), .IN2(n2639), .IN3(n2640), .Q(n2626) );
  AOI22X1 U2271 ( .IN1(n2629), .IN2(n2628), .IN3(n2630), .IN4(n2641), .QN(
        n2625) );
  OR2X1 U2272 ( .IN1(n2628), .IN2(n2629), .Q(n2641) );
  XOR3X1 U2273 ( .IN1(\i_m4stg_frac/ps[73] ), .IN2(\i_m4stg_frac/pc[72] ), 
        .IN3(n1086), .Q(n2630) );
  AO22X1 U2274 ( .IN1(\i_m4stg_frac/pc[71] ), .IN2(n1085), .IN3(
        \i_m4stg_frac/ps[72] ), .IN4(n2642), .Q(n2628) );
  OR2X1 U2275 ( .IN1(n1085), .IN2(\i_m4stg_frac/pc[71] ), .Q(n2642) );
  OAI22X1 U2276 ( .IN1(\i_m4stg_frac/n450 ), .IN2(\i_m4stg_frac/n763 ), .IN3(
        n2643), .IN4(\i_m4stg_frac/n917 ), .QN(n2629) );
  AND2X1 U2277 ( .IN1(\i_m4stg_frac/n763 ), .IN2(\i_m4stg_frac/n450 ), .Q(
        n2643) );
  NOR2X0 U2278 ( .IN1(se_mul64), .IN2(n2050), .QN(\i_m4stg_frac/n415 ) );
  XNOR2X1 U2279 ( .IN1(n2180), .IN2(n2179), .Q(n2050) );
  XOR3X1 U2280 ( .IN1(n2644), .IN2(n2645), .IN3(n2646), .Q(n2179) );
  AO22X1 U2281 ( .IN1(n2635), .IN2(n2636), .IN3(n2634), .IN4(n2647), .Q(n2180)
         );
  OR2X1 U2282 ( .IN1(n2636), .IN2(n2635), .Q(n2647) );
  XOR3X1 U2283 ( .IN1(\i_m4stg_frac/n911 ), .IN2(\i_m4stg_frac/n757 ), .IN3(
        \i_m4stg_frac/n444 ), .Q(n2634) );
  XNOR3X1 U2284 ( .IN1(n2648), .IN2(n2649), .IN3(n2650), .Q(n2636) );
  AOI22X1 U2285 ( .IN1(n2639), .IN2(n2638), .IN3(n2640), .IN4(n2651), .QN(
        n2635) );
  OR2X1 U2286 ( .IN1(n2638), .IN2(n2639), .Q(n2651) );
  XOR3X1 U2287 ( .IN1(\i_m4stg_frac/ps[74] ), .IN2(\i_m4stg_frac/pc[73] ), 
        .IN3(n1087), .Q(n2640) );
  AO22X1 U2288 ( .IN1(\i_m4stg_frac/pc[72] ), .IN2(n1086), .IN3(
        \i_m4stg_frac/ps[73] ), .IN4(n2652), .Q(n2638) );
  OR2X1 U2289 ( .IN1(n1086), .IN2(\i_m4stg_frac/pc[72] ), .Q(n2652) );
  OAI22X1 U2290 ( .IN1(\i_m4stg_frac/n448 ), .IN2(\i_m4stg_frac/n761 ), .IN3(
        n2653), .IN4(\i_m4stg_frac/n915 ), .QN(n2639) );
  AND2X1 U2291 ( .IN1(\i_m4stg_frac/n761 ), .IN2(\i_m4stg_frac/n448 ), .Q(
        n2653) );
  NOR2X0 U2292 ( .IN1(se_mul64), .IN2(n2049), .QN(\i_m4stg_frac/n413 ) );
  XNOR2X1 U2293 ( .IN1(n2178), .IN2(n2177), .Q(n2049) );
  XOR3X1 U2294 ( .IN1(n2654), .IN2(n2655), .IN3(n2656), .Q(n2177) );
  AO22X1 U2295 ( .IN1(n2645), .IN2(n2646), .IN3(n2644), .IN4(n2657), .Q(n2178)
         );
  OR2X1 U2296 ( .IN1(n2646), .IN2(n2645), .Q(n2657) );
  XOR3X1 U2297 ( .IN1(\i_m4stg_frac/n909 ), .IN2(\i_m4stg_frac/n755 ), .IN3(
        \i_m4stg_frac/n442 ), .Q(n2644) );
  XNOR3X1 U2298 ( .IN1(n2658), .IN2(n2659), .IN3(n2660), .Q(n2646) );
  AOI22X1 U2299 ( .IN1(n2649), .IN2(n2648), .IN3(n2650), .IN4(n2661), .QN(
        n2645) );
  OR2X1 U2300 ( .IN1(n2648), .IN2(n2649), .Q(n2661) );
  XOR3X1 U2301 ( .IN1(\i_m4stg_frac/ps[75] ), .IN2(\i_m4stg_frac/pc[74] ), 
        .IN3(n1088), .Q(n2650) );
  AO22X1 U2302 ( .IN1(\i_m4stg_frac/pc[73] ), .IN2(n1087), .IN3(
        \i_m4stg_frac/ps[74] ), .IN4(n2662), .Q(n2648) );
  OR2X1 U2303 ( .IN1(n1087), .IN2(\i_m4stg_frac/pc[73] ), .Q(n2662) );
  OAI22X1 U2304 ( .IN1(\i_m4stg_frac/n446 ), .IN2(\i_m4stg_frac/n759 ), .IN3(
        n2663), .IN4(\i_m4stg_frac/n913 ), .QN(n2649) );
  AND2X1 U2305 ( .IN1(\i_m4stg_frac/n759 ), .IN2(\i_m4stg_frac/n446 ), .Q(
        n2663) );
  NOR2X0 U2306 ( .IN1(se_mul64), .IN2(n2048), .QN(\i_m4stg_frac/n411 ) );
  XNOR2X1 U2307 ( .IN1(n2176), .IN2(n2175), .Q(n2048) );
  XOR3X1 U2308 ( .IN1(n2664), .IN2(n2665), .IN3(n2666), .Q(n2175) );
  AO22X1 U2309 ( .IN1(n2655), .IN2(n2656), .IN3(n2654), .IN4(n2667), .Q(n2176)
         );
  OR2X1 U2310 ( .IN1(n2656), .IN2(n2655), .Q(n2667) );
  XOR3X1 U2311 ( .IN1(\i_m4stg_frac/n907 ), .IN2(\i_m4stg_frac/n753 ), .IN3(
        \i_m4stg_frac/n440 ), .Q(n2654) );
  XNOR3X1 U2312 ( .IN1(n2668), .IN2(n2669), .IN3(n2670), .Q(n2656) );
  AOI22X1 U2313 ( .IN1(n2659), .IN2(n2658), .IN3(n2660), .IN4(n2671), .QN(
        n2655) );
  OR2X1 U2314 ( .IN1(n2658), .IN2(n2659), .Q(n2671) );
  XOR3X1 U2315 ( .IN1(\i_m4stg_frac/ps[76] ), .IN2(\i_m4stg_frac/pc[75] ), 
        .IN3(n1089), .Q(n2660) );
  AO22X1 U2316 ( .IN1(\i_m4stg_frac/pc[74] ), .IN2(n1088), .IN3(
        \i_m4stg_frac/ps[75] ), .IN4(n2672), .Q(n2658) );
  OR2X1 U2317 ( .IN1(n1088), .IN2(\i_m4stg_frac/pc[74] ), .Q(n2672) );
  OAI22X1 U2318 ( .IN1(\i_m4stg_frac/n444 ), .IN2(\i_m4stg_frac/n757 ), .IN3(
        n2673), .IN4(\i_m4stg_frac/n911 ), .QN(n2659) );
  AND2X1 U2319 ( .IN1(\i_m4stg_frac/n757 ), .IN2(\i_m4stg_frac/n444 ), .Q(
        n2673) );
  NOR2X0 U2320 ( .IN1(se_mul64), .IN2(n2047), .QN(\i_m4stg_frac/n409 ) );
  XNOR2X1 U2321 ( .IN1(n2174), .IN2(n2173), .Q(n2047) );
  XOR3X1 U2322 ( .IN1(n2674), .IN2(n2675), .IN3(n2676), .Q(n2173) );
  AO22X1 U2323 ( .IN1(n2665), .IN2(n2666), .IN3(n2664), .IN4(n2677), .Q(n2174)
         );
  OR2X1 U2324 ( .IN1(n2666), .IN2(n2665), .Q(n2677) );
  XOR3X1 U2325 ( .IN1(\i_m4stg_frac/n905 ), .IN2(\i_m4stg_frac/n751 ), .IN3(
        \i_m4stg_frac/n438 ), .Q(n2664) );
  XNOR3X1 U2326 ( .IN1(n2678), .IN2(n2679), .IN3(n2680), .Q(n2666) );
  AOI22X1 U2327 ( .IN1(n2669), .IN2(n2668), .IN3(n2670), .IN4(n2681), .QN(
        n2665) );
  OR2X1 U2328 ( .IN1(n2668), .IN2(n2669), .Q(n2681) );
  XOR3X1 U2329 ( .IN1(\i_m4stg_frac/ps[77] ), .IN2(\i_m4stg_frac/pc[76] ), 
        .IN3(n1090), .Q(n2670) );
  AO22X1 U2330 ( .IN1(\i_m4stg_frac/pc[75] ), .IN2(n1089), .IN3(
        \i_m4stg_frac/ps[76] ), .IN4(n2682), .Q(n2668) );
  OR2X1 U2331 ( .IN1(n1089), .IN2(\i_m4stg_frac/pc[75] ), .Q(n2682) );
  OAI22X1 U2332 ( .IN1(\i_m4stg_frac/n442 ), .IN2(\i_m4stg_frac/n755 ), .IN3(
        n2683), .IN4(\i_m4stg_frac/n909 ), .QN(n2669) );
  AND2X1 U2333 ( .IN1(\i_m4stg_frac/n755 ), .IN2(\i_m4stg_frac/n442 ), .Q(
        n2683) );
  NOR2X0 U2334 ( .IN1(se_mul64), .IN2(n2046), .QN(\i_m4stg_frac/n407 ) );
  XNOR2X1 U2335 ( .IN1(n2172), .IN2(n2171), .Q(n2046) );
  XOR3X1 U2336 ( .IN1(n2684), .IN2(n2685), .IN3(n2686), .Q(n2171) );
  AO22X1 U2337 ( .IN1(n2675), .IN2(n2676), .IN3(n2674), .IN4(n2687), .Q(n2172)
         );
  OR2X1 U2338 ( .IN1(n2676), .IN2(n2675), .Q(n2687) );
  XOR3X1 U2339 ( .IN1(\i_m4stg_frac/n903 ), .IN2(\i_m4stg_frac/n749 ), .IN3(
        \i_m4stg_frac/n436 ), .Q(n2674) );
  XNOR3X1 U2340 ( .IN1(n2688), .IN2(n2689), .IN3(n2690), .Q(n2676) );
  AOI22X1 U2341 ( .IN1(n2679), .IN2(n2678), .IN3(n2680), .IN4(n2691), .QN(
        n2675) );
  OR2X1 U2342 ( .IN1(n2678), .IN2(n2679), .Q(n2691) );
  XOR3X1 U2343 ( .IN1(\i_m4stg_frac/ps[78] ), .IN2(\i_m4stg_frac/pc[77] ), 
        .IN3(n1091), .Q(n2680) );
  AO22X1 U2344 ( .IN1(\i_m4stg_frac/pc[76] ), .IN2(n1090), .IN3(
        \i_m4stg_frac/ps[77] ), .IN4(n2692), .Q(n2678) );
  OR2X1 U2345 ( .IN1(n1090), .IN2(\i_m4stg_frac/pc[76] ), .Q(n2692) );
  OAI22X1 U2346 ( .IN1(\i_m4stg_frac/n440 ), .IN2(\i_m4stg_frac/n753 ), .IN3(
        n2693), .IN4(\i_m4stg_frac/n907 ), .QN(n2679) );
  AND2X1 U2347 ( .IN1(\i_m4stg_frac/n753 ), .IN2(\i_m4stg_frac/n440 ), .Q(
        n2693) );
  NOR2X0 U2348 ( .IN1(se_mul64), .IN2(n2045), .QN(\i_m4stg_frac/n405 ) );
  XNOR2X1 U2349 ( .IN1(n2170), .IN2(n2169), .Q(n2045) );
  XOR3X1 U2350 ( .IN1(n2694), .IN2(n2695), .IN3(n2696), .Q(n2169) );
  AO22X1 U2351 ( .IN1(n2685), .IN2(n2686), .IN3(n2684), .IN4(n2697), .Q(n2170)
         );
  OR2X1 U2352 ( .IN1(n2686), .IN2(n2685), .Q(n2697) );
  XOR3X1 U2353 ( .IN1(\i_m4stg_frac/n901 ), .IN2(\i_m4stg_frac/n747 ), .IN3(
        \i_m4stg_frac/n434 ), .Q(n2684) );
  XNOR3X1 U2354 ( .IN1(n2698), .IN2(n2699), .IN3(n2700), .Q(n2686) );
  AOI22X1 U2355 ( .IN1(n2689), .IN2(n2688), .IN3(n2690), .IN4(n2701), .QN(
        n2685) );
  OR2X1 U2356 ( .IN1(n2688), .IN2(n2689), .Q(n2701) );
  XOR3X1 U2357 ( .IN1(\i_m4stg_frac/ps[79] ), .IN2(\i_m4stg_frac/pc[78] ), 
        .IN3(n1092), .Q(n2690) );
  AO22X1 U2358 ( .IN1(\i_m4stg_frac/pc[77] ), .IN2(n1091), .IN3(
        \i_m4stg_frac/ps[78] ), .IN4(n2702), .Q(n2688) );
  OR2X1 U2359 ( .IN1(n1091), .IN2(\i_m4stg_frac/pc[77] ), .Q(n2702) );
  OAI22X1 U2360 ( .IN1(\i_m4stg_frac/n438 ), .IN2(\i_m4stg_frac/n751 ), .IN3(
        n2703), .IN4(\i_m4stg_frac/n905 ), .QN(n2689) );
  AND2X1 U2361 ( .IN1(\i_m4stg_frac/n751 ), .IN2(\i_m4stg_frac/n438 ), .Q(
        n2703) );
  NOR2X0 U2362 ( .IN1(se_mul64), .IN2(n2044), .QN(\i_m4stg_frac/n403 ) );
  XNOR2X1 U2363 ( .IN1(n2168), .IN2(n2167), .Q(n2044) );
  XOR3X1 U2364 ( .IN1(n2704), .IN2(n2705), .IN3(n2706), .Q(n2167) );
  AO22X1 U2365 ( .IN1(n2695), .IN2(n2696), .IN3(n2694), .IN4(n2707), .Q(n2168)
         );
  OR2X1 U2366 ( .IN1(n2696), .IN2(n2695), .Q(n2707) );
  XOR3X1 U2367 ( .IN1(\i_m4stg_frac/n899 ), .IN2(\i_m4stg_frac/n745 ), .IN3(
        \i_m4stg_frac/n432 ), .Q(n2694) );
  XNOR3X1 U2368 ( .IN1(n2708), .IN2(n2709), .IN3(n2710), .Q(n2696) );
  AOI22X1 U2369 ( .IN1(n2699), .IN2(n2698), .IN3(n2700), .IN4(n2711), .QN(
        n2695) );
  OR2X1 U2370 ( .IN1(n2698), .IN2(n2699), .Q(n2711) );
  XOR3X1 U2371 ( .IN1(\i_m4stg_frac/ps[80] ), .IN2(\i_m4stg_frac/pc[79] ), 
        .IN3(n1093), .Q(n2700) );
  AO22X1 U2372 ( .IN1(\i_m4stg_frac/pc[78] ), .IN2(n1092), .IN3(
        \i_m4stg_frac/ps[79] ), .IN4(n2712), .Q(n2698) );
  OR2X1 U2373 ( .IN1(n1092), .IN2(\i_m4stg_frac/pc[78] ), .Q(n2712) );
  OAI22X1 U2374 ( .IN1(\i_m4stg_frac/n436 ), .IN2(\i_m4stg_frac/n749 ), .IN3(
        n2713), .IN4(\i_m4stg_frac/n903 ), .QN(n2699) );
  AND2X1 U2375 ( .IN1(\i_m4stg_frac/n749 ), .IN2(\i_m4stg_frac/n436 ), .Q(
        n2713) );
  NOR2X0 U2376 ( .IN1(se_mul64), .IN2(n2043), .QN(\i_m4stg_frac/n401 ) );
  XNOR2X1 U2377 ( .IN1(n2166), .IN2(n2165), .Q(n2043) );
  XOR3X1 U2378 ( .IN1(n2714), .IN2(n2715), .IN3(n2716), .Q(n2165) );
  AO22X1 U2379 ( .IN1(n2705), .IN2(n2706), .IN3(n2704), .IN4(n2717), .Q(n2166)
         );
  OR2X1 U2380 ( .IN1(n2706), .IN2(n2705), .Q(n2717) );
  XOR3X1 U2381 ( .IN1(\i_m4stg_frac/n897 ), .IN2(\i_m4stg_frac/n743 ), .IN3(
        \i_m4stg_frac/n430 ), .Q(n2704) );
  XNOR3X1 U2382 ( .IN1(n2718), .IN2(n2719), .IN3(n2720), .Q(n2706) );
  AOI22X1 U2383 ( .IN1(n2709), .IN2(n2708), .IN3(n2710), .IN4(n2721), .QN(
        n2705) );
  OR2X1 U2384 ( .IN1(n2708), .IN2(n2709), .Q(n2721) );
  XOR3X1 U2385 ( .IN1(\i_m4stg_frac/ps[81] ), .IN2(\i_m4stg_frac/pc[80] ), 
        .IN3(n1094), .Q(n2710) );
  AO22X1 U2386 ( .IN1(\i_m4stg_frac/pc[79] ), .IN2(n1093), .IN3(
        \i_m4stg_frac/ps[80] ), .IN4(n2722), .Q(n2708) );
  OR2X1 U2387 ( .IN1(n1093), .IN2(\i_m4stg_frac/pc[79] ), .Q(n2722) );
  OAI22X1 U2388 ( .IN1(\i_m4stg_frac/n434 ), .IN2(\i_m4stg_frac/n747 ), .IN3(
        n2723), .IN4(\i_m4stg_frac/n901 ), .QN(n2709) );
  AND2X1 U2389 ( .IN1(\i_m4stg_frac/n747 ), .IN2(\i_m4stg_frac/n434 ), .Q(
        n2723) );
  NOR2X0 U2390 ( .IN1(se_mul64), .IN2(n2042), .QN(\i_m4stg_frac/n399 ) );
  XNOR2X1 U2391 ( .IN1(n2164), .IN2(n2163), .Q(n2042) );
  XOR3X1 U2392 ( .IN1(n2724), .IN2(n2725), .IN3(n2726), .Q(n2163) );
  AO22X1 U2393 ( .IN1(n2715), .IN2(n2716), .IN3(n2714), .IN4(n2727), .Q(n2164)
         );
  OR2X1 U2394 ( .IN1(n2716), .IN2(n2715), .Q(n2727) );
  XOR3X1 U2395 ( .IN1(\i_m4stg_frac/n895 ), .IN2(\i_m4stg_frac/n741 ), .IN3(
        \i_m4stg_frac/n428 ), .Q(n2714) );
  XNOR3X1 U2396 ( .IN1(n2728), .IN2(n2729), .IN3(n2730), .Q(n2716) );
  AOI22X1 U2397 ( .IN1(n2719), .IN2(n2718), .IN3(n2720), .IN4(n2731), .QN(
        n2715) );
  OR2X1 U2398 ( .IN1(n2718), .IN2(n2719), .Q(n2731) );
  XOR3X1 U2399 ( .IN1(\i_m4stg_frac/ps[82] ), .IN2(\i_m4stg_frac/pc[81] ), 
        .IN3(n1095), .Q(n2720) );
  AO22X1 U2400 ( .IN1(\i_m4stg_frac/pc[80] ), .IN2(n1094), .IN3(
        \i_m4stg_frac/ps[81] ), .IN4(n2732), .Q(n2718) );
  OR2X1 U2401 ( .IN1(n1094), .IN2(\i_m4stg_frac/pc[80] ), .Q(n2732) );
  OAI22X1 U2402 ( .IN1(\i_m4stg_frac/n432 ), .IN2(\i_m4stg_frac/n745 ), .IN3(
        n2733), .IN4(\i_m4stg_frac/n899 ), .QN(n2719) );
  AND2X1 U2403 ( .IN1(\i_m4stg_frac/n745 ), .IN2(\i_m4stg_frac/n432 ), .Q(
        n2733) );
  NOR2X0 U2404 ( .IN1(se_mul64), .IN2(n2041), .QN(\i_m4stg_frac/n397 ) );
  XNOR2X1 U2405 ( .IN1(n2162), .IN2(n2161), .Q(n2041) );
  XOR3X1 U2406 ( .IN1(n2734), .IN2(n2735), .IN3(n2736), .Q(n2161) );
  AO22X1 U2407 ( .IN1(n2725), .IN2(n2726), .IN3(n2724), .IN4(n2737), .Q(n2162)
         );
  OR2X1 U2408 ( .IN1(n2726), .IN2(n2725), .Q(n2737) );
  XOR3X1 U2409 ( .IN1(\i_m4stg_frac/n893 ), .IN2(\i_m4stg_frac/n739 ), .IN3(
        \i_m4stg_frac/n426 ), .Q(n2724) );
  XNOR3X1 U2410 ( .IN1(n2738), .IN2(n2739), .IN3(n2740), .Q(n2726) );
  AOI22X1 U2411 ( .IN1(n2729), .IN2(n2728), .IN3(n2730), .IN4(n2741), .QN(
        n2725) );
  OR2X1 U2412 ( .IN1(n2728), .IN2(n2729), .Q(n2741) );
  XOR3X1 U2413 ( .IN1(\i_m4stg_frac/ps[83] ), .IN2(\i_m4stg_frac/pc[82] ), 
        .IN3(n1096), .Q(n2730) );
  AO22X1 U2414 ( .IN1(\i_m4stg_frac/pc[81] ), .IN2(n1095), .IN3(
        \i_m4stg_frac/ps[82] ), .IN4(n2742), .Q(n2728) );
  OR2X1 U2415 ( .IN1(n1095), .IN2(\i_m4stg_frac/pc[81] ), .Q(n2742) );
  OAI22X1 U2416 ( .IN1(\i_m4stg_frac/n430 ), .IN2(\i_m4stg_frac/n743 ), .IN3(
        n2743), .IN4(\i_m4stg_frac/n897 ), .QN(n2729) );
  AND2X1 U2417 ( .IN1(\i_m4stg_frac/n743 ), .IN2(\i_m4stg_frac/n430 ), .Q(
        n2743) );
  NOR2X0 U2418 ( .IN1(se_mul64), .IN2(n2040), .QN(\i_m4stg_frac/n395 ) );
  XNOR2X1 U2419 ( .IN1(n2160), .IN2(n2159), .Q(n2040) );
  XOR3X1 U2420 ( .IN1(n2744), .IN2(n2745), .IN3(n2746), .Q(n2159) );
  AO22X1 U2421 ( .IN1(n2735), .IN2(n2736), .IN3(n2734), .IN4(n2747), .Q(n2160)
         );
  OR2X1 U2422 ( .IN1(n2736), .IN2(n2735), .Q(n2747) );
  XOR3X1 U2423 ( .IN1(\i_m4stg_frac/n891 ), .IN2(\i_m4stg_frac/n737 ), .IN3(
        \i_m4stg_frac/n424 ), .Q(n2734) );
  XNOR3X1 U2424 ( .IN1(n2748), .IN2(n2749), .IN3(n2750), .Q(n2736) );
  AOI22X1 U2425 ( .IN1(n2739), .IN2(n2738), .IN3(n2740), .IN4(n2751), .QN(
        n2735) );
  OR2X1 U2426 ( .IN1(n2738), .IN2(n2739), .Q(n2751) );
  XOR3X1 U2427 ( .IN1(\i_m4stg_frac/ps[84] ), .IN2(\i_m4stg_frac/pc[83] ), 
        .IN3(n1097), .Q(n2740) );
  AO22X1 U2428 ( .IN1(\i_m4stg_frac/pc[82] ), .IN2(n1096), .IN3(
        \i_m4stg_frac/ps[83] ), .IN4(n2752), .Q(n2738) );
  OR2X1 U2429 ( .IN1(n1096), .IN2(\i_m4stg_frac/pc[82] ), .Q(n2752) );
  OAI22X1 U2430 ( .IN1(\i_m4stg_frac/n428 ), .IN2(\i_m4stg_frac/n741 ), .IN3(
        n2753), .IN4(\i_m4stg_frac/n895 ), .QN(n2739) );
  AND2X1 U2431 ( .IN1(\i_m4stg_frac/n741 ), .IN2(\i_m4stg_frac/n428 ), .Q(
        n2753) );
  NOR2X0 U2432 ( .IN1(se_mul64), .IN2(n2039), .QN(\i_m4stg_frac/n393 ) );
  XNOR2X1 U2433 ( .IN1(n2158), .IN2(n2157), .Q(n2039) );
  XOR3X1 U2434 ( .IN1(n2754), .IN2(n2755), .IN3(n2756), .Q(n2157) );
  AO22X1 U2435 ( .IN1(n2745), .IN2(n2746), .IN3(n2744), .IN4(n2757), .Q(n2158)
         );
  OR2X1 U2436 ( .IN1(n2746), .IN2(n2745), .Q(n2757) );
  XOR3X1 U2437 ( .IN1(\i_m4stg_frac/n889 ), .IN2(\i_m4stg_frac/n735 ), .IN3(
        \i_m4stg_frac/n422 ), .Q(n2744) );
  XNOR3X1 U2438 ( .IN1(n2758), .IN2(n2759), .IN3(n2760), .Q(n2746) );
  AOI22X1 U2439 ( .IN1(n2749), .IN2(n2748), .IN3(n2750), .IN4(n2761), .QN(
        n2745) );
  OR2X1 U2440 ( .IN1(n2748), .IN2(n2749), .Q(n2761) );
  XOR3X1 U2441 ( .IN1(\i_m4stg_frac/ps[85] ), .IN2(\i_m4stg_frac/pc[84] ), 
        .IN3(n1098), .Q(n2750) );
  AO22X1 U2442 ( .IN1(\i_m4stg_frac/pc[83] ), .IN2(n1097), .IN3(
        \i_m4stg_frac/ps[84] ), .IN4(n2762), .Q(n2748) );
  OR2X1 U2443 ( .IN1(n1097), .IN2(\i_m4stg_frac/pc[83] ), .Q(n2762) );
  OAI22X1 U2444 ( .IN1(\i_m4stg_frac/n426 ), .IN2(\i_m4stg_frac/n739 ), .IN3(
        n2763), .IN4(\i_m4stg_frac/n893 ), .QN(n2749) );
  AND2X1 U2445 ( .IN1(\i_m4stg_frac/n739 ), .IN2(\i_m4stg_frac/n426 ), .Q(
        n2763) );
  NOR2X0 U2446 ( .IN1(se_mul64), .IN2(n2038), .QN(\i_m4stg_frac/n391 ) );
  XNOR2X1 U2447 ( .IN1(n2156), .IN2(n2155), .Q(n2038) );
  XOR3X1 U2448 ( .IN1(n2764), .IN2(n2765), .IN3(n2766), .Q(n2155) );
  AO22X1 U2449 ( .IN1(n2755), .IN2(n2756), .IN3(n2754), .IN4(n2767), .Q(n2156)
         );
  OR2X1 U2450 ( .IN1(n2756), .IN2(n2755), .Q(n2767) );
  XOR3X1 U2451 ( .IN1(\i_m4stg_frac/n887 ), .IN2(\i_m4stg_frac/n733 ), .IN3(
        \i_m4stg_frac/n420 ), .Q(n2754) );
  XNOR3X1 U2452 ( .IN1(n2768), .IN2(n2769), .IN3(n2770), .Q(n2756) );
  AOI22X1 U2453 ( .IN1(n2759), .IN2(n2758), .IN3(n2760), .IN4(n2771), .QN(
        n2755) );
  OR2X1 U2454 ( .IN1(n2758), .IN2(n2759), .Q(n2771) );
  XOR3X1 U2455 ( .IN1(\i_m4stg_frac/ps[86] ), .IN2(\i_m4stg_frac/pc[85] ), 
        .IN3(n1099), .Q(n2760) );
  AO22X1 U2456 ( .IN1(\i_m4stg_frac/pc[84] ), .IN2(n1098), .IN3(
        \i_m4stg_frac/ps[85] ), .IN4(n2772), .Q(n2758) );
  OR2X1 U2457 ( .IN1(n1098), .IN2(\i_m4stg_frac/pc[84] ), .Q(n2772) );
  OAI22X1 U2458 ( .IN1(\i_m4stg_frac/n424 ), .IN2(\i_m4stg_frac/n737 ), .IN3(
        n2773), .IN4(\i_m4stg_frac/n891 ), .QN(n2759) );
  AND2X1 U2459 ( .IN1(\i_m4stg_frac/n737 ), .IN2(\i_m4stg_frac/n424 ), .Q(
        n2773) );
  NOR2X0 U2460 ( .IN1(se_mul64), .IN2(n2037), .QN(\i_m4stg_frac/n389 ) );
  XNOR2X1 U2461 ( .IN1(n2154), .IN2(n2153), .Q(n2037) );
  XOR3X1 U2462 ( .IN1(n2774), .IN2(n2775), .IN3(n2776), .Q(n2153) );
  AO22X1 U2463 ( .IN1(n2765), .IN2(n2766), .IN3(n2764), .IN4(n2777), .Q(n2154)
         );
  OR2X1 U2464 ( .IN1(n2766), .IN2(n2765), .Q(n2777) );
  XOR3X1 U2465 ( .IN1(\i_m4stg_frac/n885 ), .IN2(\i_m4stg_frac/n731 ), .IN3(
        \i_m4stg_frac/n418 ), .Q(n2764) );
  XNOR3X1 U2466 ( .IN1(n2778), .IN2(n2779), .IN3(n2780), .Q(n2766) );
  AOI22X1 U2467 ( .IN1(n2769), .IN2(n2768), .IN3(n2770), .IN4(n2781), .QN(
        n2765) );
  OR2X1 U2468 ( .IN1(n2768), .IN2(n2769), .Q(n2781) );
  XOR3X1 U2469 ( .IN1(\i_m4stg_frac/ps[87] ), .IN2(\i_m4stg_frac/pc[86] ), 
        .IN3(n1100), .Q(n2770) );
  AO22X1 U2470 ( .IN1(\i_m4stg_frac/pc[85] ), .IN2(n1099), .IN3(
        \i_m4stg_frac/ps[86] ), .IN4(n2782), .Q(n2768) );
  OR2X1 U2471 ( .IN1(n1099), .IN2(\i_m4stg_frac/pc[85] ), .Q(n2782) );
  OAI22X1 U2472 ( .IN1(\i_m4stg_frac/n422 ), .IN2(\i_m4stg_frac/n735 ), .IN3(
        n2783), .IN4(\i_m4stg_frac/n889 ), .QN(n2769) );
  AND2X1 U2473 ( .IN1(\i_m4stg_frac/n735 ), .IN2(\i_m4stg_frac/n422 ), .Q(
        n2783) );
  NOR2X0 U2474 ( .IN1(se_mul64), .IN2(n2036), .QN(\i_m4stg_frac/n387 ) );
  XNOR2X1 U2475 ( .IN1(n2152), .IN2(n2151), .Q(n2036) );
  XOR3X1 U2476 ( .IN1(n2784), .IN2(n2785), .IN3(n2786), .Q(n2151) );
  AO22X1 U2477 ( .IN1(n2775), .IN2(n2776), .IN3(n2774), .IN4(n2787), .Q(n2152)
         );
  OR2X1 U2478 ( .IN1(n2776), .IN2(n2775), .Q(n2787) );
  XOR3X1 U2479 ( .IN1(\i_m4stg_frac/n883 ), .IN2(\i_m4stg_frac/n729 ), .IN3(
        \i_m4stg_frac/n416 ), .Q(n2774) );
  XNOR3X1 U2480 ( .IN1(n2788), .IN2(n2789), .IN3(n2790), .Q(n2776) );
  AOI22X1 U2481 ( .IN1(n2779), .IN2(n2778), .IN3(n2780), .IN4(n2791), .QN(
        n2775) );
  OR2X1 U2482 ( .IN1(n2778), .IN2(n2779), .Q(n2791) );
  XOR3X1 U2483 ( .IN1(\i_m4stg_frac/ps[88] ), .IN2(\i_m4stg_frac/pc[87] ), 
        .IN3(n1101), .Q(n2780) );
  AO22X1 U2484 ( .IN1(\i_m4stg_frac/pc[86] ), .IN2(n1100), .IN3(
        \i_m4stg_frac/ps[87] ), .IN4(n2792), .Q(n2778) );
  OR2X1 U2485 ( .IN1(n1100), .IN2(\i_m4stg_frac/pc[86] ), .Q(n2792) );
  OAI22X1 U2486 ( .IN1(\i_m4stg_frac/n420 ), .IN2(\i_m4stg_frac/n733 ), .IN3(
        n2793), .IN4(\i_m4stg_frac/n887 ), .QN(n2779) );
  AND2X1 U2487 ( .IN1(\i_m4stg_frac/n733 ), .IN2(\i_m4stg_frac/n420 ), .Q(
        n2793) );
  NOR2X0 U2488 ( .IN1(se_mul64), .IN2(n2035), .QN(\i_m4stg_frac/n385 ) );
  XNOR2X1 U2489 ( .IN1(n2150), .IN2(n2149), .Q(n2035) );
  XOR3X1 U2490 ( .IN1(n2794), .IN2(n2795), .IN3(n2796), .Q(n2149) );
  AO22X1 U2491 ( .IN1(n2785), .IN2(n2786), .IN3(n2784), .IN4(n2797), .Q(n2150)
         );
  OR2X1 U2492 ( .IN1(n2786), .IN2(n2785), .Q(n2797) );
  XOR3X1 U2493 ( .IN1(\i_m4stg_frac/n881 ), .IN2(\i_m4stg_frac/n727 ), .IN3(
        \i_m4stg_frac/n414 ), .Q(n2784) );
  XNOR3X1 U2494 ( .IN1(n2798), .IN2(n2799), .IN3(n2800), .Q(n2786) );
  AOI22X1 U2495 ( .IN1(n2789), .IN2(n2788), .IN3(n2790), .IN4(n2801), .QN(
        n2785) );
  OR2X1 U2496 ( .IN1(n2788), .IN2(n2789), .Q(n2801) );
  XOR3X1 U2497 ( .IN1(\i_m4stg_frac/ps[89] ), .IN2(\i_m4stg_frac/pc[88] ), 
        .IN3(n1102), .Q(n2790) );
  AO22X1 U2498 ( .IN1(\i_m4stg_frac/pc[87] ), .IN2(n1101), .IN3(
        \i_m4stg_frac/ps[88] ), .IN4(n2802), .Q(n2788) );
  OR2X1 U2499 ( .IN1(n1101), .IN2(\i_m4stg_frac/pc[87] ), .Q(n2802) );
  OAI22X1 U2500 ( .IN1(\i_m4stg_frac/n418 ), .IN2(\i_m4stg_frac/n731 ), .IN3(
        n2803), .IN4(\i_m4stg_frac/n885 ), .QN(n2789) );
  AND2X1 U2501 ( .IN1(\i_m4stg_frac/n731 ), .IN2(\i_m4stg_frac/n418 ), .Q(
        n2803) );
  NOR2X0 U2502 ( .IN1(se_mul64), .IN2(n2034), .QN(\i_m4stg_frac/n383 ) );
  XNOR2X1 U2503 ( .IN1(n2148), .IN2(n2147), .Q(n2034) );
  XOR3X1 U2504 ( .IN1(n2804), .IN2(n2805), .IN3(n2806), .Q(n2147) );
  AO22X1 U2505 ( .IN1(n2795), .IN2(n2796), .IN3(n2794), .IN4(n2807), .Q(n2148)
         );
  OR2X1 U2506 ( .IN1(n2796), .IN2(n2795), .Q(n2807) );
  XOR3X1 U2507 ( .IN1(\i_m4stg_frac/n879 ), .IN2(\i_m4stg_frac/n725 ), .IN3(
        \i_m4stg_frac/n412 ), .Q(n2794) );
  XNOR3X1 U2508 ( .IN1(n2808), .IN2(n2809), .IN3(n2810), .Q(n2796) );
  AOI22X1 U2509 ( .IN1(n2799), .IN2(n2798), .IN3(n2800), .IN4(n2811), .QN(
        n2795) );
  OR2X1 U2510 ( .IN1(n2798), .IN2(n2799), .Q(n2811) );
  XOR3X1 U2511 ( .IN1(\i_m4stg_frac/ps[90] ), .IN2(\i_m4stg_frac/pc[89] ), 
        .IN3(n1103), .Q(n2800) );
  AO22X1 U2512 ( .IN1(\i_m4stg_frac/pc[88] ), .IN2(n1102), .IN3(
        \i_m4stg_frac/ps[89] ), .IN4(n2812), .Q(n2798) );
  OR2X1 U2513 ( .IN1(n1102), .IN2(\i_m4stg_frac/pc[88] ), .Q(n2812) );
  OAI22X1 U2514 ( .IN1(\i_m4stg_frac/n416 ), .IN2(\i_m4stg_frac/n729 ), .IN3(
        n2813), .IN4(\i_m4stg_frac/n883 ), .QN(n2799) );
  AND2X1 U2515 ( .IN1(\i_m4stg_frac/n729 ), .IN2(\i_m4stg_frac/n416 ), .Q(
        n2813) );
  NOR2X0 U2516 ( .IN1(se_mul64), .IN2(n2033), .QN(\i_m4stg_frac/n381 ) );
  XNOR2X1 U2517 ( .IN1(n2146), .IN2(n2145), .Q(n2033) );
  XOR3X1 U2518 ( .IN1(n2814), .IN2(n2815), .IN3(n2816), .Q(n2145) );
  AO22X1 U2519 ( .IN1(n2805), .IN2(n2806), .IN3(n2804), .IN4(n2817), .Q(n2146)
         );
  OR2X1 U2520 ( .IN1(n2806), .IN2(n2805), .Q(n2817) );
  XOR3X1 U2521 ( .IN1(\i_m4stg_frac/n877 ), .IN2(\i_m4stg_frac/n723 ), .IN3(
        \i_m4stg_frac/n410 ), .Q(n2804) );
  XNOR3X1 U2522 ( .IN1(n2818), .IN2(n2819), .IN3(n2820), .Q(n2806) );
  AOI22X1 U2523 ( .IN1(n2809), .IN2(n2808), .IN3(n2810), .IN4(n2821), .QN(
        n2805) );
  OR2X1 U2524 ( .IN1(n2808), .IN2(n2809), .Q(n2821) );
  XOR3X1 U2525 ( .IN1(\i_m4stg_frac/ps[91] ), .IN2(\i_m4stg_frac/pc[90] ), 
        .IN3(n1104), .Q(n2810) );
  AO22X1 U2526 ( .IN1(\i_m4stg_frac/pc[89] ), .IN2(n1103), .IN3(
        \i_m4stg_frac/ps[90] ), .IN4(n2822), .Q(n2808) );
  OR2X1 U2527 ( .IN1(n1103), .IN2(\i_m4stg_frac/pc[89] ), .Q(n2822) );
  OAI22X1 U2528 ( .IN1(\i_m4stg_frac/n414 ), .IN2(\i_m4stg_frac/n727 ), .IN3(
        n2823), .IN4(\i_m4stg_frac/n881 ), .QN(n2809) );
  AND2X1 U2529 ( .IN1(\i_m4stg_frac/n727 ), .IN2(\i_m4stg_frac/n414 ), .Q(
        n2823) );
  NOR2X0 U2530 ( .IN1(se_mul64), .IN2(n2032), .QN(\i_m4stg_frac/n379 ) );
  XNOR2X1 U2531 ( .IN1(n2144), .IN2(n2143), .Q(n2032) );
  XOR3X1 U2532 ( .IN1(n2824), .IN2(n2825), .IN3(n2826), .Q(n2143) );
  AO22X1 U2533 ( .IN1(n2815), .IN2(n2816), .IN3(n2814), .IN4(n2827), .Q(n2144)
         );
  OR2X1 U2534 ( .IN1(n2816), .IN2(n2815), .Q(n2827) );
  XOR3X1 U2535 ( .IN1(\i_m4stg_frac/n875 ), .IN2(\i_m4stg_frac/n721 ), .IN3(
        \i_m4stg_frac/n408 ), .Q(n2814) );
  XNOR3X1 U2536 ( .IN1(n2828), .IN2(n2829), .IN3(n2830), .Q(n2816) );
  AOI22X1 U2537 ( .IN1(n2819), .IN2(n2818), .IN3(n2820), .IN4(n2831), .QN(
        n2815) );
  OR2X1 U2538 ( .IN1(n2818), .IN2(n2819), .Q(n2831) );
  XOR3X1 U2539 ( .IN1(\i_m4stg_frac/ps[92] ), .IN2(\i_m4stg_frac/pc[91] ), 
        .IN3(n1105), .Q(n2820) );
  AO22X1 U2540 ( .IN1(\i_m4stg_frac/pc[90] ), .IN2(n1104), .IN3(
        \i_m4stg_frac/ps[91] ), .IN4(n2832), .Q(n2818) );
  OR2X1 U2541 ( .IN1(n1104), .IN2(\i_m4stg_frac/pc[90] ), .Q(n2832) );
  OAI22X1 U2542 ( .IN1(\i_m4stg_frac/n412 ), .IN2(\i_m4stg_frac/n725 ), .IN3(
        n2833), .IN4(\i_m4stg_frac/n879 ), .QN(n2819) );
  AND2X1 U2543 ( .IN1(\i_m4stg_frac/n725 ), .IN2(\i_m4stg_frac/n412 ), .Q(
        n2833) );
  NOR2X0 U2544 ( .IN1(se_mul64), .IN2(n2031), .QN(\i_m4stg_frac/n377 ) );
  XNOR2X1 U2545 ( .IN1(n2142), .IN2(n2141), .Q(n2031) );
  XOR3X1 U2546 ( .IN1(n2834), .IN2(n2835), .IN3(n2836), .Q(n2141) );
  AO22X1 U2547 ( .IN1(n2825), .IN2(n2826), .IN3(n2824), .IN4(n2837), .Q(n2142)
         );
  OR2X1 U2548 ( .IN1(n2826), .IN2(n2825), .Q(n2837) );
  XOR3X1 U2549 ( .IN1(\i_m4stg_frac/n873 ), .IN2(\i_m4stg_frac/n719 ), .IN3(
        \i_m4stg_frac/n406 ), .Q(n2824) );
  XNOR3X1 U2550 ( .IN1(n2838), .IN2(n2839), .IN3(n2840), .Q(n2826) );
  AOI22X1 U2551 ( .IN1(n2829), .IN2(n2828), .IN3(n2830), .IN4(n2841), .QN(
        n2825) );
  OR2X1 U2552 ( .IN1(n2828), .IN2(n2829), .Q(n2841) );
  XOR3X1 U2553 ( .IN1(\i_m4stg_frac/ps[93] ), .IN2(\i_m4stg_frac/pc[92] ), 
        .IN3(n1106), .Q(n2830) );
  AO22X1 U2554 ( .IN1(\i_m4stg_frac/pc[91] ), .IN2(n1105), .IN3(
        \i_m4stg_frac/ps[92] ), .IN4(n2842), .Q(n2828) );
  OR2X1 U2555 ( .IN1(n1105), .IN2(\i_m4stg_frac/pc[91] ), .Q(n2842) );
  OAI22X1 U2556 ( .IN1(\i_m4stg_frac/n410 ), .IN2(\i_m4stg_frac/n723 ), .IN3(
        n2843), .IN4(\i_m4stg_frac/n877 ), .QN(n2829) );
  AND2X1 U2557 ( .IN1(\i_m4stg_frac/n723 ), .IN2(\i_m4stg_frac/n410 ), .Q(
        n2843) );
  NOR2X0 U2558 ( .IN1(se_mul64), .IN2(n2030), .QN(\i_m4stg_frac/n375 ) );
  XNOR2X1 U2559 ( .IN1(n2140), .IN2(n2139), .Q(n2030) );
  XOR3X1 U2560 ( .IN1(n2844), .IN2(n2845), .IN3(n2846), .Q(n2139) );
  AO22X1 U2561 ( .IN1(n2835), .IN2(n2836), .IN3(n2834), .IN4(n2847), .Q(n2140)
         );
  OR2X1 U2562 ( .IN1(n2836), .IN2(n2835), .Q(n2847) );
  XOR3X1 U2563 ( .IN1(\i_m4stg_frac/n871 ), .IN2(\i_m4stg_frac/n717 ), .IN3(
        \i_m4stg_frac/n404 ), .Q(n2834) );
  XNOR3X1 U2564 ( .IN1(n2848), .IN2(n2849), .IN3(n2850), .Q(n2836) );
  AOI22X1 U2565 ( .IN1(n2839), .IN2(n2838), .IN3(n2840), .IN4(n2851), .QN(
        n2835) );
  OR2X1 U2566 ( .IN1(n2838), .IN2(n2839), .Q(n2851) );
  XOR3X1 U2567 ( .IN1(\i_m4stg_frac/ps[94] ), .IN2(\i_m4stg_frac/pc[93] ), 
        .IN3(n1107), .Q(n2840) );
  AO22X1 U2568 ( .IN1(\i_m4stg_frac/pc[92] ), .IN2(n1106), .IN3(
        \i_m4stg_frac/ps[93] ), .IN4(n2852), .Q(n2838) );
  OR2X1 U2569 ( .IN1(n1106), .IN2(\i_m4stg_frac/pc[92] ), .Q(n2852) );
  OAI22X1 U2570 ( .IN1(\i_m4stg_frac/n408 ), .IN2(\i_m4stg_frac/n721 ), .IN3(
        n2853), .IN4(\i_m4stg_frac/n875 ), .QN(n2839) );
  AND2X1 U2571 ( .IN1(\i_m4stg_frac/n721 ), .IN2(\i_m4stg_frac/n408 ), .Q(
        n2853) );
  NOR2X0 U2572 ( .IN1(se_mul64), .IN2(n2029), .QN(\i_m4stg_frac/n373 ) );
  XNOR2X1 U2573 ( .IN1(n2138), .IN2(n2137), .Q(n2029) );
  XOR3X1 U2574 ( .IN1(n2854), .IN2(n2855), .IN3(n2856), .Q(n2137) );
  AO22X1 U2575 ( .IN1(n2845), .IN2(n2846), .IN3(n2844), .IN4(n2857), .Q(n2138)
         );
  OR2X1 U2576 ( .IN1(n2846), .IN2(n2845), .Q(n2857) );
  XOR3X1 U2577 ( .IN1(\i_m4stg_frac/n869 ), .IN2(\i_m4stg_frac/n715 ), .IN3(
        \i_m4stg_frac/n402 ), .Q(n2844) );
  XNOR3X1 U2578 ( .IN1(n2858), .IN2(n2859), .IN3(n2860), .Q(n2846) );
  AOI22X1 U2579 ( .IN1(n2849), .IN2(n2848), .IN3(n2850), .IN4(n2861), .QN(
        n2845) );
  OR2X1 U2580 ( .IN1(n2848), .IN2(n2849), .Q(n2861) );
  XOR3X1 U2581 ( .IN1(\i_m4stg_frac/ps[95] ), .IN2(\i_m4stg_frac/pc[94] ), 
        .IN3(n1108), .Q(n2850) );
  AO22X1 U2582 ( .IN1(\i_m4stg_frac/pc[93] ), .IN2(n1107), .IN3(
        \i_m4stg_frac/ps[94] ), .IN4(n2862), .Q(n2848) );
  OR2X1 U2583 ( .IN1(n1107), .IN2(\i_m4stg_frac/pc[93] ), .Q(n2862) );
  OAI22X1 U2584 ( .IN1(\i_m4stg_frac/n406 ), .IN2(\i_m4stg_frac/n719 ), .IN3(
        n2863), .IN4(\i_m4stg_frac/n873 ), .QN(n2849) );
  AND2X1 U2585 ( .IN1(\i_m4stg_frac/n719 ), .IN2(\i_m4stg_frac/n406 ), .Q(
        n2863) );
  NOR2X0 U2586 ( .IN1(se_mul64), .IN2(n2028), .QN(\i_m4stg_frac/n371 ) );
  XNOR2X1 U2587 ( .IN1(n2136), .IN2(n2135), .Q(n2028) );
  XOR3X1 U2588 ( .IN1(n2864), .IN2(n2865), .IN3(n2866), .Q(n2135) );
  AO22X1 U2589 ( .IN1(n2855), .IN2(n2856), .IN3(n2854), .IN4(n2867), .Q(n2136)
         );
  OR2X1 U2590 ( .IN1(n2856), .IN2(n2855), .Q(n2867) );
  XOR3X1 U2591 ( .IN1(\i_m4stg_frac/n867 ), .IN2(\i_m4stg_frac/n713 ), .IN3(
        \i_m4stg_frac/n400 ), .Q(n2854) );
  XNOR3X1 U2592 ( .IN1(n2868), .IN2(n2869), .IN3(n2870), .Q(n2856) );
  AOI22X1 U2593 ( .IN1(n2859), .IN2(n2858), .IN3(n2860), .IN4(n2871), .QN(
        n2855) );
  OR2X1 U2594 ( .IN1(n2858), .IN2(n2859), .Q(n2871) );
  XOR3X1 U2595 ( .IN1(\i_m4stg_frac/ps[96] ), .IN2(\i_m4stg_frac/pc[95] ), 
        .IN3(n1109), .Q(n2860) );
  AO22X1 U2596 ( .IN1(\i_m4stg_frac/pc[94] ), .IN2(n1108), .IN3(
        \i_m4stg_frac/ps[95] ), .IN4(n2872), .Q(n2858) );
  OR2X1 U2597 ( .IN1(n1108), .IN2(\i_m4stg_frac/pc[94] ), .Q(n2872) );
  OAI22X1 U2598 ( .IN1(\i_m4stg_frac/n404 ), .IN2(\i_m4stg_frac/n717 ), .IN3(
        n2873), .IN4(\i_m4stg_frac/n871 ), .QN(n2859) );
  AND2X1 U2599 ( .IN1(\i_m4stg_frac/n717 ), .IN2(\i_m4stg_frac/n404 ), .Q(
        n2873) );
  NOR2X0 U2600 ( .IN1(se_mul64), .IN2(n2027), .QN(\i_m4stg_frac/n369 ) );
  XNOR2X1 U2601 ( .IN1(n2131), .IN2(n2132), .Q(n2027) );
  XOR3X1 U2602 ( .IN1(n2874), .IN2(n2875), .IN3(n2876), .Q(n2132) );
  OA22X1 U2603 ( .IN1(n2866), .IN2(n2865), .IN3(n2864), .IN4(n2877), .Q(n2131)
         );
  AND2X1 U2604 ( .IN1(n2865), .IN2(n2866), .Q(n2877) );
  XOR3X1 U2605 ( .IN1(\i_m4stg_frac/n865 ), .IN2(\i_m4stg_frac/n711 ), .IN3(
        \i_m4stg_frac/n398 ), .Q(n2864) );
  AOI22X1 U2606 ( .IN1(n2869), .IN2(n2868), .IN3(n2870), .IN4(n2878), .QN(
        n2865) );
  OR2X1 U2607 ( .IN1(n2868), .IN2(n2869), .Q(n2878) );
  XOR3X1 U2608 ( .IN1(\i_m4stg_frac/ps[97] ), .IN2(\i_m4stg_frac/pc[96] ), 
        .IN3(n1110), .Q(n2870) );
  AO22X1 U2609 ( .IN1(\i_m4stg_frac/pc[95] ), .IN2(n1109), .IN3(
        \i_m4stg_frac/ps[96] ), .IN4(n2879), .Q(n2868) );
  OR2X1 U2610 ( .IN1(n1109), .IN2(\i_m4stg_frac/pc[95] ), .Q(n2879) );
  OAI22X1 U2611 ( .IN1(\i_m4stg_frac/n402 ), .IN2(\i_m4stg_frac/n715 ), .IN3(
        n2880), .IN4(\i_m4stg_frac/n869 ), .QN(n2869) );
  AND2X1 U2612 ( .IN1(\i_m4stg_frac/n715 ), .IN2(\i_m4stg_frac/n402 ), .Q(
        n2880) );
  XNOR3X1 U2613 ( .IN1(n2881), .IN2(n2882), .IN3(n2883), .Q(n2866) );
  NOR2X0 U2614 ( .IN1(se_mul64), .IN2(n2025), .QN(\i_m4stg_frac/n367 ) );
  XOR2X1 U2615 ( .IN1(n2290), .IN2(n2130), .Q(n2025) );
  INVX0 U2616 ( .INP(n2289), .ZN(n2130) );
  AO22X1 U2617 ( .IN1(n2874), .IN2(n2876), .IN3(n2884), .IN4(n2875), .Q(n2289)
         );
  AO21X1 U2618 ( .IN1(n2885), .IN2(n2886), .IN3(n2514), .Q(n2875) );
  AO21X1 U2619 ( .IN1(\i_m4stg_frac/n396 ), .IN2(\i_m4stg_frac/n550 ), .IN3(
        n2521), .Q(n2885) );
  OR2X1 U2620 ( .IN1(n2876), .IN2(n2874), .Q(n2884) );
  OAI22X1 U2621 ( .IN1(n2881), .IN2(n2882), .IN3(n2883), .IN4(n2887), .QN(
        n2876) );
  AND2X1 U2622 ( .IN1(n2881), .IN2(n2882), .Q(n2887) );
  XOR3X1 U2623 ( .IN1(\i_m4stg_frac/ps[98] ), .IN2(\i_m4stg_frac/pc[97] ), 
        .IN3(n1111), .Q(n2883) );
  OAI22X1 U2624 ( .IN1(\i_m4stg_frac/n400 ), .IN2(\i_m4stg_frac/n713 ), .IN3(
        n2888), .IN4(\i_m4stg_frac/n867 ), .QN(n2882) );
  AND2X1 U2625 ( .IN1(\i_m4stg_frac/n713 ), .IN2(\i_m4stg_frac/n400 ), .Q(
        n2888) );
  AO22X1 U2626 ( .IN1(\i_m4stg_frac/pc[96] ), .IN2(n1110), .IN3(
        \i_m4stg_frac/ps[97] ), .IN4(n2889), .Q(n2881) );
  OR2X1 U2627 ( .IN1(n1110), .IN2(\i_m4stg_frac/pc[96] ), .Q(n2889) );
  XOR3X1 U2628 ( .IN1(\i_m4stg_frac/n863 ), .IN2(n928), .IN3(n2890), .Q(n2874)
         );
  INVX0 U2629 ( .INP(n2129), .ZN(n2290) );
  XOR3X1 U2630 ( .IN1(n2512), .IN2(n2514), .IN3(n2513), .Q(n2129) );
  AO22X1 U2631 ( .IN1(n2890), .IN2(n928), .IN3(n2891), .IN4(n1330), .Q(n2513)
         );
  OR2X1 U2632 ( .IN1(n928), .IN2(n2890), .Q(n2891) );
  AO22X1 U2633 ( .IN1(\i_m4stg_frac/pc[97] ), .IN2(n1111), .IN3(
        \i_m4stg_frac/ps[98] ), .IN4(n2892), .Q(n2890) );
  OR2X1 U2634 ( .IN1(n1111), .IN2(\i_m4stg_frac/pc[97] ), .Q(n2892) );
  NOR2X0 U2635 ( .IN1(n2886), .IN2(n2893), .QN(n2514) );
  XNOR2X1 U2636 ( .IN1(\i_m4stg_frac/n550 ), .IN2(\i_m4stg_frac/n396 ), .Q(
        n2893) );
  AO22X1 U2637 ( .IN1(\i_m4stg_frac/n711 ), .IN2(\i_m4stg_frac/n398 ), .IN3(
        \i_m4stg_frac/n865 ), .IN4(n2894), .Q(n2886) );
  OR2X1 U2638 ( .IN1(\i_m4stg_frac/n711 ), .IN2(\i_m4stg_frac/n398 ), .Q(n2894) );
  XOR3X1 U2639 ( .IN1(\i_m4stg_frac/n707 ), .IN2(n2521), .IN3(n2518), .Q(n2512) );
  NOR3X0 U2640 ( .IN1(n2234), .IN2(se_mul64), .IN3(n2238), .QN(
        \i_m4stg_frac/n365 ) );
  XNOR2X1 U2641 ( .IN1(n2242), .IN2(n2243), .Q(n2238) );
  NAND2X0 U2642 ( .IN1(n2235), .IN2(n2236), .QN(n2234) );
  AO22X1 U2643 ( .IN1(\i_m4stg_frac/pc[31] ), .IN2(n1185), .IN3(
        \i_m4stg_frac/ps[32] ), .IN4(n2895), .Q(n2236) );
  OR2X1 U2644 ( .IN1(n1185), .IN2(\i_m4stg_frac/pc[31] ), .Q(n2895) );
  XOR3X1 U2645 ( .IN1(\i_m4stg_frac/ps[33] ), .IN2(\i_m4stg_frac/pc[32] ), 
        .IN3(n1120), .Q(n2235) );
  NOR2X0 U2646 ( .IN1(se_mul64), .IN2(n2240), .QN(\i_m4stg_frac/n363 ) );
  NAND4X0 U2647 ( .IN1(n2242), .IN2(n2243), .IN3(n2241), .IN4(n2205), .QN(
        n2240) );
  INVX0 U2648 ( .INP(n2896), .ZN(n2205) );
  NAND2X0 U2649 ( .IN1(n2897), .IN2(n2898), .QN(n2241) );
  OA22X1 U2650 ( .IN1(n1120), .IN2(\i_m4stg_frac/pc[32] ), .IN3(n2899), .IN4(
        \i_m4stg_frac/ps[33] ), .Q(n2243) );
  AND2X1 U2651 ( .IN1(\i_m4stg_frac/pc[32] ), .IN2(n1120), .Q(n2899) );
  XOR3X1 U2652 ( .IN1(\i_m4stg_frac/ps[34] ), .IN2(\i_m4stg_frac/pc[33] ), 
        .IN3(n1125), .Q(n2242) );
  NOR2X0 U2653 ( .IN1(se_mul64), .IN2(n2202), .QN(\i_m4stg_frac/n361 ) );
  NAND3X0 U2654 ( .IN1(n2900), .IN2(n2500), .IN3(n2896), .QN(n2202) );
  NOR2X0 U2655 ( .IN1(n2898), .IN2(n2897), .QN(n2896) );
  XNOR3X1 U2656 ( .IN1(\i_m4stg_frac/ps[35] ), .IN2(\i_m4stg_frac/pc[34] ), 
        .IN3(n1131), .Q(n2897) );
  OAI22X1 U2657 ( .IN1(n1125), .IN2(\i_m4stg_frac/pc[33] ), .IN3(n2901), .IN4(
        \i_m4stg_frac/ps[34] ), .QN(n2898) );
  AND2X1 U2658 ( .IN1(\i_m4stg_frac/pc[33] ), .IN2(n1125), .Q(n2901) );
  INVX0 U2659 ( .INP(n2203), .ZN(n2500) );
  NOR2X0 U2660 ( .IN1(n2206), .IN2(n2207), .QN(n2203) );
  NAND2X0 U2661 ( .IN1(n2207), .IN2(n2206), .QN(n2900) );
  XOR3X1 U2662 ( .IN1(\i_m4stg_frac/ps[36] ), .IN2(\i_m4stg_frac/pc[35] ), 
        .IN3(\i_m4stg_frac/n989 ), .Q(n2206) );
  AOI22X1 U2663 ( .IN1(\i_m4stg_frac/pc[34] ), .IN2(n1131), .IN3(
        \i_m4stg_frac/ps[35] ), .IN4(n2902), .QN(n2207) );
  OR2X1 U2664 ( .IN1(n1131), .IN2(\i_m4stg_frac/pc[34] ), .Q(n2902) );
  NOR3X0 U2665 ( .IN1(n2127), .IN2(se_mul64), .IN3(n2126), .QN(
        \i_m4stg_frac/n359 ) );
  XNOR2X1 U2666 ( .IN1(n2211), .IN2(n2212), .Q(n2126) );
  AO221X1 U2667 ( .IN1(\i_m4stg_frac/n707 ), .IN2(n2903), .IN3(n2518), .IN4(
        n2517), .IN5(n2519), .Q(n2127) );
  XOR3X1 U2668 ( .IN1(\i_m4stg_frac/n705 ), .IN2(n2904), .IN3(n2905), .Q(n2519) );
  INVX0 U2669 ( .INP(n2521), .ZN(n2517) );
  INVX0 U2670 ( .INP(n2520), .ZN(n2518) );
  NAND2X0 U2671 ( .IN1(n2521), .IN2(n2520), .QN(n2903) );
  XNOR3X1 U2672 ( .IN1(\i_m4stg_frac/n861 ), .IN2(\i_m4stg_frac/n548 ), .IN3(
        \i_m4stg_frac/n394 ), .Q(n2520) );
  NOR2X0 U2673 ( .IN1(\i_m4stg_frac/n550 ), .IN2(\i_m4stg_frac/n396 ), .QN(
        n2521) );
  NOR2X0 U2674 ( .IN1(se_mul64), .IN2(n2125), .QN(\i_m4stg_frac/n357 ) );
  NAND4X0 U2675 ( .IN1(n2212), .IN2(n2211), .IN3(n2213), .IN4(n2214), .QN(
        n2125) );
  INVX0 U2676 ( .INP(n2906), .ZN(n2214) );
  NAND2X0 U2677 ( .IN1(n2907), .IN2(n2908), .QN(n2213) );
  AOI22X1 U2678 ( .IN1(n2904), .IN2(n2905), .IN3(\i_m4stg_frac/n705 ), .IN4(
        n2909), .QN(n2211) );
  OR2X1 U2679 ( .IN1(n2905), .IN2(n2904), .Q(n2909) );
  XOR3X1 U2680 ( .IN1(\i_m4stg_frac/n859 ), .IN2(\i_m4stg_frac/n546 ), .IN3(
        \i_m4stg_frac/n392 ), .Q(n2905) );
  OA22X1 U2681 ( .IN1(\i_m4stg_frac/n394 ), .IN2(\i_m4stg_frac/n548 ), .IN3(
        n2910), .IN4(\i_m4stg_frac/n861 ), .Q(n2904) );
  AND2X1 U2682 ( .IN1(\i_m4stg_frac/n548 ), .IN2(\i_m4stg_frac/n394 ), .Q(
        n2910) );
  XNOR3X1 U2683 ( .IN1(\i_m4stg_frac/n703 ), .IN2(n2911), .IN3(n2912), .Q(
        n2212) );
  NOR2X0 U2684 ( .IN1(se_mul64), .IN2(n2124), .QN(\i_m4stg_frac/n355 ) );
  NAND3X0 U2685 ( .IN1(n2913), .IN2(n2220), .IN3(n2906), .QN(n2124) );
  NOR2X0 U2686 ( .IN1(n2908), .IN2(n2907), .QN(n2906) );
  XOR3X1 U2687 ( .IN1(\i_m4stg_frac/n701 ), .IN2(n2914), .IN3(n2915), .Q(n2907) );
  AO22X1 U2688 ( .IN1(n2911), .IN2(n2912), .IN3(\i_m4stg_frac/n703 ), .IN4(
        n2916), .Q(n2908) );
  OR2X1 U2689 ( .IN1(n2912), .IN2(n2911), .Q(n2916) );
  XOR3X1 U2690 ( .IN1(\i_m4stg_frac/n857 ), .IN2(\i_m4stg_frac/n544 ), .IN3(
        \i_m4stg_frac/n390 ), .Q(n2912) );
  OA22X1 U2691 ( .IN1(\i_m4stg_frac/n392 ), .IN2(\i_m4stg_frac/n546 ), .IN3(
        n2917), .IN4(\i_m4stg_frac/n859 ), .Q(n2911) );
  AND2X1 U2692 ( .IN1(\i_m4stg_frac/n546 ), .IN2(\i_m4stg_frac/n392 ), .Q(
        n2917) );
  INVX0 U2693 ( .INP(n2219), .ZN(n2220) );
  NOR2X0 U2694 ( .IN1(n2218), .IN2(n2217), .QN(n2219) );
  NAND2X0 U2695 ( .IN1(n2217), .IN2(n2218), .QN(n2913) );
  AO22X1 U2696 ( .IN1(n2914), .IN2(n2915), .IN3(\i_m4stg_frac/n701 ), .IN4(
        n2918), .Q(n2218) );
  OR2X1 U2697 ( .IN1(n2915), .IN2(n2914), .Q(n2918) );
  XOR3X1 U2698 ( .IN1(\i_m4stg_frac/n855 ), .IN2(\i_m4stg_frac/n542 ), .IN3(
        \i_m4stg_frac/n388 ), .Q(n2915) );
  OA22X1 U2699 ( .IN1(\i_m4stg_frac/n390 ), .IN2(\i_m4stg_frac/n544 ), .IN3(
        n2919), .IN4(\i_m4stg_frac/n857 ), .Q(n2914) );
  AND2X1 U2700 ( .IN1(\i_m4stg_frac/n544 ), .IN2(\i_m4stg_frac/n390 ), .Q(
        n2919) );
  XOR3X1 U2701 ( .IN1(\i_m4stg_frac/n699 ), .IN2(n2226), .IN3(n2227), .Q(n2217) );
  XOR3X1 U2702 ( .IN1(\i_m4stg_frac/n853 ), .IN2(\i_m4stg_frac/n540 ), .IN3(
        \i_m4stg_frac/n386 ), .Q(n2227) );
  OA22X1 U2703 ( .IN1(\i_m4stg_frac/n388 ), .IN2(\i_m4stg_frac/n542 ), .IN3(
        n2920), .IN4(\i_m4stg_frac/n855 ), .Q(n2226) );
  AND2X1 U2704 ( .IN1(\i_m4stg_frac/n542 ), .IN2(\i_m4stg_frac/n388 ), .Q(
        n2920) );
  OA22X1 U2705 ( .IN1(n2921), .IN2(n2922), .IN3(n2923), .IN4(n2924), .Q(
        \i_m4stg_frac/n1693 ) );
  MUX21X1 U2706 ( .IN1(n2925), .IN2(n2926), .S(\i_m4stg_frac/n300 ), .Q(n2922)
         );
  NOR2X0 U2707 ( .IN1(\i_m4stg_frac/n345 ), .IN2(\i_m4stg_frac/n207 ), .QN(
        n2926) );
  AND2X1 U2708 ( .IN1(\i_m4stg_frac/n207 ), .IN2(\i_m4stg_frac/n345 ), .Q(
        n2925) );
  NOR2X0 U2709 ( .IN1(mul_rst_l), .IN2(n1375), .QN(\i_m4stg_frac/cyc3_dff/N7 )
         );
  NOR3X0 U2710 ( .IN1(\i_m4stg_frac/n1464 ), .IN2(se_mul64), .IN3(mul_rst_l), 
        .QN(\i_m4stg_frac/cyc2_dff/N7 ) );
  NOR2X0 U2711 ( .IN1(mul_rst_l), .IN2(n2924), .QN(\i_m4stg_frac/cyc1_dff/N7 )
         );
  NOR3X0 U2712 ( .IN1(n2927), .IN2(se_mul64), .IN3(\i_m4stg_frac/n1462 ), .QN(
        \i_m4stg_frac/co31_dff/N3 ) );
  AO21X1 U2713 ( .IN1(n2928), .IN2(n2929), .IN3(se_mul64), .Q(
        \i_m4stg_frac/ckbuf_1/N1 ) );
  NAND2X0 U2714 ( .IN1(n603), .IN2(\i_m4stg_frac/n854 ), .QN(
        \i_m4stg_frac/ckbuf_0/N1 ) );
  NAND2X0 U2715 ( .IN1(n2930), .IN2(n2931), .QN(
        \i_m4stg_frac/booth/out_dff9/N5 ) );
  OAI22X1 U2716 ( .IN1(n2932), .IN2(n2921), .IN3(n2933), .IN4(n2924), .QN(
        \i_m4stg_frac/booth/out_dff9/N4 ) );
  OA21X1 U2717 ( .IN1(n2934), .IN2(n2935), .IN3(n2936), .Q(n2933) );
  INVX0 U2718 ( .INP(n2937), .ZN(n2936) );
  MUX21X1 U2719 ( .IN1(n2934), .IN2(n2935), .S(n2938), .Q(n2937) );
  OA21X1 U2720 ( .IN1(\i_m4stg_frac/n334 ), .IN2(n1161), .IN3(n2939), .Q(n2932) );
  INVX0 U2721 ( .INP(n2940), .ZN(n2939) );
  MUX21X1 U2722 ( .IN1(n1161), .IN2(\i_m4stg_frac/n334 ), .S(
        \i_m4stg_frac/n201 ), .Q(n2940) );
  NAND2X0 U2723 ( .IN1(n2941), .IN2(n2942), .QN(
        \i_m4stg_frac/booth/out_dff9/N3 ) );
  MUX21X1 U2724 ( .IN1(n2943), .IN2(n2944), .S(\i_m4stg_frac/n334 ), .Q(n2942)
         );
  NAND2X0 U2725 ( .IN1(n2945), .IN2(n1172), .QN(n2944) );
  NAND2X0 U2726 ( .IN1(n2946), .IN2(\i_m4stg_frac/n215 ), .QN(n2943) );
  MUX21X1 U2727 ( .IN1(n2947), .IN2(n2948), .S(n2935), .Q(n2941) );
  AO221X1 U2728 ( .IN1(n1814), .IN2(n1136), .IN3(n1810), .IN4(n930), .IN5(
        n2949), .Q(n2935) );
  NAND2X0 U2729 ( .IN1(n2950), .IN2(n2938), .QN(n2948) );
  NAND2X0 U2730 ( .IN1(n2951), .IN2(n2934), .QN(n2947) );
  OR2X1 U2731 ( .IN1(n2950), .IN2(n2946), .Q(\i_m4stg_frac/booth/out_dff8/N5 )
         );
  OAI22X1 U2732 ( .IN1(n2952), .IN2(n2921), .IN3(n2953), .IN4(n2924), .QN(
        \i_m4stg_frac/booth/out_dff8/N4 ) );
  OA21X1 U2733 ( .IN1(n2954), .IN2(n2955), .IN3(n2956), .Q(n2953) );
  MUX21X1 U2734 ( .IN1(n2957), .IN2(n2934), .S(n2958), .Q(n2956) );
  OA21X1 U2735 ( .IN1(\i_m4stg_frac/n343 ), .IN2(\i_m4stg_frac/n211 ), .IN3(
        n2959), .Q(n2952) );
  INVX0 U2736 ( .INP(n2960), .ZN(n2959) );
  MUX21X1 U2737 ( .IN1(\i_m4stg_frac/n211 ), .IN2(\i_m4stg_frac/n343 ), .S(
        \i_m4stg_frac/n201 ), .Q(n2960) );
  NAND2X0 U2738 ( .IN1(n2961), .IN2(n2962), .QN(
        \i_m4stg_frac/booth/out_dff8/N3 ) );
  MUX21X1 U2739 ( .IN1(n2963), .IN2(n2964), .S(\i_m4stg_frac/n343 ), .Q(n2962)
         );
  NAND2X0 U2740 ( .IN1(n2946), .IN2(n944), .QN(n2964) );
  NOR2X0 U2741 ( .IN1(n1172), .IN2(n2921), .QN(n2946) );
  NAND2X0 U2742 ( .IN1(n2965), .IN2(n1172), .QN(n2963) );
  MUX21X1 U2743 ( .IN1(n2966), .IN2(n2967), .S(n2958), .Q(n2961) );
  AOI221X1 U2744 ( .IN1(n1814), .IN2(n1141), .IN3(n1810), .IN4(n892), .IN5(
        n2949), .QN(n2958) );
  NAND2X0 U2745 ( .IN1(n2954), .IN2(n2950), .QN(n2967) );
  NOR2X0 U2746 ( .IN1(n2924), .IN2(n2934), .QN(n2950) );
  NAND2X0 U2747 ( .IN1(n2968), .IN2(n2934), .QN(n2966) );
  INVX0 U2748 ( .INP(n2955), .ZN(n2934) );
  AO221X1 U2749 ( .IN1(n1814), .IN2(n930), .IN3(n1810), .IN4(n1141), .IN5(
        n2949), .Q(n2955) );
  OR2X1 U2750 ( .IN1(n2968), .IN2(n2965), .Q(\i_m4stg_frac/booth/out_dff7/N5 )
         );
  OAI22X1 U2751 ( .IN1(n2969), .IN2(n2921), .IN3(n2970), .IN4(n2924), .QN(
        \i_m4stg_frac/booth/out_dff7/N4 ) );
  OA21X1 U2752 ( .IN1(n2971), .IN2(n2957), .IN3(n2972), .Q(n2970) );
  MUX21X1 U2753 ( .IN1(n2973), .IN2(n2954), .S(n2974), .Q(n2972) );
  OA21X1 U2754 ( .IN1(n944), .IN2(n1323), .IN3(n2975), .Q(n2969) );
  MUX21X1 U2755 ( .IN1(\i_m4stg_frac/n341 ), .IN2(\i_m4stg_frac/n211 ), .S(
        \i_m4stg_frac/n205 ), .Q(n2975) );
  NAND2X0 U2756 ( .IN1(n2976), .IN2(n2977), .QN(
        \i_m4stg_frac/booth/out_dff7/N3 ) );
  MUX21X1 U2757 ( .IN1(n2978), .IN2(n2979), .S(\i_m4stg_frac/n341 ), .Q(n2977)
         );
  NAND2X0 U2758 ( .IN1(n2965), .IN2(n1173), .QN(n2979) );
  NOR2X0 U2759 ( .IN1(n944), .IN2(n2921), .QN(n2965) );
  NAND2X0 U2760 ( .IN1(n2980), .IN2(n944), .QN(n2978) );
  MUX21X1 U2761 ( .IN1(n2981), .IN2(n2982), .S(n2974), .Q(n2976) );
  AOI221X1 U2762 ( .IN1(n1814), .IN2(n1054), .IN3(n1810), .IN4(n927), .IN5(
        n2949), .QN(n2974) );
  NAND2X0 U2763 ( .IN1(n2971), .IN2(n2968), .QN(n2982) );
  NOR2X0 U2764 ( .IN1(n2924), .IN2(n2954), .QN(n2968) );
  NAND2X0 U2765 ( .IN1(n2983), .IN2(n2954), .QN(n2981) );
  INVX0 U2766 ( .INP(n2957), .ZN(n2954) );
  AO221X1 U2767 ( .IN1(n1814), .IN2(n892), .IN3(n1810), .IN4(n1054), .IN5(
        n2949), .Q(n2957) );
  OR2X1 U2768 ( .IN1(n2983), .IN2(n2980), .Q(\i_m4stg_frac/booth/out_dff6/N5 )
         );
  OAI22X1 U2769 ( .IN1(n2984), .IN2(n2921), .IN3(n2985), .IN4(n2924), .QN(
        \i_m4stg_frac/booth/out_dff6/N4 ) );
  OA21X1 U2770 ( .IN1(n2986), .IN2(n2973), .IN3(n2987), .Q(n2985) );
  MUX21X1 U2771 ( .IN1(n2988), .IN2(n2971), .S(n2989), .Q(n2987) );
  OA21X1 U2772 ( .IN1(\i_m4stg_frac/n339 ), .IN2(\i_m4stg_frac/n209 ), .IN3(
        n2990), .Q(n2984) );
  INVX0 U2773 ( .INP(n2991), .ZN(n2990) );
  MUX21X1 U2774 ( .IN1(\i_m4stg_frac/n209 ), .IN2(\i_m4stg_frac/n339 ), .S(
        \i_m4stg_frac/n205 ), .Q(n2991) );
  NAND2X0 U2775 ( .IN1(n2992), .IN2(n2993), .QN(
        \i_m4stg_frac/booth/out_dff6/N3 ) );
  MUX21X1 U2776 ( .IN1(n2994), .IN2(n2995), .S(\i_m4stg_frac/n339 ), .Q(n2993)
         );
  NAND2X0 U2777 ( .IN1(n2980), .IN2(n945), .QN(n2995) );
  NOR2X0 U2778 ( .IN1(n1173), .IN2(n2921), .QN(n2980) );
  NAND2X0 U2779 ( .IN1(n2996), .IN2(n1173), .QN(n2994) );
  MUX21X1 U2780 ( .IN1(n2997), .IN2(n2998), .S(n2989), .Q(n2992) );
  AOI221X1 U2781 ( .IN1(n1814), .IN2(n1113), .IN3(n1810), .IN4(n925), .IN5(
        n2949), .QN(n2989) );
  NAND2X0 U2782 ( .IN1(n2986), .IN2(n2983), .QN(n2998) );
  NOR2X0 U2783 ( .IN1(n2924), .IN2(n2971), .QN(n2983) );
  NAND2X0 U2784 ( .IN1(n2999), .IN2(n2971), .QN(n2997) );
  INVX0 U2785 ( .INP(n2973), .ZN(n2971) );
  AO221X1 U2786 ( .IN1(n1814), .IN2(n927), .IN3(n1810), .IN4(n1113), .IN5(
        n2949), .Q(n2973) );
  OR2X1 U2787 ( .IN1(n2999), .IN2(n2996), .Q(\i_m4stg_frac/booth/out_dff5/N5 )
         );
  OAI22X1 U2788 ( .IN1(n3000), .IN2(n2921), .IN3(n3001), .IN4(n2924), .QN(
        \i_m4stg_frac/booth/out_dff5/N4 ) );
  OA21X1 U2789 ( .IN1(n3002), .IN2(n2988), .IN3(n3003), .Q(n3001) );
  MUX21X1 U2790 ( .IN1(n3004), .IN2(n2986), .S(n3005), .Q(n3003) );
  OA21X1 U2791 ( .IN1(n945), .IN2(n1324), .IN3(n3006), .Q(n3000) );
  MUX21X1 U2792 ( .IN1(\i_m4stg_frac/n337 ), .IN2(\i_m4stg_frac/n209 ), .S(
        \i_m4stg_frac/n203 ), .Q(n3006) );
  NAND2X0 U2793 ( .IN1(n3007), .IN2(n3008), .QN(
        \i_m4stg_frac/booth/out_dff5/N3 ) );
  MUX21X1 U2794 ( .IN1(n3009), .IN2(n3010), .S(\i_m4stg_frac/n337 ), .Q(n3008)
         );
  NAND2X0 U2795 ( .IN1(n2996), .IN2(n946), .QN(n3010) );
  NOR2X0 U2796 ( .IN1(n945), .IN2(n2921), .QN(n2996) );
  NAND2X0 U2797 ( .IN1(n3011), .IN2(n945), .QN(n3009) );
  MUX21X1 U2798 ( .IN1(n3012), .IN2(n3013), .S(n3005), .Q(n3007) );
  AOI221X1 U2799 ( .IN1(n1814), .IN2(n881), .IN3(n1810), .IN4(n1137), .IN5(
        n2949), .QN(n3005) );
  NAND2X0 U2800 ( .IN1(n3002), .IN2(n2999), .QN(n3013) );
  NOR2X0 U2801 ( .IN1(n2924), .IN2(n2986), .QN(n2999) );
  NAND2X0 U2802 ( .IN1(n3014), .IN2(n2986), .QN(n3012) );
  INVX0 U2803 ( .INP(n2988), .ZN(n2986) );
  AO221X1 U2804 ( .IN1(n1814), .IN2(n925), .IN3(n1810), .IN4(n881), .IN5(n2949), .Q(n2988) );
  OR2X1 U2805 ( .IN1(n3014), .IN2(n3011), .Q(\i_m4stg_frac/booth/out_dff4/N5 )
         );
  OAI22X1 U2806 ( .IN1(n3015), .IN2(n2921), .IN3(n3016), .IN4(n2924), .QN(
        \i_m4stg_frac/booth/out_dff4/N4 ) );
  OA21X1 U2807 ( .IN1(n3017), .IN2(n3004), .IN3(n3018), .Q(n3016) );
  MUX21X1 U2808 ( .IN1(n3019), .IN2(n3002), .S(n3020), .Q(n3018) );
  OA21X1 U2809 ( .IN1(n946), .IN2(n1325), .IN3(n3021), .Q(n3015) );
  MUX21X1 U2810 ( .IN1(\i_m4stg_frac/n336 ), .IN2(\i_m4stg_frac/n203 ), .S(
        \i_m4stg_frac/n199 ), .Q(n3021) );
  NAND2X0 U2811 ( .IN1(n3022), .IN2(n3023), .QN(
        \i_m4stg_frac/booth/out_dff4/N3 ) );
  MUX21X1 U2812 ( .IN1(n3024), .IN2(n3025), .S(\i_m4stg_frac/n336 ), .Q(n3023)
         );
  NAND2X0 U2813 ( .IN1(n3011), .IN2(n1174), .QN(n3025) );
  NOR2X0 U2814 ( .IN1(n946), .IN2(n2921), .QN(n3011) );
  NAND2X0 U2815 ( .IN1(n3026), .IN2(n946), .QN(n3024) );
  MUX21X1 U2816 ( .IN1(n3027), .IN2(n3028), .S(n3020), .Q(n3022) );
  AOI221X1 U2817 ( .IN1(n1814), .IN2(n898), .IN3(n1810), .IN4(n953), .IN5(
        n2949), .QN(n3020) );
  NAND2X0 U2818 ( .IN1(n3017), .IN2(n3014), .QN(n3028) );
  NOR2X0 U2819 ( .IN1(n2924), .IN2(n3002), .QN(n3014) );
  NAND2X0 U2820 ( .IN1(n3029), .IN2(n3002), .QN(n3027) );
  INVX0 U2821 ( .INP(n3004), .ZN(n3002) );
  AO221X1 U2822 ( .IN1(n1814), .IN2(n1137), .IN3(n1810), .IN4(n898), .IN5(
        n2949), .Q(n3004) );
  OR2X1 U2823 ( .IN1(n3029), .IN2(n3026), .Q(\i_m4stg_frac/booth/out_dff3/N5 )
         );
  OAI22X1 U2824 ( .IN1(n3030), .IN2(n2921), .IN3(n3031), .IN4(n2924), .QN(
        \i_m4stg_frac/booth/out_dff3/N4 ) );
  OA21X1 U2825 ( .IN1(n3032), .IN2(n3019), .IN3(n3033), .Q(n3031) );
  MUX21X1 U2826 ( .IN1(n3034), .IN2(n3017), .S(n3035), .Q(n3033) );
  OA21X1 U2827 ( .IN1(\i_m4stg_frac/n335 ), .IN2(\i_m4stg_frac/n213 ), .IN3(
        n3036), .Q(n3030) );
  INVX0 U2828 ( .INP(n3037), .ZN(n3036) );
  MUX21X1 U2829 ( .IN1(\i_m4stg_frac/n213 ), .IN2(\i_m4stg_frac/n335 ), .S(
        \i_m4stg_frac/n199 ), .Q(n3037) );
  NAND2X0 U2830 ( .IN1(n3038), .IN2(n3039), .QN(
        \i_m4stg_frac/booth/out_dff3/N3 ) );
  MUX21X1 U2831 ( .IN1(n3040), .IN2(n3041), .S(\i_m4stg_frac/n335 ), .Q(n3039)
         );
  NAND2X0 U2832 ( .IN1(n3026), .IN2(n1127), .QN(n3041) );
  NOR2X0 U2833 ( .IN1(n1174), .IN2(n2921), .QN(n3026) );
  NAND2X0 U2834 ( .IN1(n3042), .IN2(n1174), .QN(n3040) );
  MUX21X1 U2835 ( .IN1(n3043), .IN2(n3044), .S(n3035), .Q(n3038) );
  AOI221X1 U2836 ( .IN1(n1814), .IN2(n1149), .IN3(n1810), .IN4(n941), .IN5(
        n2949), .QN(n3035) );
  NAND2X0 U2837 ( .IN1(n3032), .IN2(n3029), .QN(n3044) );
  NOR2X0 U2838 ( .IN1(n2924), .IN2(n3017), .QN(n3029) );
  NAND2X0 U2839 ( .IN1(n3045), .IN2(n3017), .QN(n3043) );
  INVX0 U2840 ( .INP(n3019), .ZN(n3017) );
  AO221X1 U2841 ( .IN1(n1814), .IN2(n953), .IN3(n1810), .IN4(n1149), .IN5(
        n2949), .Q(n3019) );
  OR2X1 U2842 ( .IN1(n3045), .IN2(n3042), .Q(\i_m4stg_frac/booth/out_dff2/N5 )
         );
  AO221X1 U2843 ( .IN1(\i_m4stg_frac/n850 ), .IN2(n3046), .IN3(n3047), .IN4(
        n1127), .IN5(n3048), .Q(\i_m4stg_frac/booth/out_dff2/N4 ) );
  MUX21X1 U2844 ( .IN1(n3049), .IN2(n3042), .S(\i_m4stg_frac/n1277 ), .Q(n3048) );
  NOR2X0 U2845 ( .IN1(\i_m4stg_frac/n333 ), .IN2(n2921), .QN(n3049) );
  AO21X1 U2846 ( .IN1(n3032), .IN2(m2stg_frac2_array_in[3]), .IN3(n3050), .Q(
        n3046) );
  MUX21X1 U2847 ( .IN1(n3051), .IN2(n3034), .S(n3052), .Q(n3050) );
  NAND2X0 U2848 ( .IN1(n3053), .IN2(n3054), .QN(
        \i_m4stg_frac/booth/out_dff2/N3 ) );
  MUX21X1 U2849 ( .IN1(n3055), .IN2(n3056), .S(\i_m4stg_frac/n1277 ), .Q(n3054) );
  NAND2X0 U2850 ( .IN1(n3042), .IN2(n1352), .QN(n3056) );
  NOR2X0 U2851 ( .IN1(n1127), .IN2(n2921), .QN(n3042) );
  NAND2X0 U2852 ( .IN1(n3047), .IN2(n1127), .QN(n3055) );
  MUX21X1 U2853 ( .IN1(n3057), .IN2(n3058), .S(n3052), .Q(n3053) );
  AOI221X1 U2854 ( .IN1(n1814), .IN2(n1155), .IN3(n1810), .IN4(n896), .IN5(
        n2949), .QN(n3052) );
  NAND2X0 U2855 ( .IN1(n3045), .IN2(n3051), .QN(n3058) );
  NOR2X0 U2856 ( .IN1(n2924), .IN2(n3032), .QN(n3045) );
  NAND2X0 U2857 ( .IN1(n3059), .IN2(n3032), .QN(n3057) );
  INVX0 U2858 ( .INP(n3034), .ZN(n3032) );
  AO221X1 U2859 ( .IN1(n1814), .IN2(n941), .IN3(n1810), .IN4(n1155), .IN5(
        n2949), .Q(n3034) );
  AO21X1 U2860 ( .IN1(\i_m4stg_frac/booth/out_dff15/N5 ), .IN2(n3060), .IN3(
        n3061), .Q(\i_m4stg_frac/booth/out_dff15/N4 ) );
  MUX21X1 U2861 ( .IN1(n3062), .IN2(\i_m4stg_frac/booth/out_dff14/N5 ), .S(
        n3063), .Q(n3061) );
  NOR2X0 U2862 ( .IN1(m2stg_frac2_array_in[31]), .IN2(n2924), .QN(n3062) );
  INVX0 U2863 ( .INP(n3064), .ZN(n3060) );
  INVX0 U2864 ( .INP(n3065), .ZN(\i_m4stg_frac/booth/out_dff15/N5 ) );
  MUX21X1 U2865 ( .IN1(n3066), .IN2(n3067), .S(n3063), .Q(
        \i_m4stg_frac/booth/out_dff15/N3 ) );
  AOI221X1 U2866 ( .IN1(n1814), .IN2(n1160), .IN3(n1810), .IN4(n959), .IN5(
        n3068), .QN(n3063) );
  AO221X1 U2867 ( .IN1(n1809), .IN2(n887), .IN3(n1812), .IN4(n1045), .IN5(
        n1816), .Q(n3068) );
  NOR2X0 U2868 ( .IN1(n3064), .IN2(n3065), .QN(n3067) );
  NAND2X0 U2869 ( .IN1(\i_m4stg_frac/n850 ), .IN2(m2stg_frac2_array_in[31]), 
        .QN(n3065) );
  NOR2X0 U2870 ( .IN1(m2stg_frac2_array_in[31]), .IN2(n3069), .QN(n3066) );
  AO221X1 U2871 ( .IN1(n1814), .IN2(n958), .IN3(n1810), .IN4(n1160), .IN5(
        n3070), .Q(m2stg_frac2_array_in[31]) );
  AO221X1 U2872 ( .IN1(n1809), .IN2(n1045), .IN3(n1812), .IN4(n919), .IN5(
        n1816), .Q(n3070) );
  NOR3X0 U2873 ( .IN1(n1880), .IN2(\fpu_mul_ctl/n117 ), .IN3(n1058), .QN(n1809) );
  AO21X1 U2874 ( .IN1(n3071), .IN2(\i_m4stg_frac/booth/out_dff14/N5 ), .IN3(
        n3072), .Q(\i_m4stg_frac/booth/out_dff14/N4 ) );
  MUX21X1 U2875 ( .IN1(n3073), .IN2(\i_m4stg_frac/booth/out_dff13/N5 ), .S(
        n3074), .Q(n3072) );
  NOR2X0 U2876 ( .IN1(n2924), .IN2(n3064), .QN(n3073) );
  INVX0 U2877 ( .INP(n3069), .ZN(\i_m4stg_frac/booth/out_dff14/N5 ) );
  INVX0 U2878 ( .INP(n3075), .ZN(n3071) );
  MUX21X1 U2879 ( .IN1(n3076), .IN2(n3077), .S(n3074), .Q(
        \i_m4stg_frac/booth/out_dff14/N3 ) );
  AOI221X1 U2880 ( .IN1(\fpu_mul_frac_dp/n837 ), .IN2(n1814), .IN3(n1810), 
        .IN4(n1148), .IN5(n2949), .QN(n3074) );
  NOR2X0 U2881 ( .IN1(n3069), .IN2(n3075), .QN(n3077) );
  NAND2X0 U2882 ( .IN1(\i_m4stg_frac/n850 ), .IN2(n3064), .QN(n3069) );
  NOR2X0 U2883 ( .IN1(n3064), .IN2(n3078), .QN(n3076) );
  AO221X1 U2884 ( .IN1(n1814), .IN2(n959), .IN3(\fpu_mul_frac_dp/n837 ), .IN4(
        n1810), .IN5(n3079), .Q(n3064) );
  AO21X1 U2885 ( .IN1(n1812), .IN2(n887), .IN3(n1816), .Q(n3079) );
  INVX0 U2886 ( .INP(n1803), .ZN(n1812) );
  NAND3X0 U2887 ( .IN1(n910), .IN2(n1058), .IN3(n3080), .QN(n1803) );
  NAND3X0 U2888 ( .IN1(n3081), .IN2(n1818), .IN3(n1880), .QN(n3080) );
  INVX0 U2889 ( .INP(n1876), .ZN(n1880) );
  OR2X1 U2890 ( .IN1(n3082), .IN2(n1853), .Q(n3081) );
  AO21X1 U2891 ( .IN1(n3083), .IN2(\i_m4stg_frac/booth/out_dff13/N5 ), .IN3(
        n3084), .Q(\i_m4stg_frac/booth/out_dff13/N4 ) );
  MUX21X1 U2892 ( .IN1(n3085), .IN2(\i_m4stg_frac/booth/out_dff12/N5 ), .S(
        n3086), .Q(n3084) );
  NOR2X0 U2893 ( .IN1(n2924), .IN2(n3075), .QN(n3085) );
  INVX0 U2894 ( .INP(n3078), .ZN(\i_m4stg_frac/booth/out_dff13/N5 ) );
  INVX0 U2895 ( .INP(n3087), .ZN(n3083) );
  MUX21X1 U2896 ( .IN1(n3088), .IN2(n3089), .S(n3086), .Q(
        \i_m4stg_frac/booth/out_dff13/N3 ) );
  AOI221X1 U2897 ( .IN1(n1814), .IN2(n897), .IN3(n1810), .IN4(n957), .IN5(
        n2949), .QN(n3086) );
  NOR2X0 U2898 ( .IN1(n3078), .IN2(n3087), .QN(n3089) );
  NAND2X0 U2899 ( .IN1(\i_m4stg_frac/n850 ), .IN2(n3075), .QN(n3078) );
  NOR2X0 U2900 ( .IN1(n3075), .IN2(n3090), .QN(n3088) );
  AO221X1 U2901 ( .IN1(n1814), .IN2(n1148), .IN3(n1810), .IN4(n897), .IN5(
        n2949), .Q(n3075) );
  AO21X1 U2902 ( .IN1(n3091), .IN2(\i_m4stg_frac/booth/out_dff12/N5 ), .IN3(
        n3092), .Q(\i_m4stg_frac/booth/out_dff12/N4 ) );
  MUX21X1 U2903 ( .IN1(n3093), .IN2(\i_m4stg_frac/booth/out_dff11/N5 ), .S(
        n3094), .Q(n3092) );
  NOR2X0 U2904 ( .IN1(n2924), .IN2(n3087), .QN(n3093) );
  INVX0 U2905 ( .INP(n3090), .ZN(\i_m4stg_frac/booth/out_dff12/N5 ) );
  INVX0 U2906 ( .INP(n3095), .ZN(n3091) );
  MUX21X1 U2907 ( .IN1(n3096), .IN2(n3097), .S(n3094), .Q(
        \i_m4stg_frac/booth/out_dff12/N3 ) );
  AOI221X1 U2908 ( .IN1(n1814), .IN2(n1157), .IN3(n1810), .IN4(n955), .IN5(
        n2949), .QN(n3094) );
  NOR2X0 U2909 ( .IN1(n3090), .IN2(n3095), .QN(n3097) );
  NAND2X0 U2910 ( .IN1(\i_m4stg_frac/n850 ), .IN2(n3087), .QN(n3090) );
  NOR2X0 U2911 ( .IN1(n3087), .IN2(n3098), .QN(n3096) );
  AO221X1 U2912 ( .IN1(n1814), .IN2(n957), .IN3(n1810), .IN4(n1157), .IN5(
        n2949), .Q(n3087) );
  AO21X1 U2913 ( .IN1(n3099), .IN2(\i_m4stg_frac/booth/out_dff11/N5 ), .IN3(
        n3100), .Q(\i_m4stg_frac/booth/out_dff11/N4 ) );
  MUX21X1 U2914 ( .IN1(n3101), .IN2(\i_m4stg_frac/n1283 ), .S(n3102), .Q(n3100) );
  INVX0 U2915 ( .INP(n3103), .ZN(\i_m4stg_frac/n1283 ) );
  NOR2X0 U2916 ( .IN1(n2924), .IN2(n3095), .QN(n3101) );
  INVX0 U2917 ( .INP(n3098), .ZN(\i_m4stg_frac/booth/out_dff11/N5 ) );
  MUX21X1 U2918 ( .IN1(n3104), .IN2(n3105), .S(n3102), .Q(
        \i_m4stg_frac/booth/out_dff11/N3 ) );
  AOI221X1 U2919 ( .IN1(n1814), .IN2(n1146), .IN3(n1810), .IN4(n940), .IN5(
        n2949), .QN(n3102) );
  NOR2X0 U2920 ( .IN1(n3098), .IN2(n3106), .QN(n3105) );
  NAND2X0 U2921 ( .IN1(\i_m4stg_frac/n850 ), .IN2(n3095), .QN(n3098) );
  NOR2X0 U2922 ( .IN1(n3095), .IN2(n3103), .QN(n3104) );
  AO221X1 U2923 ( .IN1(n1814), .IN2(n955), .IN3(n1810), .IN4(n1146), .IN5(
        n2949), .Q(n3095) );
  NAND4X0 U2924 ( .IN1(n3107), .IN2(n3108), .IN3(n3109), .IN4(n2931), .QN(
        \i_m4stg_frac/booth/out_dff10/N4 ) );
  NAND2X0 U2925 ( .IN1(n3099), .IN2(n2951), .QN(n3109) );
  INVX0 U2926 ( .INP(n2930), .ZN(n2951) );
  INVX0 U2927 ( .INP(n3106), .ZN(n3099) );
  NAND2X0 U2928 ( .IN1(\i_m4stg_frac/n1285 ), .IN2(n1278), .QN(n3108) );
  MUX21X1 U2929 ( .IN1(n3110), .IN2(n3103), .S(n3111), .Q(n3107) );
  NAND2X0 U2930 ( .IN1(n2938), .IN2(\i_m4stg_frac/n850 ), .QN(n3110) );
  INVX0 U2931 ( .INP(n3112), .ZN(n2938) );
  AO21X1 U2932 ( .IN1(n2945), .IN2(n1278), .IN3(n3113), .Q(
        \i_m4stg_frac/booth/out_dff10/N3 ) );
  MUX21X1 U2933 ( .IN1(n3114), .IN2(n3115), .S(n3111), .Q(n3113) );
  AOI221X1 U2934 ( .IN1(n1814), .IN2(n1156), .IN3(n1810), .IN4(n932), .IN5(
        n2949), .QN(n3111) );
  NOR2X0 U2935 ( .IN1(n3112), .IN2(n3103), .QN(n3115) );
  NAND2X0 U2936 ( .IN1(\i_m4stg_frac/n850 ), .IN2(n3106), .QN(n3103) );
  NOR2X0 U2937 ( .IN1(n2930), .IN2(n3106), .QN(n3114) );
  AO221X1 U2938 ( .IN1(n1814), .IN2(n940), .IN3(n1810), .IN4(n1156), .IN5(
        n2949), .Q(n3106) );
  NAND2X0 U2939 ( .IN1(\i_m4stg_frac/n850 ), .IN2(n3112), .QN(n2930) );
  AO221X1 U2940 ( .IN1(n1814), .IN2(n932), .IN3(n1810), .IN4(n1136), .IN5(
        n2949), .Q(n3112) );
  INVX0 U2941 ( .INP(n2931), .ZN(n2945) );
  NAND2X0 U2942 ( .IN1(\i_m4stg_frac/n1285 ), .IN2(n1161), .QN(n2931) );
  NAND4X0 U2943 ( .IN1(n3116), .IN2(n3117), .IN3(n3118), .IN4(n3119), .QN(
        \i_m4stg_frac/booth/out_dff1/N4 ) );
  MUX21X1 U2944 ( .IN1(n3120), .IN2(n3121), .S(n3122), .Q(n3117) );
  NAND2X0 U2945 ( .IN1(\i_m4stg_frac/n850 ), .IN2(n3123), .QN(n3120) );
  MUX21X1 U2946 ( .IN1(n3124), .IN2(\i_m4stg_frac/n1684 ), .S(
        \i_m4stg_frac/n1281 ), .Q(n3116) );
  NAND2X0 U2947 ( .IN1(\i_m4stg_frac/n1285 ), .IN2(\i_m4stg_frac/n207 ), .QN(
        n3124) );
  NAND2X0 U2948 ( .IN1(n3125), .IN2(n3126), .QN(
        \i_m4stg_frac/booth/out_dff1/N3 ) );
  MUX21X1 U2949 ( .IN1(n3118), .IN2(n3127), .S(n3122), .Q(n3126) );
  AOI221X1 U2950 ( .IN1(n1814), .IN2(n1147), .IN3(n1810), .IN4(n939), .IN5(
        n2949), .QN(n3122) );
  NAND2X0 U2951 ( .IN1(n3059), .IN2(n3123), .QN(n3127) );
  INVX0 U2952 ( .INP(m2stg_frac2_array_in[1]), .ZN(n3123) );
  INVX0 U2953 ( .INP(n3121), .ZN(n3059) );
  NAND2X0 U2954 ( .IN1(\i_m4stg_frac/n850 ), .IN2(m2stg_frac2_array_in[3]), 
        .QN(n3121) );
  NAND2X0 U2955 ( .IN1(n3128), .IN2(n3051), .QN(n3118) );
  INVX0 U2956 ( .INP(m2stg_frac2_array_in[3]), .ZN(n3051) );
  AO221X1 U2957 ( .IN1(n1814), .IN2(n896), .IN3(n1810), .IN4(n1147), .IN5(
        n2949), .Q(m2stg_frac2_array_in[3]) );
  MUX21X1 U2958 ( .IN1(n3119), .IN2(n3129), .S(\i_m4stg_frac/n1281 ), .Q(n3125) );
  NAND2X0 U2959 ( .IN1(\i_m4stg_frac/n207 ), .IN2(n3047), .QN(n3129) );
  INVX0 U2960 ( .INP(\i_m4stg_frac/n1684 ), .ZN(n3047) );
  NAND2X0 U2961 ( .IN1(\i_m4stg_frac/n333 ), .IN2(\i_m4stg_frac/n1285 ), .QN(
        \i_m4stg_frac/n1684 ) );
  OR3X1 U2962 ( .IN1(\i_m4stg_frac/n207 ), .IN2(\i_m4stg_frac/n333 ), .IN3(
        n2921), .Q(n3119) );
  AO22X1 U2963 ( .IN1(n2923), .IN2(n3128), .IN3(n3130), .IN4(
        \i_m4stg_frac/n1285 ), .Q(\i_m4stg_frac/booth/out_dff0/N3 ) );
  INVX0 U2964 ( .INP(n2921), .ZN(\i_m4stg_frac/n1285 ) );
  NAND2X0 U2965 ( .IN1(n3131), .IN2(\i_m4stg_frac/n854 ), .QN(n2921) );
  MUX21X1 U2966 ( .IN1(n3132), .IN2(n3133), .S(\i_m4stg_frac/n345 ), .Q(n3130)
         );
  NOR2X0 U2967 ( .IN1(\i_m4stg_frac/n300 ), .IN2(\i_m4stg_frac/n207 ), .QN(
        n3133) );
  AND2X1 U2968 ( .IN1(\i_m4stg_frac/n300 ), .IN2(\i_m4stg_frac/n207 ), .Q(
        n3132) );
  INVX0 U2969 ( .INP(\i_m4stg_frac/n1692 ), .ZN(n3128) );
  NAND2X0 U2970 ( .IN1(\i_m4stg_frac/n850 ), .IN2(m2stg_frac2_array_in[1]), 
        .QN(\i_m4stg_frac/n1692 ) );
  AO221X1 U2971 ( .IN1(n1814), .IN2(n939), .IN3(n1810), .IN4(n1158), .IN5(
        n2949), .Q(m2stg_frac2_array_in[1]) );
  INVX0 U2972 ( .INP(n1807), .ZN(n1810) );
  NAND3X0 U2973 ( .IN1(n1882), .IN2(n886), .IN3(\fpu_mul_ctl/n264 ), .QN(n1807) );
  INVX0 U2974 ( .INP(n2924), .ZN(\i_m4stg_frac/n850 ) );
  NAND2X0 U2975 ( .IN1(\i_m4stg_frac/n854 ), .IN2(n2928), .QN(n2924) );
  INVX0 U2976 ( .INP(se_mul64), .ZN(\i_m4stg_frac/n854 ) );
  AOI21X1 U2977 ( .IN1(n1814), .IN2(n1158), .IN3(n2949), .QN(n2923) );
  AND2X1 U2978 ( .IN1(n1816), .IN2(n3134), .Q(n2949) );
  AOI21X1 U2979 ( .IN1(n3135), .IN2(n3136), .IN3(n1808), .QN(n1816) );
  AND3X1 U2980 ( .IN1(n3137), .IN2(n1845), .IN3(n3138), .Q(n1808) );
  NAND3X0 U2981 ( .IN1(n1817), .IN2(n3139), .IN3(n1818), .QN(n3138) );
  AO221X1 U2982 ( .IN1(n3140), .IN2(n3141), .IN3(\fpu_mul_ctl/n256 ), .IN4(
        n3142), .IN5(n3143), .Q(n1845) );
  OAI22X1 U2983 ( .IN1(n3144), .IN2(\fpu_mul_ctl/n259 ), .IN3(n1338), .IN4(
        n3145), .QN(n3142) );
  NAND2X0 U2984 ( .IN1(n885), .IN2(n3146), .QN(n3140) );
  OR3X1 U2985 ( .IN1(n1037), .IN2(n3147), .IN3(n3143), .Q(n3137) );
  NAND3X0 U2986 ( .IN1(n3146), .IN2(n885), .IN3(n3148), .QN(n3136) );
  NAND2X0 U2987 ( .IN1(n3149), .IN2(n3150), .QN(n3135) );
  INVX0 U2988 ( .INP(n1804), .ZN(n1814) );
  NAND3X0 U2989 ( .IN1(n886), .IN2(n1058), .IN3(n3151), .QN(n1804) );
  NAND3X0 U2990 ( .IN1(n3152), .IN2(n1817), .IN3(n1886), .QN(n3151) );
  INVX0 U2991 ( .INP(n1882), .ZN(n1886) );
  OR2X1 U2992 ( .IN1(n3153), .IN2(n1854), .Q(n3152) );
  XNOR3X1 U2993 ( .IN1(\i_m4stg_frac/n158 ), .IN2(\i_m4stg_frac/n323 ), .IN3(
        n3154), .Q(\i_m4stg_frac/addout[9] ) );
  XNOR3X1 U2994 ( .IN1(\i_m4stg_frac/n159 ), .IN2(\i_m4stg_frac/n324 ), .IN3(
        n3155), .Q(\i_m4stg_frac/addout[8] ) );
  XNOR3X1 U2995 ( .IN1(\i_m4stg_frac/n160 ), .IN2(\i_m4stg_frac/n325 ), .IN3(
        n3156), .Q(\i_m4stg_frac/addout[7] ) );
  XOR3X1 U2996 ( .IN1(\i_m4stg_frac/n52 ), .IN2(\i_m4stg_frac/n217 ), .IN3(
        n3157), .Q(\i_m4stg_frac/addout[73] ) );
  AOI22X1 U2997 ( .IN1(n3158), .IN2(\i_m4stg_frac/n54 ), .IN3(n3159), .IN4(
        \i_m4stg_frac/n219 ), .QN(n3157) );
  OR2X1 U2998 ( .IN1(\i_m4stg_frac/n219 ), .IN2(n3159), .Q(n3158) );
  XNOR3X1 U2999 ( .IN1(\i_m4stg_frac/n219 ), .IN2(\i_m4stg_frac/n54 ), .IN3(
        n3159), .Q(\i_m4stg_frac/addout[72] ) );
  AO22X1 U3000 ( .IN1(\i_m4stg_frac/n221 ), .IN2(n3160), .IN3(
        \i_m4stg_frac/n56 ), .IN4(n3161), .Q(n3159) );
  OR2X1 U3001 ( .IN1(n3160), .IN2(\i_m4stg_frac/n221 ), .Q(n3161) );
  XNOR3X1 U3002 ( .IN1(\i_m4stg_frac/n56 ), .IN2(\i_m4stg_frac/n221 ), .IN3(
        n3160), .Q(\i_m4stg_frac/addout[71] ) );
  AO22X1 U3003 ( .IN1(\i_m4stg_frac/n223 ), .IN2(n3162), .IN3(
        \i_m4stg_frac/n58 ), .IN4(n3163), .Q(n3160) );
  OR2X1 U3004 ( .IN1(n3162), .IN2(\i_m4stg_frac/n223 ), .Q(n3163) );
  XNOR3X1 U3005 ( .IN1(\i_m4stg_frac/n223 ), .IN2(\i_m4stg_frac/n58 ), .IN3(
        n3162), .Q(\i_m4stg_frac/addout[70] ) );
  AO22X1 U3006 ( .IN1(\i_m4stg_frac/n225 ), .IN2(n3164), .IN3(
        \i_m4stg_frac/n60 ), .IN4(n3165), .Q(n3162) );
  OR2X1 U3007 ( .IN1(n3164), .IN2(\i_m4stg_frac/n225 ), .Q(n3165) );
  XNOR3X1 U3008 ( .IN1(\i_m4stg_frac/n161 ), .IN2(\i_m4stg_frac/n326 ), .IN3(
        n3166), .Q(\i_m4stg_frac/addout[6] ) );
  XNOR3X1 U3009 ( .IN1(\i_m4stg_frac/n60 ), .IN2(\i_m4stg_frac/n225 ), .IN3(
        n3164), .Q(\i_m4stg_frac/addout[69] ) );
  AO22X1 U3010 ( .IN1(\i_m4stg_frac/n227 ), .IN2(n3167), .IN3(
        \i_m4stg_frac/n62 ), .IN4(n3168), .Q(n3164) );
  OR2X1 U3011 ( .IN1(n3167), .IN2(\i_m4stg_frac/n227 ), .Q(n3168) );
  XNOR3X1 U3012 ( .IN1(\i_m4stg_frac/n227 ), .IN2(\i_m4stg_frac/n62 ), .IN3(
        n3167), .Q(\i_m4stg_frac/addout[68] ) );
  AO22X1 U3013 ( .IN1(\i_m4stg_frac/n229 ), .IN2(n3169), .IN3(
        \i_m4stg_frac/n64 ), .IN4(n3170), .Q(n3167) );
  OR2X1 U3014 ( .IN1(n3169), .IN2(\i_m4stg_frac/n229 ), .Q(n3170) );
  XNOR3X1 U3015 ( .IN1(\i_m4stg_frac/n64 ), .IN2(\i_m4stg_frac/n229 ), .IN3(
        n3169), .Q(\i_m4stg_frac/addout[67] ) );
  AO22X1 U3016 ( .IN1(\i_m4stg_frac/n231 ), .IN2(n3171), .IN3(
        \i_m4stg_frac/n66 ), .IN4(n3172), .Q(n3169) );
  OR2X1 U3017 ( .IN1(n3171), .IN2(\i_m4stg_frac/n231 ), .Q(n3172) );
  XNOR3X1 U3018 ( .IN1(\i_m4stg_frac/n231 ), .IN2(\i_m4stg_frac/n66 ), .IN3(
        n3171), .Q(\i_m4stg_frac/addout[66] ) );
  AO22X1 U3019 ( .IN1(\i_m4stg_frac/n233 ), .IN2(n3173), .IN3(
        \i_m4stg_frac/n68 ), .IN4(n3174), .Q(n3171) );
  OR2X1 U3020 ( .IN1(n3173), .IN2(\i_m4stg_frac/n233 ), .Q(n3174) );
  XNOR3X1 U3021 ( .IN1(\i_m4stg_frac/n68 ), .IN2(\i_m4stg_frac/n233 ), .IN3(
        n3173), .Q(\i_m4stg_frac/addout[65] ) );
  AO22X1 U3022 ( .IN1(\i_m4stg_frac/n235 ), .IN2(n3175), .IN3(
        \i_m4stg_frac/n70 ), .IN4(n3176), .Q(n3173) );
  OR2X1 U3023 ( .IN1(n3175), .IN2(\i_m4stg_frac/n235 ), .Q(n3176) );
  XNOR3X1 U3024 ( .IN1(\i_m4stg_frac/n235 ), .IN2(\i_m4stg_frac/n70 ), .IN3(
        n3175), .Q(\i_m4stg_frac/addout[64] ) );
  AO22X1 U3025 ( .IN1(\i_m4stg_frac/n237 ), .IN2(n3177), .IN3(
        \i_m4stg_frac/n72 ), .IN4(n3178), .Q(n3175) );
  OR2X1 U3026 ( .IN1(n3177), .IN2(\i_m4stg_frac/n237 ), .Q(n3178) );
  XNOR3X1 U3027 ( .IN1(\i_m4stg_frac/n72 ), .IN2(\i_m4stg_frac/n237 ), .IN3(
        n3177), .Q(\i_m4stg_frac/addout[63] ) );
  AO22X1 U3028 ( .IN1(\i_m4stg_frac/n239 ), .IN2(n3179), .IN3(
        \i_m4stg_frac/n74 ), .IN4(n3180), .Q(n3177) );
  OR2X1 U3029 ( .IN1(n3179), .IN2(\i_m4stg_frac/n239 ), .Q(n3180) );
  XNOR3X1 U3030 ( .IN1(\i_m4stg_frac/n239 ), .IN2(\i_m4stg_frac/n74 ), .IN3(
        n3179), .Q(\i_m4stg_frac/addout[62] ) );
  AO22X1 U3031 ( .IN1(\i_m4stg_frac/n241 ), .IN2(n3181), .IN3(
        \i_m4stg_frac/n76 ), .IN4(n3182), .Q(n3179) );
  OR2X1 U3032 ( .IN1(n3181), .IN2(\i_m4stg_frac/n241 ), .Q(n3182) );
  XNOR3X1 U3033 ( .IN1(\i_m4stg_frac/n76 ), .IN2(\i_m4stg_frac/n241 ), .IN3(
        n3181), .Q(\i_m4stg_frac/addout[61] ) );
  AO22X1 U3034 ( .IN1(\i_m4stg_frac/n243 ), .IN2(n3183), .IN3(
        \i_m4stg_frac/n78 ), .IN4(n3184), .Q(n3181) );
  OR2X1 U3035 ( .IN1(n3183), .IN2(\i_m4stg_frac/n243 ), .Q(n3184) );
  XNOR3X1 U3036 ( .IN1(\i_m4stg_frac/n243 ), .IN2(\i_m4stg_frac/n78 ), .IN3(
        n3183), .Q(\i_m4stg_frac/addout[60] ) );
  AO22X1 U3037 ( .IN1(\i_m4stg_frac/n245 ), .IN2(n3185), .IN3(
        \i_m4stg_frac/n80 ), .IN4(n3186), .Q(n3183) );
  OR2X1 U3038 ( .IN1(n3185), .IN2(\i_m4stg_frac/n245 ), .Q(n3186) );
  XNOR3X1 U3039 ( .IN1(\i_m4stg_frac/n162 ), .IN2(\i_m4stg_frac/n327 ), .IN3(
        n3187), .Q(\i_m4stg_frac/addout[5] ) );
  XNOR3X1 U3040 ( .IN1(\i_m4stg_frac/n80 ), .IN2(\i_m4stg_frac/n245 ), .IN3(
        n3185), .Q(\i_m4stg_frac/addout[59] ) );
  AO22X1 U3041 ( .IN1(\i_m4stg_frac/n247 ), .IN2(n3188), .IN3(
        \i_m4stg_frac/n82 ), .IN4(n3189), .Q(n3185) );
  OR2X1 U3042 ( .IN1(n3188), .IN2(\i_m4stg_frac/n247 ), .Q(n3189) );
  XNOR3X1 U3043 ( .IN1(\i_m4stg_frac/n247 ), .IN2(\i_m4stg_frac/n82 ), .IN3(
        n3188), .Q(\i_m4stg_frac/addout[58] ) );
  AO22X1 U3044 ( .IN1(\i_m4stg_frac/n249 ), .IN2(n3190), .IN3(
        \i_m4stg_frac/n84 ), .IN4(n3191), .Q(n3188) );
  OR2X1 U3045 ( .IN1(n3190), .IN2(\i_m4stg_frac/n249 ), .Q(n3191) );
  XNOR3X1 U3046 ( .IN1(\i_m4stg_frac/n84 ), .IN2(\i_m4stg_frac/n249 ), .IN3(
        n3190), .Q(\i_m4stg_frac/addout[57] ) );
  AO22X1 U3047 ( .IN1(\i_m4stg_frac/n251 ), .IN2(n3192), .IN3(
        \i_m4stg_frac/n86 ), .IN4(n3193), .Q(n3190) );
  OR2X1 U3048 ( .IN1(n3192), .IN2(\i_m4stg_frac/n251 ), .Q(n3193) );
  XNOR3X1 U3049 ( .IN1(\i_m4stg_frac/n251 ), .IN2(\i_m4stg_frac/n86 ), .IN3(
        n3192), .Q(\i_m4stg_frac/addout[56] ) );
  AO22X1 U3050 ( .IN1(\i_m4stg_frac/n253 ), .IN2(n3194), .IN3(
        \i_m4stg_frac/n88 ), .IN4(n3195), .Q(n3192) );
  OR2X1 U3051 ( .IN1(n3194), .IN2(\i_m4stg_frac/n253 ), .Q(n3195) );
  XNOR3X1 U3052 ( .IN1(\i_m4stg_frac/n88 ), .IN2(\i_m4stg_frac/n253 ), .IN3(
        n3194), .Q(\i_m4stg_frac/addout[55] ) );
  AO22X1 U3053 ( .IN1(\i_m4stg_frac/n255 ), .IN2(n3196), .IN3(
        \i_m4stg_frac/n90 ), .IN4(n3197), .Q(n3194) );
  OR2X1 U3054 ( .IN1(n3196), .IN2(\i_m4stg_frac/n255 ), .Q(n3197) );
  XNOR3X1 U3055 ( .IN1(\i_m4stg_frac/n255 ), .IN2(\i_m4stg_frac/n90 ), .IN3(
        n3196), .Q(\i_m4stg_frac/addout[54] ) );
  AO22X1 U3056 ( .IN1(\i_m4stg_frac/n257 ), .IN2(n3198), .IN3(
        \i_m4stg_frac/n92 ), .IN4(n3199), .Q(n3196) );
  OR2X1 U3057 ( .IN1(n3198), .IN2(\i_m4stg_frac/n257 ), .Q(n3199) );
  XNOR3X1 U3058 ( .IN1(\i_m4stg_frac/n92 ), .IN2(\i_m4stg_frac/n257 ), .IN3(
        n3198), .Q(\i_m4stg_frac/addout[53] ) );
  AO22X1 U3059 ( .IN1(\i_m4stg_frac/n259 ), .IN2(n3200), .IN3(
        \i_m4stg_frac/n94 ), .IN4(n3201), .Q(n3198) );
  OR2X1 U3060 ( .IN1(n3200), .IN2(\i_m4stg_frac/n259 ), .Q(n3201) );
  XNOR3X1 U3061 ( .IN1(\i_m4stg_frac/n259 ), .IN2(\i_m4stg_frac/n94 ), .IN3(
        n3200), .Q(\i_m4stg_frac/addout[52] ) );
  AO22X1 U3062 ( .IN1(\i_m4stg_frac/n261 ), .IN2(n3202), .IN3(
        \i_m4stg_frac/n96 ), .IN4(n3203), .Q(n3200) );
  OR2X1 U3063 ( .IN1(n3202), .IN2(\i_m4stg_frac/n261 ), .Q(n3203) );
  XNOR3X1 U3064 ( .IN1(\i_m4stg_frac/n96 ), .IN2(\i_m4stg_frac/n261 ), .IN3(
        n3202), .Q(\i_m4stg_frac/addout[51] ) );
  AO22X1 U3065 ( .IN1(\i_m4stg_frac/n263 ), .IN2(n3204), .IN3(
        \i_m4stg_frac/n98 ), .IN4(n3205), .Q(n3202) );
  OR2X1 U3066 ( .IN1(n3204), .IN2(\i_m4stg_frac/n263 ), .Q(n3205) );
  XNOR3X1 U3067 ( .IN1(\i_m4stg_frac/n263 ), .IN2(\i_m4stg_frac/n98 ), .IN3(
        n3204), .Q(\i_m4stg_frac/addout[50] ) );
  AO22X1 U3068 ( .IN1(\i_m4stg_frac/n100 ), .IN2(n3206), .IN3(
        \i_m4stg_frac/n265 ), .IN4(n3207), .Q(n3204) );
  OR2X1 U3069 ( .IN1(n3206), .IN2(\i_m4stg_frac/n100 ), .Q(n3207) );
  XNOR3X1 U3070 ( .IN1(\i_m4stg_frac/n163 ), .IN2(\i_m4stg_frac/n328 ), .IN3(
        n3208), .Q(\i_m4stg_frac/addout[4] ) );
  XNOR3X1 U3071 ( .IN1(\i_m4stg_frac/n265 ), .IN2(\i_m4stg_frac/n100 ), .IN3(
        n3206), .Q(\i_m4stg_frac/addout[49] ) );
  AO22X1 U3072 ( .IN1(\i_m4stg_frac/n102 ), .IN2(n3209), .IN3(
        \i_m4stg_frac/n267 ), .IN4(n3210), .Q(n3206) );
  OR2X1 U3073 ( .IN1(n3209), .IN2(\i_m4stg_frac/n102 ), .Q(n3210) );
  XNOR3X1 U3074 ( .IN1(\i_m4stg_frac/n102 ), .IN2(\i_m4stg_frac/n267 ), .IN3(
        n3209), .Q(\i_m4stg_frac/addout[48] ) );
  AO22X1 U3075 ( .IN1(\i_m4stg_frac/n104 ), .IN2(n3211), .IN3(
        \i_m4stg_frac/n269 ), .IN4(n3212), .Q(n3209) );
  OR2X1 U3076 ( .IN1(n3211), .IN2(\i_m4stg_frac/n104 ), .Q(n3212) );
  XNOR3X1 U3077 ( .IN1(\i_m4stg_frac/n269 ), .IN2(\i_m4stg_frac/n104 ), .IN3(
        n3211), .Q(\i_m4stg_frac/addout[47] ) );
  AO22X1 U3078 ( .IN1(\i_m4stg_frac/n106 ), .IN2(n3213), .IN3(
        \i_m4stg_frac/n271 ), .IN4(n3214), .Q(n3211) );
  OR2X1 U3079 ( .IN1(n3213), .IN2(\i_m4stg_frac/n106 ), .Q(n3214) );
  XNOR3X1 U3080 ( .IN1(\i_m4stg_frac/n106 ), .IN2(\i_m4stg_frac/n271 ), .IN3(
        n3213), .Q(\i_m4stg_frac/addout[46] ) );
  AO22X1 U3081 ( .IN1(\i_m4stg_frac/n108 ), .IN2(n3215), .IN3(
        \i_m4stg_frac/n273 ), .IN4(n3216), .Q(n3213) );
  OR2X1 U3082 ( .IN1(n3215), .IN2(\i_m4stg_frac/n108 ), .Q(n3216) );
  XNOR3X1 U3083 ( .IN1(\i_m4stg_frac/n273 ), .IN2(\i_m4stg_frac/n108 ), .IN3(
        n3215), .Q(\i_m4stg_frac/addout[45] ) );
  AO22X1 U3084 ( .IN1(\i_m4stg_frac/n110 ), .IN2(n3217), .IN3(
        \i_m4stg_frac/n275 ), .IN4(n3218), .Q(n3215) );
  OR2X1 U3085 ( .IN1(n3217), .IN2(\i_m4stg_frac/n110 ), .Q(n3218) );
  XNOR3X1 U3086 ( .IN1(\i_m4stg_frac/n110 ), .IN2(\i_m4stg_frac/n275 ), .IN3(
        n3217), .Q(\i_m4stg_frac/addout[44] ) );
  AO22X1 U3087 ( .IN1(\i_m4stg_frac/n112 ), .IN2(n3219), .IN3(
        \i_m4stg_frac/n277 ), .IN4(n3220), .Q(n3217) );
  OR2X1 U3088 ( .IN1(n3219), .IN2(\i_m4stg_frac/n112 ), .Q(n3220) );
  XNOR3X1 U3089 ( .IN1(\i_m4stg_frac/n277 ), .IN2(\i_m4stg_frac/n112 ), .IN3(
        n3219), .Q(\i_m4stg_frac/addout[43] ) );
  AO22X1 U3090 ( .IN1(\i_m4stg_frac/n114 ), .IN2(n3221), .IN3(
        \i_m4stg_frac/n279 ), .IN4(n3222), .Q(n3219) );
  OR2X1 U3091 ( .IN1(n3221), .IN2(\i_m4stg_frac/n114 ), .Q(n3222) );
  XNOR3X1 U3092 ( .IN1(\i_m4stg_frac/n114 ), .IN2(\i_m4stg_frac/n279 ), .IN3(
        n3221), .Q(\i_m4stg_frac/addout[42] ) );
  AO22X1 U3093 ( .IN1(\i_m4stg_frac/n116 ), .IN2(n3223), .IN3(
        \i_m4stg_frac/n281 ), .IN4(n3224), .Q(n3221) );
  OR2X1 U3094 ( .IN1(n3223), .IN2(\i_m4stg_frac/n116 ), .Q(n3224) );
  XNOR3X1 U3095 ( .IN1(\i_m4stg_frac/n281 ), .IN2(\i_m4stg_frac/n116 ), .IN3(
        n3223), .Q(\i_m4stg_frac/addout[41] ) );
  AO22X1 U3096 ( .IN1(\i_m4stg_frac/n118 ), .IN2(n3225), .IN3(
        \i_m4stg_frac/n283 ), .IN4(n3226), .Q(n3223) );
  OR2X1 U3097 ( .IN1(n3225), .IN2(\i_m4stg_frac/n118 ), .Q(n3226) );
  XNOR3X1 U3098 ( .IN1(\i_m4stg_frac/n118 ), .IN2(\i_m4stg_frac/n283 ), .IN3(
        n3225), .Q(\i_m4stg_frac/addout[40] ) );
  AO22X1 U3099 ( .IN1(\i_m4stg_frac/n120 ), .IN2(n3227), .IN3(
        \i_m4stg_frac/n285 ), .IN4(n3228), .Q(n3225) );
  OR2X1 U3100 ( .IN1(n3227), .IN2(\i_m4stg_frac/n120 ), .Q(n3228) );
  XNOR3X1 U3101 ( .IN1(\i_m4stg_frac/n164 ), .IN2(\i_m4stg_frac/n329 ), .IN3(
        n3229), .Q(\i_m4stg_frac/addout[3] ) );
  XNOR3X1 U3102 ( .IN1(\i_m4stg_frac/n285 ), .IN2(\i_m4stg_frac/n120 ), .IN3(
        n3227), .Q(\i_m4stg_frac/addout[39] ) );
  AO22X1 U3103 ( .IN1(\i_m4stg_frac/n122 ), .IN2(n3230), .IN3(
        \i_m4stg_frac/n287 ), .IN4(n3231), .Q(n3227) );
  OR2X1 U3104 ( .IN1(n3230), .IN2(\i_m4stg_frac/n122 ), .Q(n3231) );
  XNOR3X1 U3105 ( .IN1(\i_m4stg_frac/n122 ), .IN2(\i_m4stg_frac/n287 ), .IN3(
        n3230), .Q(\i_m4stg_frac/addout[38] ) );
  AO22X1 U3106 ( .IN1(\i_m4stg_frac/n124 ), .IN2(n3232), .IN3(
        \i_m4stg_frac/n289 ), .IN4(n3233), .Q(n3230) );
  OR2X1 U3107 ( .IN1(n3232), .IN2(\i_m4stg_frac/n124 ), .Q(n3233) );
  XNOR3X1 U3108 ( .IN1(\i_m4stg_frac/n289 ), .IN2(\i_m4stg_frac/n124 ), .IN3(
        n3232), .Q(\i_m4stg_frac/addout[37] ) );
  AO22X1 U3109 ( .IN1(\i_m4stg_frac/n126 ), .IN2(n3234), .IN3(
        \i_m4stg_frac/n291 ), .IN4(n3235), .Q(n3232) );
  OR2X1 U3110 ( .IN1(n3234), .IN2(\i_m4stg_frac/n126 ), .Q(n3235) );
  XNOR3X1 U3111 ( .IN1(\i_m4stg_frac/n126 ), .IN2(\i_m4stg_frac/n291 ), .IN3(
        n3234), .Q(\i_m4stg_frac/addout[36] ) );
  AO22X1 U3112 ( .IN1(\i_m4stg_frac/n128 ), .IN2(n3236), .IN3(
        \i_m4stg_frac/n293 ), .IN4(n3237), .Q(n3234) );
  OR2X1 U3113 ( .IN1(n3236), .IN2(\i_m4stg_frac/n128 ), .Q(n3237) );
  XNOR3X1 U3114 ( .IN1(\i_m4stg_frac/n293 ), .IN2(\i_m4stg_frac/n128 ), .IN3(
        n3236), .Q(\i_m4stg_frac/addout[35] ) );
  AO22X1 U3115 ( .IN1(\i_m4stg_frac/n130 ), .IN2(n3238), .IN3(
        \i_m4stg_frac/n295 ), .IN4(n3239), .Q(n3236) );
  OR2X1 U3116 ( .IN1(n3238), .IN2(\i_m4stg_frac/n130 ), .Q(n3239) );
  XNOR3X1 U3117 ( .IN1(\i_m4stg_frac/n130 ), .IN2(\i_m4stg_frac/n295 ), .IN3(
        n3238), .Q(\i_m4stg_frac/addout[34] ) );
  AO22X1 U3118 ( .IN1(\i_m4stg_frac/n132 ), .IN2(n3240), .IN3(
        \i_m4stg_frac/n297 ), .IN4(n3241), .Q(n3238) );
  OR2X1 U3119 ( .IN1(n3240), .IN2(\i_m4stg_frac/n132 ), .Q(n3241) );
  XNOR3X1 U3120 ( .IN1(\i_m4stg_frac/n297 ), .IN2(\i_m4stg_frac/n132 ), .IN3(
        n3240), .Q(\i_m4stg_frac/addout[33] ) );
  AO22X1 U3121 ( .IN1(\i_m4stg_frac/n134 ), .IN2(n2927), .IN3(
        \i_m4stg_frac/n299 ), .IN4(n3242), .Q(n3240) );
  OR2X1 U3122 ( .IN1(n2927), .IN2(\i_m4stg_frac/n134 ), .Q(n3242) );
  XNOR3X1 U3123 ( .IN1(\i_m4stg_frac/n134 ), .IN2(\i_m4stg_frac/n299 ), .IN3(
        n2927), .Q(\i_m4stg_frac/addout[32] ) );
  AO22X1 U3124 ( .IN1(\i_m4stg_frac/n136 ), .IN2(n3243), .IN3(
        \i_m4stg_frac/n301 ), .IN4(n3244), .Q(n2927) );
  OR2X1 U3125 ( .IN1(n3243), .IN2(\i_m4stg_frac/n136 ), .Q(n3244) );
  XNOR3X1 U3126 ( .IN1(\i_m4stg_frac/n301 ), .IN2(\i_m4stg_frac/n136 ), .IN3(
        n3243), .Q(\i_m4stg_frac/addout[31] ) );
  AO22X1 U3127 ( .IN1(\i_m4stg_frac/n137 ), .IN2(n3245), .IN3(
        \i_m4stg_frac/n302 ), .IN4(n3246), .Q(n3243) );
  OR2X1 U3128 ( .IN1(n3245), .IN2(\i_m4stg_frac/n137 ), .Q(n3246) );
  XNOR3X1 U3129 ( .IN1(\i_m4stg_frac/n137 ), .IN2(\i_m4stg_frac/n302 ), .IN3(
        n3245), .Q(\i_m4stg_frac/addout[30] ) );
  AO22X1 U3130 ( .IN1(\i_m4stg_frac/n138 ), .IN2(n3247), .IN3(
        \i_m4stg_frac/n303 ), .IN4(n3248), .Q(n3245) );
  OR2X1 U3131 ( .IN1(n3247), .IN2(\i_m4stg_frac/n138 ), .Q(n3248) );
  XOR2X1 U3132 ( .IN1(n1165), .IN2(n3249), .Q(\i_m4stg_frac/addout[2] ) );
  XNOR3X1 U3133 ( .IN1(\i_m4stg_frac/n303 ), .IN2(\i_m4stg_frac/n138 ), .IN3(
        n3247), .Q(\i_m4stg_frac/addout[29] ) );
  AO22X1 U3134 ( .IN1(\i_m4stg_frac/n139 ), .IN2(n3250), .IN3(
        \i_m4stg_frac/n304 ), .IN4(n3251), .Q(n3247) );
  OR2X1 U3135 ( .IN1(n3250), .IN2(\i_m4stg_frac/n139 ), .Q(n3251) );
  XNOR3X1 U3136 ( .IN1(\i_m4stg_frac/n139 ), .IN2(\i_m4stg_frac/n304 ), .IN3(
        n3250), .Q(\i_m4stg_frac/addout[28] ) );
  AO22X1 U3137 ( .IN1(\i_m4stg_frac/n140 ), .IN2(n3252), .IN3(
        \i_m4stg_frac/n305 ), .IN4(n3253), .Q(n3250) );
  OR2X1 U3138 ( .IN1(n3252), .IN2(\i_m4stg_frac/n140 ), .Q(n3253) );
  XNOR3X1 U3139 ( .IN1(\i_m4stg_frac/n305 ), .IN2(\i_m4stg_frac/n140 ), .IN3(
        n3252), .Q(\i_m4stg_frac/addout[27] ) );
  AO22X1 U3140 ( .IN1(\i_m4stg_frac/n141 ), .IN2(n3254), .IN3(
        \i_m4stg_frac/n306 ), .IN4(n3255), .Q(n3252) );
  OR2X1 U3141 ( .IN1(n3254), .IN2(\i_m4stg_frac/n141 ), .Q(n3255) );
  XNOR3X1 U3142 ( .IN1(\i_m4stg_frac/n141 ), .IN2(\i_m4stg_frac/n306 ), .IN3(
        n3254), .Q(\i_m4stg_frac/addout[26] ) );
  AO22X1 U3143 ( .IN1(\i_m4stg_frac/n142 ), .IN2(n3256), .IN3(
        \i_m4stg_frac/n307 ), .IN4(n3257), .Q(n3254) );
  OR2X1 U3144 ( .IN1(n3256), .IN2(\i_m4stg_frac/n142 ), .Q(n3257) );
  XNOR3X1 U3145 ( .IN1(\i_m4stg_frac/n307 ), .IN2(\i_m4stg_frac/n142 ), .IN3(
        n3256), .Q(\i_m4stg_frac/addout[25] ) );
  AO22X1 U3146 ( .IN1(\i_m4stg_frac/n143 ), .IN2(n3258), .IN3(
        \i_m4stg_frac/n308 ), .IN4(n3259), .Q(n3256) );
  OR2X1 U3147 ( .IN1(n3258), .IN2(\i_m4stg_frac/n143 ), .Q(n3259) );
  XNOR3X1 U3148 ( .IN1(\i_m4stg_frac/n143 ), .IN2(\i_m4stg_frac/n308 ), .IN3(
        n3258), .Q(\i_m4stg_frac/addout[24] ) );
  AO22X1 U3149 ( .IN1(\i_m4stg_frac/n144 ), .IN2(n3260), .IN3(
        \i_m4stg_frac/n309 ), .IN4(n3261), .Q(n3258) );
  OR2X1 U3150 ( .IN1(n3260), .IN2(\i_m4stg_frac/n144 ), .Q(n3261) );
  XNOR3X1 U3151 ( .IN1(\i_m4stg_frac/n309 ), .IN2(\i_m4stg_frac/n144 ), .IN3(
        n3260), .Q(\i_m4stg_frac/addout[23] ) );
  AO22X1 U3152 ( .IN1(\i_m4stg_frac/n145 ), .IN2(n3262), .IN3(
        \i_m4stg_frac/n310 ), .IN4(n3263), .Q(n3260) );
  OR2X1 U3153 ( .IN1(n3262), .IN2(\i_m4stg_frac/n145 ), .Q(n3263) );
  XNOR3X1 U3154 ( .IN1(\i_m4stg_frac/n145 ), .IN2(\i_m4stg_frac/n310 ), .IN3(
        n3262), .Q(\i_m4stg_frac/addout[22] ) );
  AO22X1 U3155 ( .IN1(\i_m4stg_frac/n146 ), .IN2(n3264), .IN3(
        \i_m4stg_frac/n311 ), .IN4(n3265), .Q(n3262) );
  OR2X1 U3156 ( .IN1(n3264), .IN2(\i_m4stg_frac/n146 ), .Q(n3265) );
  XNOR3X1 U3157 ( .IN1(\i_m4stg_frac/n311 ), .IN2(\i_m4stg_frac/n146 ), .IN3(
        n3264), .Q(\i_m4stg_frac/addout[21] ) );
  AO22X1 U3158 ( .IN1(\i_m4stg_frac/n147 ), .IN2(n3266), .IN3(
        \i_m4stg_frac/n312 ), .IN4(n3267), .Q(n3264) );
  OR2X1 U3159 ( .IN1(n3266), .IN2(\i_m4stg_frac/n147 ), .Q(n3267) );
  XNOR3X1 U3160 ( .IN1(\i_m4stg_frac/n147 ), .IN2(\i_m4stg_frac/n312 ), .IN3(
        n3266), .Q(\i_m4stg_frac/addout[20] ) );
  AO22X1 U3161 ( .IN1(\i_m4stg_frac/n148 ), .IN2(n3268), .IN3(
        \i_m4stg_frac/n313 ), .IN4(n3269), .Q(n3266) );
  OR2X1 U3162 ( .IN1(n3268), .IN2(\i_m4stg_frac/n148 ), .Q(n3269) );
  NOR2X0 U3163 ( .IN1(n3249), .IN2(n3270), .QN(\i_m4stg_frac/addout[1] ) );
  OA21X1 U3164 ( .IN1(\i_m4stg_frac/n332 ), .IN2(\i_m4stg_frac/n1329 ), .IN3(
        \i_m4stg_frac/n331 ), .Q(n3270) );
  XNOR3X1 U3165 ( .IN1(\i_m4stg_frac/n313 ), .IN2(\i_m4stg_frac/n148 ), .IN3(
        n3268), .Q(\i_m4stg_frac/addout[19] ) );
  AO22X1 U3166 ( .IN1(\i_m4stg_frac/n149 ), .IN2(n3271), .IN3(
        \i_m4stg_frac/n314 ), .IN4(n3272), .Q(n3268) );
  OR2X1 U3167 ( .IN1(n3271), .IN2(\i_m4stg_frac/n149 ), .Q(n3272) );
  XNOR3X1 U3168 ( .IN1(\i_m4stg_frac/n149 ), .IN2(\i_m4stg_frac/n314 ), .IN3(
        n3271), .Q(\i_m4stg_frac/addout[18] ) );
  AO22X1 U3169 ( .IN1(\i_m4stg_frac/n150 ), .IN2(n3273), .IN3(
        \i_m4stg_frac/n315 ), .IN4(n3274), .Q(n3271) );
  OR2X1 U3170 ( .IN1(n3273), .IN2(\i_m4stg_frac/n150 ), .Q(n3274) );
  XNOR3X1 U3171 ( .IN1(\i_m4stg_frac/n315 ), .IN2(\i_m4stg_frac/n150 ), .IN3(
        n3273), .Q(\i_m4stg_frac/addout[17] ) );
  OR2X1 U3172 ( .IN1(\i_m4stg_frac/n316 ), .IN2(n3275), .Q(n3273) );
  XOR2X1 U3173 ( .IN1(\i_m4stg_frac/n316 ), .IN2(n3275), .Q(
        \i_m4stg_frac/addout[16] ) );
  OA22X1 U3174 ( .IN1(n3276), .IN2(\i_m4stg_frac/n152 ), .IN3(n3277), .IN4(
        \i_m4stg_frac/n317 ), .Q(n3275) );
  AND2X1 U3175 ( .IN1(\i_m4stg_frac/n152 ), .IN2(n3276), .Q(n3277) );
  XNOR3X1 U3176 ( .IN1(\i_m4stg_frac/n152 ), .IN2(\i_m4stg_frac/n317 ), .IN3(
        n3276), .Q(\i_m4stg_frac/addout[15] ) );
  AO22X1 U3177 ( .IN1(\i_m4stg_frac/n153 ), .IN2(n3278), .IN3(
        \i_m4stg_frac/n318 ), .IN4(n3279), .Q(n3276) );
  OR2X1 U3178 ( .IN1(n3278), .IN2(\i_m4stg_frac/n153 ), .Q(n3279) );
  XNOR3X1 U3179 ( .IN1(\i_m4stg_frac/n153 ), .IN2(\i_m4stg_frac/n318 ), .IN3(
        n3278), .Q(\i_m4stg_frac/addout[14] ) );
  AO22X1 U3180 ( .IN1(\i_m4stg_frac/n154 ), .IN2(n3280), .IN3(
        \i_m4stg_frac/n319 ), .IN4(n3281), .Q(n3278) );
  OR2X1 U3181 ( .IN1(n3280), .IN2(\i_m4stg_frac/n154 ), .Q(n3281) );
  XNOR3X1 U3182 ( .IN1(\i_m4stg_frac/n154 ), .IN2(\i_m4stg_frac/n319 ), .IN3(
        n3280), .Q(\i_m4stg_frac/addout[13] ) );
  AO22X1 U3183 ( .IN1(\i_m4stg_frac/n155 ), .IN2(n3282), .IN3(
        \i_m4stg_frac/n320 ), .IN4(n3283), .Q(n3280) );
  OR2X1 U3184 ( .IN1(n3282), .IN2(\i_m4stg_frac/n155 ), .Q(n3283) );
  XNOR3X1 U3185 ( .IN1(\i_m4stg_frac/n155 ), .IN2(\i_m4stg_frac/n320 ), .IN3(
        n3282), .Q(\i_m4stg_frac/addout[12] ) );
  AO22X1 U3186 ( .IN1(\i_m4stg_frac/n156 ), .IN2(n3284), .IN3(
        \i_m4stg_frac/n321 ), .IN4(n3285), .Q(n3282) );
  OR2X1 U3187 ( .IN1(n3284), .IN2(\i_m4stg_frac/n156 ), .Q(n3285) );
  XNOR3X1 U3188 ( .IN1(\i_m4stg_frac/n156 ), .IN2(\i_m4stg_frac/n321 ), .IN3(
        n3284), .Q(\i_m4stg_frac/addout[11] ) );
  AO22X1 U3189 ( .IN1(\i_m4stg_frac/n157 ), .IN2(n3286), .IN3(
        \i_m4stg_frac/n322 ), .IN4(n3287), .Q(n3284) );
  OR2X1 U3190 ( .IN1(n3286), .IN2(\i_m4stg_frac/n157 ), .Q(n3287) );
  XNOR3X1 U3191 ( .IN1(\i_m4stg_frac/n157 ), .IN2(\i_m4stg_frac/n322 ), .IN3(
        n3286), .Q(\i_m4stg_frac/addout[10] ) );
  AO22X1 U3192 ( .IN1(\i_m4stg_frac/n158 ), .IN2(n3154), .IN3(
        \i_m4stg_frac/n323 ), .IN4(n3288), .Q(n3286) );
  OR2X1 U3193 ( .IN1(n3154), .IN2(\i_m4stg_frac/n158 ), .Q(n3288) );
  AO22X1 U3194 ( .IN1(\i_m4stg_frac/n159 ), .IN2(n3155), .IN3(
        \i_m4stg_frac/n324 ), .IN4(n3289), .Q(n3154) );
  OR2X1 U3195 ( .IN1(n3155), .IN2(\i_m4stg_frac/n159 ), .Q(n3289) );
  AO22X1 U3196 ( .IN1(\i_m4stg_frac/n160 ), .IN2(n3156), .IN3(
        \i_m4stg_frac/n325 ), .IN4(n3290), .Q(n3155) );
  OR2X1 U3197 ( .IN1(n3156), .IN2(\i_m4stg_frac/n160 ), .Q(n3290) );
  AO22X1 U3198 ( .IN1(\i_m4stg_frac/n161 ), .IN2(n3166), .IN3(
        \i_m4stg_frac/n326 ), .IN4(n3291), .Q(n3156) );
  OR2X1 U3199 ( .IN1(n3166), .IN2(\i_m4stg_frac/n161 ), .Q(n3291) );
  AO22X1 U3200 ( .IN1(\i_m4stg_frac/n162 ), .IN2(n3187), .IN3(
        \i_m4stg_frac/n327 ), .IN4(n3292), .Q(n3166) );
  OR2X1 U3201 ( .IN1(n3187), .IN2(\i_m4stg_frac/n162 ), .Q(n3292) );
  AO22X1 U3202 ( .IN1(\i_m4stg_frac/n163 ), .IN2(n3208), .IN3(
        \i_m4stg_frac/n328 ), .IN4(n3293), .Q(n3187) );
  OR2X1 U3203 ( .IN1(n3208), .IN2(\i_m4stg_frac/n163 ), .Q(n3293) );
  AO22X1 U3204 ( .IN1(\i_m4stg_frac/n164 ), .IN2(n3229), .IN3(
        \i_m4stg_frac/n329 ), .IN4(n3294), .Q(n3208) );
  OR2X1 U3205 ( .IN1(n3229), .IN2(\i_m4stg_frac/n164 ), .Q(n3294) );
  NAND2X0 U3206 ( .IN1(n3249), .IN2(n1165), .QN(n3229) );
  NOR3X0 U3207 ( .IN1(\i_m4stg_frac/n331 ), .IN2(\i_m4stg_frac/n332 ), .IN3(
        \i_m4stg_frac/n1329 ), .QN(n3249) );
  XOR2X1 U3208 ( .IN1(\i_m4stg_frac/n332 ), .IN2(\i_m4stg_frac/n1329 ), .Q(
        \i_m4stg_frac/addout[0] ) );
  NOR3X0 U3209 ( .IN1(n2342), .IN2(se_mul64), .IN3(n2341), .QN(
        \i_m4stg_frac/a2cot_dff/N19 ) );
  XOR3X1 U3210 ( .IN1(n2350), .IN2(n2352), .IN3(n2351), .Q(n2341) );
  XNOR3X1 U3211 ( .IN1(\i_m4stg_frac/n965 ), .IN2(\i_m4stg_frac/n811 ), .IN3(
        n2359), .Q(n2351) );
  XOR3X1 U3212 ( .IN1(\i_m4stg_frac/ps[48] ), .IN2(\i_m4stg_frac/pc[47] ), 
        .IN3(\i_m4stg_frac/n652 ), .Q(n2359) );
  AO22X1 U3213 ( .IN1(n3295), .IN2(n929), .IN3(n3296), .IN4(n1189), .Q(n2352)
         );
  OR2X1 U3214 ( .IN1(n929), .IN2(n3295), .Q(n3296) );
  OAI22X1 U3215 ( .IN1(n2245), .IN2(n2246), .IN3(n2247), .IN4(n3297), .QN(
        n2342) );
  AND2X1 U3216 ( .IN1(n2245), .IN2(n2246), .Q(n3297) );
  AO22X1 U3217 ( .IN1(n2495), .IN2(n2494), .IN3(n3298), .IN4(n1331), .Q(n2247)
         );
  OR2X1 U3218 ( .IN1(n2494), .IN2(n2495), .Q(n3298) );
  AO22X1 U3219 ( .IN1(\i_m4stg_frac/pc[44] ), .IN2(n1112), .IN3(
        \i_m4stg_frac/ps[45] ), .IN4(n3299), .Q(n2494) );
  OR2X1 U3220 ( .IN1(n1112), .IN2(\i_m4stg_frac/pc[44] ), .Q(n3299) );
  XNOR3X1 U3221 ( .IN1(\i_m4stg_frac/ps[46] ), .IN2(\i_m4stg_frac/pc[45] ), 
        .IN3(\i_m4stg_frac/n969 ), .Q(n2495) );
  AO22X1 U3222 ( .IN1(\i_m4stg_frac/pc[45] ), .IN2(n1192), .IN3(
        \i_m4stg_frac/ps[46] ), .IN4(n3300), .Q(n2246) );
  OR2X1 U3223 ( .IN1(n1192), .IN2(\i_m4stg_frac/pc[45] ), .Q(n3300) );
  XOR3X1 U3224 ( .IN1(n1189), .IN2(n929), .IN3(n3295), .Q(n2245) );
  OA21X1 U3225 ( .IN1(\i_m4stg_frac/ps[47] ), .IN2(\i_m4stg_frac/pc[46] ), 
        .IN3(n2350), .Q(n3295) );
  NAND2X0 U3226 ( .IN1(\i_m4stg_frac/ps[47] ), .IN2(\i_m4stg_frac/pc[46] ), 
        .QN(n2350) );
  XOR3X1 U3227 ( .IN1(n3301), .IN2(n3302), .IN3(n3303), .Q(
        \i_m4stg_frac/a1sum[9] ) );
  XNOR3X1 U3228 ( .IN1(n3304), .IN2(n3305), .IN3(n3306), .Q(
        \i_m4stg_frac/a1sum[8] ) );
  XOR2X1 U3229 ( .IN1(n3307), .IN2(n3308), .Q(\i_m4stg_frac/a1sum[7] ) );
  XOR2X1 U3230 ( .IN1(n3309), .IN2(n3310), .Q(\i_m4stg_frac/a1sum[79] ) );
  XOR2X1 U3231 ( .IN1(n3310), .IN2(n3311), .Q(\i_m4stg_frac/a1sum[78] ) );
  NOR2X0 U3232 ( .IN1(n3312), .IN2(n3313), .QN(n3311) );
  XOR3X1 U3233 ( .IN1(n3314), .IN2(n3315), .IN3(n3316), .Q(
        \i_m4stg_frac/a1sum[77] ) );
  XNOR2X1 U3234 ( .IN1(n3317), .IN2(n3318), .Q(\i_m4stg_frac/a1sum[76] ) );
  NAND2X0 U3235 ( .IN1(n3319), .IN2(n3320), .QN(n3318) );
  XOR2X1 U3236 ( .IN1(n3321), .IN2(n3322), .Q(\i_m4stg_frac/a1sum[75] ) );
  AND2X1 U3237 ( .IN1(n3323), .IN2(n3324), .Q(n3321) );
  XOR3X1 U3238 ( .IN1(n3325), .IN2(n3326), .IN3(n3327), .Q(
        \i_m4stg_frac/a1sum[74] ) );
  XNOR2X1 U3239 ( .IN1(n3328), .IN2(n3329), .Q(\i_m4stg_frac/a1sum[73] ) );
  NOR2X0 U3240 ( .IN1(n3330), .IN2(n3331), .QN(n3329) );
  XNOR3X1 U3241 ( .IN1(n3332), .IN2(n3333), .IN3(n3334), .Q(
        \i_m4stg_frac/a1sum[72] ) );
  XOR3X1 U3242 ( .IN1(n3335), .IN2(n3336), .IN3(n3337), .Q(
        \i_m4stg_frac/a1sum[71] ) );
  XOR3X1 U3243 ( .IN1(n3338), .IN2(n3339), .IN3(n3340), .Q(
        \i_m4stg_frac/a1sum[70] ) );
  XOR2X1 U3244 ( .IN1(n3341), .IN2(n3342), .Q(\i_m4stg_frac/a1sum[6] ) );
  XOR3X1 U3245 ( .IN1(n3343), .IN2(n3344), .IN3(n3345), .Q(
        \i_m4stg_frac/a1sum[69] ) );
  XOR3X1 U3246 ( .IN1(n3346), .IN2(n3347), .IN3(n3348), .Q(
        \i_m4stg_frac/a1sum[68] ) );
  XOR3X1 U3247 ( .IN1(n3349), .IN2(n3350), .IN3(n3351), .Q(
        \i_m4stg_frac/a1sum[67] ) );
  XOR3X1 U3248 ( .IN1(n3352), .IN2(n3353), .IN3(n3354), .Q(
        \i_m4stg_frac/a1sum[66] ) );
  XOR3X1 U3249 ( .IN1(n3355), .IN2(n3356), .IN3(n3357), .Q(
        \i_m4stg_frac/a1sum[65] ) );
  XOR3X1 U3250 ( .IN1(n3358), .IN2(n3359), .IN3(n3360), .Q(
        \i_m4stg_frac/a1sum[64] ) );
  XOR3X1 U3251 ( .IN1(n3361), .IN2(n3362), .IN3(n3363), .Q(
        \i_m4stg_frac/a1sum[63] ) );
  XOR3X1 U3252 ( .IN1(n3364), .IN2(n3365), .IN3(n3366), .Q(
        \i_m4stg_frac/a1sum[62] ) );
  XOR3X1 U3253 ( .IN1(n3367), .IN2(n3368), .IN3(n3369), .Q(
        \i_m4stg_frac/a1sum[61] ) );
  XOR3X1 U3254 ( .IN1(n3370), .IN2(n3371), .IN3(n3372), .Q(
        \i_m4stg_frac/a1sum[60] ) );
  XOR2X1 U3255 ( .IN1(n3373), .IN2(n3374), .Q(\i_m4stg_frac/a1sum[5] ) );
  XOR3X1 U3256 ( .IN1(n3375), .IN2(n3376), .IN3(n3377), .Q(
        \i_m4stg_frac/a1sum[59] ) );
  XOR3X1 U3257 ( .IN1(n3378), .IN2(n3379), .IN3(n3380), .Q(
        \i_m4stg_frac/a1sum[58] ) );
  XOR3X1 U3258 ( .IN1(n3381), .IN2(n3382), .IN3(n3383), .Q(
        \i_m4stg_frac/a1sum[57] ) );
  XOR3X1 U3259 ( .IN1(n3384), .IN2(n3385), .IN3(n3386), .Q(
        \i_m4stg_frac/a1sum[56] ) );
  XOR3X1 U3260 ( .IN1(n3387), .IN2(n3388), .IN3(n3389), .Q(
        \i_m4stg_frac/a1sum[55] ) );
  XOR3X1 U3261 ( .IN1(n3390), .IN2(n3391), .IN3(n3392), .Q(
        \i_m4stg_frac/a1sum[54] ) );
  XOR3X1 U3262 ( .IN1(n3393), .IN2(n3394), .IN3(n3395), .Q(
        \i_m4stg_frac/a1sum[53] ) );
  XOR3X1 U3263 ( .IN1(n3396), .IN2(n3397), .IN3(n3398), .Q(
        \i_m4stg_frac/a1sum[52] ) );
  XOR3X1 U3264 ( .IN1(n3399), .IN2(n3400), .IN3(n3401), .Q(
        \i_m4stg_frac/a1sum[51] ) );
  XOR3X1 U3265 ( .IN1(n3402), .IN2(n3403), .IN3(n3404), .Q(
        \i_m4stg_frac/a1sum[50] ) );
  XOR2X1 U3266 ( .IN1(n3405), .IN2(n3406), .Q(\i_m4stg_frac/a1sum[4] ) );
  XOR3X1 U3267 ( .IN1(n3407), .IN2(n3408), .IN3(n3409), .Q(
        \i_m4stg_frac/a1sum[49] ) );
  XOR3X1 U3268 ( .IN1(n3410), .IN2(n3411), .IN3(n3412), .Q(
        \i_m4stg_frac/a1sum[48] ) );
  XOR3X1 U3269 ( .IN1(n3413), .IN2(n3414), .IN3(n3415), .Q(
        \i_m4stg_frac/a1sum[47] ) );
  XOR3X1 U3270 ( .IN1(n3416), .IN2(n3417), .IN3(n3418), .Q(
        \i_m4stg_frac/a1sum[46] ) );
  XOR3X1 U3271 ( .IN1(n3419), .IN2(n3420), .IN3(n3421), .Q(
        \i_m4stg_frac/a1sum[45] ) );
  XOR3X1 U3272 ( .IN1(n3422), .IN2(n3423), .IN3(n3424), .Q(
        \i_m4stg_frac/a1sum[44] ) );
  XOR3X1 U3273 ( .IN1(n3425), .IN2(n3426), .IN3(n3427), .Q(
        \i_m4stg_frac/a1sum[43] ) );
  XOR3X1 U3274 ( .IN1(n3428), .IN2(n3429), .IN3(n3430), .Q(
        \i_m4stg_frac/a1sum[42] ) );
  XOR3X1 U3275 ( .IN1(n3431), .IN2(n3432), .IN3(n3433), .Q(
        \i_m4stg_frac/a1sum[41] ) );
  XOR3X1 U3276 ( .IN1(n3434), .IN2(n3435), .IN3(n3436), .Q(
        \i_m4stg_frac/a1sum[40] ) );
  XOR3X1 U3277 ( .IN1(n3437), .IN2(n3438), .IN3(n3439), .Q(
        \i_m4stg_frac/a1sum[3] ) );
  XOR3X1 U3278 ( .IN1(n3440), .IN2(n3441), .IN3(n3442), .Q(
        \i_m4stg_frac/a1sum[39] ) );
  XOR3X1 U3279 ( .IN1(n3443), .IN2(n3444), .IN3(n3445), .Q(
        \i_m4stg_frac/a1sum[38] ) );
  XOR3X1 U3280 ( .IN1(n3446), .IN2(n3447), .IN3(n3448), .Q(
        \i_m4stg_frac/a1sum[37] ) );
  XOR3X1 U3281 ( .IN1(n3449), .IN2(n3450), .IN3(n3451), .Q(
        \i_m4stg_frac/a1sum[36] ) );
  XOR3X1 U3282 ( .IN1(n3452), .IN2(n3453), .IN3(n3454), .Q(
        \i_m4stg_frac/a1sum[35] ) );
  XOR3X1 U3283 ( .IN1(n3455), .IN2(n3456), .IN3(n3457), .Q(
        \i_m4stg_frac/a1sum[34] ) );
  XOR3X1 U3284 ( .IN1(n3458), .IN2(n3459), .IN3(n3460), .Q(
        \i_m4stg_frac/a1sum[33] ) );
  XOR3X1 U3285 ( .IN1(n3461), .IN2(n3462), .IN3(n3463), .Q(
        \i_m4stg_frac/a1sum[32] ) );
  XOR3X1 U3286 ( .IN1(n3464), .IN2(n3465), .IN3(n3466), .Q(
        \i_m4stg_frac/a1sum[31] ) );
  XOR3X1 U3287 ( .IN1(n3467), .IN2(n3468), .IN3(n3469), .Q(
        \i_m4stg_frac/a1sum[30] ) );
  OA21X1 U3288 ( .IN1(n3470), .IN2(n3471), .IN3(n3438), .Q(
        \i_m4stg_frac/a1sum[2] ) );
  XOR3X1 U3289 ( .IN1(n3472), .IN2(n3473), .IN3(n3474), .Q(
        \i_m4stg_frac/a1sum[29] ) );
  XOR3X1 U3290 ( .IN1(n3475), .IN2(n3476), .IN3(n3477), .Q(
        \i_m4stg_frac/a1sum[28] ) );
  XOR3X1 U3291 ( .IN1(n3478), .IN2(n3479), .IN3(n3480), .Q(
        \i_m4stg_frac/a1sum[27] ) );
  XOR3X1 U3292 ( .IN1(n3481), .IN2(n3482), .IN3(n3483), .Q(
        \i_m4stg_frac/a1sum[26] ) );
  XOR3X1 U3293 ( .IN1(n3484), .IN2(n3485), .IN3(n3486), .Q(
        \i_m4stg_frac/a1sum[25] ) );
  XOR3X1 U3294 ( .IN1(n3487), .IN2(n3488), .IN3(n3489), .Q(
        \i_m4stg_frac/a1sum[24] ) );
  XOR3X1 U3295 ( .IN1(n3490), .IN2(n3491), .IN3(n3492), .Q(
        \i_m4stg_frac/a1sum[23] ) );
  XOR3X1 U3296 ( .IN1(n3493), .IN2(n3494), .IN3(n3495), .Q(
        \i_m4stg_frac/a1sum[22] ) );
  XOR3X1 U3297 ( .IN1(n3496), .IN2(n3497), .IN3(n3498), .Q(
        \i_m4stg_frac/a1sum[21] ) );
  XOR3X1 U3298 ( .IN1(n3499), .IN2(n3500), .IN3(n3501), .Q(
        \i_m4stg_frac/a1sum[20] ) );
  OA21X1 U3299 ( .IN1(n3502), .IN2(n3503), .IN3(n3504), .Q(
        \i_m4stg_frac/a1sum[1] ) );
  AND2X1 U3300 ( .IN1(n3505), .IN2(n3506), .Q(n3502) );
  XOR3X1 U3301 ( .IN1(n3507), .IN2(n3508), .IN3(n3509), .Q(
        \i_m4stg_frac/a1sum[19] ) );
  XOR3X1 U3302 ( .IN1(n3510), .IN2(n3511), .IN3(n3512), .Q(
        \i_m4stg_frac/a1sum[18] ) );
  XOR3X1 U3303 ( .IN1(n3513), .IN2(n3514), .IN3(n3515), .Q(
        \i_m4stg_frac/a1sum[17] ) );
  XOR3X1 U3304 ( .IN1(n3516), .IN2(n3517), .IN3(n3518), .Q(
        \i_m4stg_frac/a1sum[16] ) );
  XOR3X1 U3305 ( .IN1(n3519), .IN2(n3520), .IN3(n3521), .Q(
        \i_m4stg_frac/a1sum[15] ) );
  XOR3X1 U3306 ( .IN1(n3522), .IN2(n3523), .IN3(n3524), .Q(
        \i_m4stg_frac/a1sum[14] ) );
  XOR3X1 U3307 ( .IN1(n3525), .IN2(n3526), .IN3(n3527), .Q(
        \i_m4stg_frac/a1sum[13] ) );
  XOR3X1 U3308 ( .IN1(n3528), .IN2(n3529), .IN3(n3530), .Q(
        \i_m4stg_frac/a1sum[12] ) );
  XOR2X1 U3309 ( .IN1(n3531), .IN2(n3532), .Q(\i_m4stg_frac/a1sum[11] ) );
  XOR3X1 U3310 ( .IN1(n3533), .IN2(n3534), .IN3(n3535), .Q(
        \i_m4stg_frac/a1sum[10] ) );
  NOR2X0 U3311 ( .IN1(\i_m4stg_frac/n676 ), .IN2(n3505), .QN(
        \i_m4stg_frac/a1sum[0] ) );
  AO22X1 U3312 ( .IN1(n3536), .IN2(n3537), .IN3(n3303), .IN4(n3538), .Q(
        \i_m4stg_frac/a1cout[9] ) );
  NAND2X0 U3313 ( .IN1(n3302), .IN2(n3301), .QN(n3538) );
  INVX0 U3314 ( .INP(n3536), .ZN(n3302) );
  XOR3X1 U3315 ( .IN1(n3539), .IN2(n3540), .IN3(n3541), .Q(n3303) );
  INVX0 U3316 ( .INP(n3301), .ZN(n3537) );
  OA22X1 U3317 ( .IN1(n3542), .IN2(n3543), .IN3(n3544), .IN4(n3545), .Q(n3301)
         );
  AND2X1 U3318 ( .IN1(n3543), .IN2(n3542), .Q(n3545) );
  NAND2X0 U3319 ( .IN1(n3546), .IN2(n3547), .QN(n3536) );
  NAND3X0 U3320 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(n3548), .IN3(n3549), .QN(
        n3547) );
  INVX0 U3321 ( .INP(n3550), .ZN(n3549) );
  OAI21X1 U3322 ( .IN1(n3548), .IN2(n1034), .IN3(n3551), .QN(n3546) );
  OAI22X1 U3323 ( .IN1(n3306), .IN2(n3305), .IN3(n3304), .IN4(n3552), .QN(
        \i_m4stg_frac/a1cout[8] ) );
  AND2X1 U3324 ( .IN1(n3305), .IN2(n3306), .Q(n3552) );
  AOI22X1 U3325 ( .IN1(n3553), .IN2(n3554), .IN3(n3555), .IN4(n3556), .QN(
        n3305) );
  OR2X1 U3326 ( .IN1(n3554), .IN2(n3553), .Q(n3556) );
  XOR3X1 U3327 ( .IN1(n3544), .IN2(n3543), .IN3(n3542), .Q(n3306) );
  XNOR3X1 U3328 ( .IN1(n3557), .IN2(n3558), .IN3(n3559), .Q(n3542) );
  AOI22X1 U3329 ( .IN1(n3560), .IN2(n3561), .IN3(n3562), .IN4(n3563), .QN(
        n3543) );
  OR2X1 U3330 ( .IN1(n3561), .IN2(n3560), .Q(n3562) );
  XOR2X1 U3331 ( .IN1(n3564), .IN2(n3548), .Q(n3544) );
  NAND2X0 U3332 ( .IN1(n3565), .IN2(n3566), .QN(n3548) );
  MUX21X1 U3333 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1468 ), .Q(n3566) );
  MUX21X1 U3334 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1469 ), .Q(n3565) );
  NAND3X0 U3335 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(n1116), .IN3(
        \i_m4stg_frac/n665 ), .QN(n3564) );
  NOR2X0 U3336 ( .IN1(n3308), .IN2(n3307), .QN(\i_m4stg_frac/a1cout[7] ) );
  AO22X1 U3337 ( .IN1(n3571), .IN2(n3572), .IN3(n3573), .IN4(n3574), .Q(n3307)
         );
  NAND2X0 U3338 ( .IN1(n3575), .IN2(n3576), .QN(n3573) );
  INVX0 U3339 ( .INP(n3575), .ZN(n3572) );
  INVX0 U3340 ( .INP(n3576), .ZN(n3571) );
  XNOR3X1 U3341 ( .IN1(n3555), .IN2(n3554), .IN3(n3553), .Q(n3308) );
  XOR3X1 U3342 ( .IN1(n3563), .IN2(n3561), .IN3(n3560), .Q(n3553) );
  NAND2X0 U3343 ( .IN1(n3577), .IN2(n3578), .QN(n3560) );
  MUX21X1 U3344 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1472 ), .Q(n3578) );
  MUX21X1 U3345 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1471 ), .Q(n3577) );
  NAND2X0 U3346 ( .IN1(n3583), .IN2(n3584), .QN(n3561) );
  MUX21X1 U3347 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1474 ), .Q(n3584) );
  MUX21X1 U3348 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1473 ), .Q(n3583) );
  NAND2X0 U3349 ( .IN1(n3589), .IN2(n3590), .QN(n3563) );
  MUX21X1 U3350 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1469 ), .Q(n3590) );
  MUX21X1 U3351 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1470 ), .Q(n3589) );
  AO22X1 U3352 ( .IN1(n3595), .IN2(n3596), .IN3(n3597), .IN4(n3598), .Q(n3554)
         );
  OR2X1 U3353 ( .IN1(n3596), .IN2(n3595), .Q(n3597) );
  AND2X1 U3354 ( .IN1(n3599), .IN2(n3304), .Q(n3555) );
  NAND3X0 U3355 ( .IN1(n3600), .IN2(n3601), .IN3(n3602), .QN(n3304) );
  AO21X1 U3356 ( .IN1(n3602), .IN2(n3600), .IN3(n3601), .Q(n3599) );
  NAND2X0 U3357 ( .IN1(n3603), .IN2(n3604), .QN(n3601) );
  MUX21X1 U3358 ( .IN1(n3605), .IN2(n3570), .S(\i_m4stg_frac/n1468 ), .Q(n3604) );
  NAND2X0 U3359 ( .IN1(n3606), .IN2(n912), .QN(n3605) );
  MUX21X1 U3360 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1467 ), .Q(n3603) );
  NAND2X0 U3361 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(\i_m4stg_frac/n668 ), .QN(
        n3600) );
  NOR2X0 U3362 ( .IN1(n3309), .IN2(n3310), .QN(\i_m4stg_frac/a1cout[79] ) );
  AND3X1 U3363 ( .IN1(n3310), .IN2(n3607), .IN3(n3608), .Q(
        \i_m4stg_frac/a1cout[78] ) );
  OA21X1 U3364 ( .IN1(n3313), .IN2(\i_m4stg_frac/n656 ), .IN3(n3609), .Q(n3310) );
  AO21X1 U3365 ( .IN1(n3316), .IN2(n3314), .IN3(n3315), .Q(
        \i_m4stg_frac/a1cout[77] ) );
  XOR2X1 U3366 ( .IN1(n3607), .IN2(n3608), .Q(n3316) );
  INVX0 U3367 ( .INP(n3312), .ZN(n3607) );
  OAI22X1 U3368 ( .IN1(n3319), .IN2(n3317), .IN3(n3317), .IN4(n3320), .QN(
        \i_m4stg_frac/a1cout[76] ) );
  NAND2X0 U3369 ( .IN1(n3322), .IN2(n3610), .QN(n3320) );
  OA21X1 U3370 ( .IN1(n3611), .IN2(n3612), .IN3(n3314), .Q(n3317) );
  OAI21X1 U3371 ( .IN1(n3315), .IN2(n3613), .IN3(n3611), .QN(n3314) );
  NOR2X0 U3372 ( .IN1(n3612), .IN2(n3608), .QN(n3613) );
  AND2X1 U3373 ( .IN1(n3608), .IN2(n3612), .Q(n3315) );
  AO21X1 U3374 ( .IN1(n3614), .IN2(n3615), .IN3(n3616), .Q(n3612) );
  NAND2X0 U3375 ( .IN1(n3617), .IN2(n3618), .QN(n3319) );
  OAI22X1 U3376 ( .IN1(n3322), .IN2(n3324), .IN3(n3322), .IN4(n3323), .QN(
        \i_m4stg_frac/a1cout[75] ) );
  INVX0 U3377 ( .INP(n3619), .ZN(n3323) );
  NAND2X0 U3378 ( .IN1(n3618), .IN2(n3620), .QN(n3324) );
  XOR3X1 U3379 ( .IN1(n3621), .IN2(n3610), .IN3(n3622), .Q(n3322) );
  XOR2X1 U3380 ( .IN1(n3617), .IN2(n3623), .Q(n3622) );
  OA21X1 U3381 ( .IN1(n3327), .IN2(n3326), .IN3(n3325), .Q(
        \i_m4stg_frac/a1cout[74] ) );
  AOI21X1 U3382 ( .IN1(n3624), .IN2(n3617), .IN3(n3619), .QN(n3325) );
  NOR2X0 U3383 ( .IN1(n3624), .IN2(n3617), .QN(n3619) );
  AND2X1 U3384 ( .IN1(n3625), .IN2(n3626), .Q(n3617) );
  MUX21X1 U3385 ( .IN1(n3627), .IN2(n934), .S(\i_m4stg_frac/n662 ), .Q(n3625)
         );
  NAND2X0 U3386 ( .IN1(\i_m4stg_frac/n1530 ), .IN2(n934), .QN(n3627) );
  XOR2X1 U3387 ( .IN1(n3628), .IN2(n3620), .Q(n3624) );
  NOR2X0 U3388 ( .IN1(n3629), .IN2(n3630), .QN(n3620) );
  AND2X1 U3389 ( .IN1(n3631), .IN2(n3618), .Q(n3326) );
  NOR2X0 U3390 ( .IN1(n3328), .IN2(n3632), .QN(n3327) );
  AO22X1 U3391 ( .IN1(n3328), .IN2(n3331), .IN3(n3330), .IN4(n3328), .Q(
        \i_m4stg_frac/a1cout[73] ) );
  AND2X1 U3392 ( .IN1(n3332), .IN2(n3633), .Q(n3330) );
  AND2X1 U3393 ( .IN1(n3634), .IN2(n3618), .Q(n3331) );
  XOR3X1 U3394 ( .IN1(n3635), .IN2(n3621), .IN3(n3636), .Q(n3328) );
  XOR2X1 U3395 ( .IN1(n3637), .IN2(n3632), .Q(n3635) );
  XOR2X1 U3396 ( .IN1(n3630), .IN2(n3638), .Q(n3632) );
  OAI22X1 U3397 ( .IN1(n3332), .IN2(n3333), .IN3(n3334), .IN4(n3639), .QN(
        \i_m4stg_frac/a1cout[72] ) );
  AND2X1 U3398 ( .IN1(n3332), .IN2(n3333), .Q(n3639) );
  MUX21X1 U3399 ( .IN1(n3640), .IN2(n3641), .S(n3642), .Q(n3334) );
  INVX0 U3400 ( .INP(n3643), .ZN(n3642) );
  NAND2X0 U3401 ( .IN1(n3644), .IN2(n3618), .QN(n3333) );
  XOR3X1 U3402 ( .IN1(n3645), .IN2(n3621), .IN3(n3633), .Q(n3332) );
  AO221X1 U3403 ( .IN1(n3646), .IN2(n914), .IN3(n3638), .IN4(n3551), .IN5(
        n3636), .Q(n3633) );
  INVX0 U3404 ( .INP(n3631), .ZN(n3636) );
  NAND3X0 U3405 ( .IN1(n3629), .IN2(n3647), .IN3(n3648), .QN(n3631) );
  NAND2X0 U3406 ( .IN1(n3649), .IN2(n914), .QN(n3648) );
  INVX0 U3407 ( .INP(n3647), .ZN(n3551) );
  XOR2X1 U3408 ( .IN1(n3634), .IN2(n3623), .Q(n3645) );
  AO21X1 U3409 ( .IN1(n3650), .IN2(n3651), .IN3(n3646), .Q(n3634) );
  AO22X1 U3410 ( .IN1(n3335), .IN2(n3336), .IN3(n3337), .IN4(n3652), .Q(
        \i_m4stg_frac/a1cout[71] ) );
  NAND2X0 U3411 ( .IN1(n3653), .IN2(n3339), .QN(n3652) );
  XOR2X1 U3412 ( .IN1(n3643), .IN2(n3641), .Q(n3337) );
  INVX0 U3413 ( .INP(n3654), .ZN(n3641) );
  XOR3X1 U3414 ( .IN1(n3655), .IN2(n3621), .IN3(n3644), .Q(n3643) );
  AO21X1 U3415 ( .IN1(n3656), .IN2(n3650), .IN3(n3646), .Q(n3644) );
  XOR2X1 U3416 ( .IN1(n3637), .IN2(n3640), .Q(n3655) );
  XOR2X1 U3417 ( .IN1(n3602), .IN2(n3657), .Q(n3640) );
  INVX0 U3418 ( .INP(n3653), .ZN(n3335) );
  MUX21X1 U3419 ( .IN1(n3658), .IN2(n3654), .S(n3659), .Q(n3653) );
  AO22X1 U3420 ( .IN1(n3660), .IN2(n3336), .IN3(n3338), .IN4(n3661), .Q(
        \i_m4stg_frac/a1cout[70] ) );
  NAND2X0 U3421 ( .IN1(n3340), .IN2(n3339), .QN(n3661) );
  XOR2X1 U3422 ( .IN1(n3659), .IN2(n3658), .Q(n3338) );
  AOI22X1 U3423 ( .IN1(n3662), .IN2(n3663), .IN3(n3664), .IN4(n3665), .QN(
        n3658) );
  NAND2X0 U3424 ( .IN1(n3666), .IN2(n3667), .QN(n3664) );
  XNOR3X1 U3425 ( .IN1(n3668), .IN2(n3637), .IN3(n3654), .Q(n3659) );
  XOR2X1 U3426 ( .IN1(n3657), .IN2(n3656), .Q(n3654) );
  AO21X1 U3427 ( .IN1(n3669), .IN2(n3670), .IN3(n3671), .Q(n3656) );
  INVX0 U3428 ( .INP(n3569), .ZN(n3671) );
  XOR2X1 U3429 ( .IN1(n3621), .IN2(n3672), .Q(n3668) );
  INVX0 U3430 ( .INP(n3339), .ZN(n3336) );
  NAND2X0 U3431 ( .IN1(n3673), .IN2(n3618), .QN(n3339) );
  NAND2X0 U3432 ( .IN1(n3623), .IN2(n3611), .QN(n3618) );
  INVX0 U3433 ( .INP(n3340), .ZN(n3660) );
  MUX21X1 U3434 ( .IN1(n3674), .IN2(n3675), .S(n3676), .Q(n3340) );
  NOR2X0 U3435 ( .IN1(n3342), .IN2(n3341), .QN(\i_m4stg_frac/a1cout[6] ) );
  XOR3X1 U3436 ( .IN1(n3574), .IN2(n3576), .IN3(n3575), .Q(n3341) );
  XOR3X1 U3437 ( .IN1(n3598), .IN2(n3596), .IN3(n3595), .Q(n3575) );
  NAND2X0 U3438 ( .IN1(n3677), .IN2(n3678), .QN(n3595) );
  MUX21X1 U3439 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1470 ), .Q(n3678) );
  MUX21X1 U3440 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1471 ), .Q(n3677) );
  NAND2X0 U3441 ( .IN1(n3679), .IN2(n3680), .QN(n3596) );
  MUX21X1 U3442 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1472 ), .Q(n3680) );
  MUX21X1 U3443 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1473 ), .Q(n3679) );
  NAND2X0 U3444 ( .IN1(n3681), .IN2(n3682), .QN(n3598) );
  MUX21X1 U3445 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1468 ), .Q(n3682) );
  MUX21X1 U3446 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1469 ), .Q(n3681) );
  AO22X1 U3447 ( .IN1(n3683), .IN2(n3684), .IN3(n3685), .IN4(n3686), .Q(n3576)
         );
  OR2X1 U3448 ( .IN1(n3684), .IN2(n3683), .Q(n3685) );
  NAND2X0 U3449 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(n3606), .QN(n3574) );
  AOI22X1 U3450 ( .IN1(n3687), .IN2(n3688), .IN3(n3689), .IN4(n3690), .QN(
        n3342) );
  NAND2X0 U3451 ( .IN1(n3691), .IN2(n3591), .QN(n3690) );
  AO22X1 U3452 ( .IN1(n3344), .IN2(n3345), .IN3(n3692), .IN4(n3343), .Q(
        \i_m4stg_frac/a1cout[69] ) );
  AO22X1 U3453 ( .IN1(n3637), .IN2(n3673), .IN3(n3693), .IN4(n3694), .Q(n3343)
         );
  AOI21X1 U3454 ( .IN1(n3623), .IN2(n3672), .IN3(n3695), .QN(n3693) );
  OR2X1 U3455 ( .IN1(n3345), .IN2(n3344), .Q(n3692) );
  INVX0 U3456 ( .INP(n3696), .ZN(n3345) );
  MUX21X1 U3457 ( .IN1(n3697), .IN2(n3698), .S(n3699), .Q(n3696) );
  XOR2X1 U3458 ( .IN1(n3676), .IN2(n3674), .Q(n3344) );
  AOI22X1 U3459 ( .IN1(n3700), .IN2(n3667), .IN3(n3663), .IN4(n3701), .QN(
        n3674) );
  OR2X1 U3460 ( .IN1(n3667), .IN2(n3700), .Q(n3701) );
  XOR3X1 U3461 ( .IN1(n3672), .IN2(n3628), .IN3(n3675), .Q(n3676) );
  XOR2X1 U3462 ( .IN1(n3702), .IN2(n3665), .Q(n3675) );
  NOR2X0 U3463 ( .IN1(n3637), .IN2(n3621), .QN(n3628) );
  INVX0 U3464 ( .INP(n3611), .ZN(n3621) );
  NAND2X0 U3465 ( .IN1(n3694), .IN2(n3608), .QN(n3611) );
  INVX0 U3466 ( .INP(n3313), .ZN(n3608) );
  AO22X1 U3467 ( .IN1(n3703), .IN2(n3704), .IN3(n3705), .IN4(n3347), .Q(
        \i_m4stg_frac/a1cout[68] ) );
  AO22X1 U3468 ( .IN1(n3706), .IN2(n3673), .IN3(n3707), .IN4(n3694), .Q(n3347)
         );
  OA21X1 U3469 ( .IN1(n3706), .IN2(n3673), .IN3(n3708), .Q(n3707) );
  NAND2X0 U3470 ( .IN1(n3348), .IN2(n3346), .QN(n3705) );
  INVX0 U3471 ( .INP(n3703), .ZN(n3346) );
  INVX0 U3472 ( .INP(n3348), .ZN(n3704) );
  MUX21X1 U3473 ( .IN1(n3709), .IN2(n3710), .S(n3711), .Q(n3348) );
  INVX0 U3474 ( .INP(n3712), .ZN(n3711) );
  XNOR2X1 U3475 ( .IN1(n3699), .IN2(n3698), .Q(n3703) );
  OA22X1 U3476 ( .IN1(n3713), .IN2(n3714), .IN3(n3666), .IN4(n3715), .Q(n3698)
         );
  AND2X1 U3477 ( .IN1(n3714), .IN2(n3713), .Q(n3715) );
  INVX0 U3478 ( .INP(n3716), .ZN(n3714) );
  XOR3X1 U3479 ( .IN1(n3623), .IN2(n3697), .IN3(n3717), .Q(n3699) );
  XOR2X1 U3480 ( .IN1(n3673), .IN2(n3718), .Q(n3717) );
  NOR2X0 U3481 ( .IN1(n3695), .IN2(n3719), .QN(n3718) );
  XNOR2X1 U3482 ( .IN1(n3702), .IN2(n3700), .Q(n3697) );
  NOR2X0 U3483 ( .IN1(n3720), .IN2(n3721), .QN(n3700) );
  XOR2X1 U3484 ( .IN1(n3666), .IN2(n3662), .Q(n3702) );
  INVX0 U3485 ( .INP(n3667), .ZN(n3662) );
  NAND2X0 U3486 ( .IN1(n3722), .IN2(n3723), .QN(n3667) );
  MUX21X1 U3487 ( .IN1(n3724), .IN2(n937), .S(\i_m4stg_frac/n671 ), .Q(n3722)
         );
  NAND2X0 U3488 ( .IN1(\i_m4stg_frac/n1530 ), .IN2(n937), .QN(n3724) );
  INVX0 U3489 ( .INP(n3637), .ZN(n3623) );
  XNOR2X1 U3490 ( .IN1(n3313), .IN2(n3694), .Q(n3637) );
  AO22X1 U3491 ( .IN1(n3725), .IN2(n3726), .IN3(n3727), .IN4(n3350), .Q(
        \i_m4stg_frac/a1cout[67] ) );
  AO22X1 U3492 ( .IN1(n3728), .IN2(n3673), .IN3(n3729), .IN4(n3730), .Q(n3350)
         );
  OR2X1 U3493 ( .IN1(n3673), .IN2(n3728), .Q(n3730) );
  NAND2X0 U3494 ( .IN1(n3351), .IN2(n3349), .QN(n3727) );
  INVX0 U3495 ( .INP(n3725), .ZN(n3349) );
  INVX0 U3496 ( .INP(n3351), .ZN(n3726) );
  MUX21X1 U3497 ( .IN1(n3731), .IN2(n3732), .S(n3733), .Q(n3351) );
  INVX0 U3498 ( .INP(n3734), .ZN(n3733) );
  XOR2X1 U3499 ( .IN1(n3712), .IN2(n3710), .Q(n3725) );
  OA22X1 U3500 ( .IN1(n3735), .IN2(n3736), .IN3(n3666), .IN4(n3737), .Q(n3710)
         );
  AND2X1 U3501 ( .IN1(n3736), .IN2(n3735), .Q(n3737) );
  XOR3X1 U3502 ( .IN1(n3673), .IN2(n3738), .IN3(n3739), .Q(n3712) );
  XNOR2X1 U3503 ( .IN1(n3709), .IN2(n3706), .Q(n3739) );
  XNOR2X1 U3504 ( .IN1(n3694), .IN2(n3695), .Q(n3706) );
  OA21X1 U3505 ( .IN1(n1123), .IN2(n3313), .IN3(n3740), .Q(n3695) );
  MUX21X1 U3506 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1519 ), .Q(n3740) );
  NAND2X0 U3507 ( .IN1(n3743), .IN2(n938), .QN(n3313) );
  XOR2X1 U3508 ( .IN1(\i_m4stg_frac/n654 ), .IN2(n907), .Q(n3743) );
  XOR3X1 U3509 ( .IN1(n3713), .IN2(n3663), .IN3(n3716), .Q(n3709) );
  XNOR2X1 U3510 ( .IN1(n3721), .IN2(n3720), .Q(n3713) );
  NAND2X0 U3511 ( .IN1(n3694), .IN2(n3708), .QN(n3738) );
  AO22X1 U3512 ( .IN1(n3744), .IN2(n3745), .IN3(n3746), .IN4(n3353), .Q(
        \i_m4stg_frac/a1cout[66] ) );
  AO22X1 U3513 ( .IN1(n3747), .IN2(n3673), .IN3(n3748), .IN4(n3749), .Q(n3353)
         );
  OR2X1 U3514 ( .IN1(n3747), .IN2(n3673), .Q(n3749) );
  NAND2X0 U3515 ( .IN1(n3354), .IN2(n3352), .QN(n3746) );
  INVX0 U3516 ( .INP(n3744), .ZN(n3352) );
  INVX0 U3517 ( .INP(n3745), .ZN(n3354) );
  MUX21X1 U3518 ( .IN1(n3750), .IN2(n3751), .S(n3752), .Q(n3745) );
  XOR2X1 U3519 ( .IN1(n3734), .IN2(n3732), .Q(n3744) );
  AOI22X1 U3520 ( .IN1(n3753), .IN2(n3754), .IN3(n3663), .IN4(n3755), .QN(
        n3732) );
  OR2X1 U3521 ( .IN1(n3754), .IN2(n3753), .Q(n3755) );
  XOR3X1 U3522 ( .IN1(n3672), .IN2(n3729), .IN3(n3756), .Q(n3734) );
  XNOR2X1 U3523 ( .IN1(n3731), .IN2(n3728), .Q(n3756) );
  XOR2X1 U3524 ( .IN1(n3708), .IN2(n3694), .Q(n3728) );
  INVX0 U3525 ( .INP(n3719), .ZN(n3694) );
  NAND2X0 U3526 ( .IN1(n3757), .IN2(n3758), .QN(n3708) );
  MUX21X1 U3527 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1518 ), .Q(n3758) );
  MUX21X1 U3528 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1519 ), .Q(n3757) );
  XOR3X1 U3529 ( .IN1(n3666), .IN2(n3735), .IN3(n3736), .Q(n3731) );
  OA221X1 U3530 ( .IN1(n3760), .IN2(\i_m4stg_frac/n674 ), .IN3(n3720), .IN4(
        n3579), .IN5(n3716), .Q(n3736) );
  NAND3X0 U3531 ( .IN1(n3720), .IN2(n3579), .IN3(n3761), .QN(n3716) );
  NAND2X0 U3532 ( .IN1(n3762), .IN2(n924), .QN(n3761) );
  OA21X1 U3533 ( .IN1(n3763), .IN2(n3506), .IN3(n3760), .Q(n3735) );
  INVX0 U3534 ( .INP(n3764), .ZN(n3763) );
  NOR2X0 U3535 ( .IN1(n3765), .IN2(n3766), .QN(n3729) );
  INVX0 U3536 ( .INP(n3673), .ZN(n3672) );
  AO22X1 U3537 ( .IN1(n3356), .IN2(n3357), .IN3(n3767), .IN4(n3355), .Q(
        \i_m4stg_frac/a1cout[65] ) );
  AO22X1 U3538 ( .IN1(n3768), .IN2(n3769), .IN3(n3770), .IN4(n3771), .Q(n3355)
         );
  OR2X1 U3539 ( .IN1(n3768), .IN2(n3769), .Q(n3771) );
  AND2X1 U3540 ( .IN1(n3772), .IN2(n3773), .Q(n3770) );
  OR2X1 U3541 ( .IN1(n3357), .IN2(n3356), .Q(n3767) );
  INVX0 U3542 ( .INP(n3774), .ZN(n3357) );
  MUX21X1 U3543 ( .IN1(n3775), .IN2(n3776), .S(n3777), .Q(n3774) );
  INVX0 U3544 ( .INP(n3778), .ZN(n3777) );
  XNOR2X1 U3545 ( .IN1(n3750), .IN2(n3752), .Q(n3356) );
  XOR3X1 U3546 ( .IN1(n3673), .IN2(n3748), .IN3(n3779), .Q(n3752) );
  XNOR2X1 U3547 ( .IN1(n3751), .IN2(n3747), .Q(n3779) );
  XOR2X1 U3548 ( .IN1(n3765), .IN2(n3766), .Q(n3747) );
  OA21X1 U3549 ( .IN1(n1313), .IN2(n3719), .IN3(n3780), .Q(n3766) );
  MUX21X1 U3550 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1519 ), .Q(n3780) );
  NAND2X0 U3551 ( .IN1(n3615), .IN2(n1133), .QN(n3719) );
  XOR2X1 U3552 ( .IN1(n1039), .IN2(\i_m4stg_frac/n1530 ), .Q(n3615) );
  AND2X1 U3553 ( .IN1(n3783), .IN2(n3784), .Q(n3765) );
  MUX21X1 U3554 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1517 ), .Q(n3784) );
  MUX21X1 U3555 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1518 ), .Q(n3783) );
  XOR3X1 U3556 ( .IN1(n3753), .IN2(n3663), .IN3(n3754), .Q(n3751) );
  AO21X1 U3557 ( .IN1(n3785), .IN2(n3764), .IN3(n3786), .Q(n3754) );
  XOR2X1 U3558 ( .IN1(n3506), .IN2(n3787), .Q(n3753) );
  NOR2X0 U3559 ( .IN1(n3788), .IN2(n3789), .QN(n3748) );
  AO21X1 U3560 ( .IN1(n3790), .IN2(n3650), .IN3(n3646), .Q(n3673) );
  INVX0 U3561 ( .INP(n3791), .ZN(n3650) );
  AO22X1 U3562 ( .IN1(n3792), .IN2(n3663), .IN3(n3793), .IN4(n3794), .Q(n3750)
         );
  NAND2X0 U3563 ( .IN1(n3666), .IN2(n3795), .QN(n3793) );
  INVX0 U3564 ( .INP(n3666), .ZN(n3663) );
  INVX0 U3565 ( .INP(n3795), .ZN(n3792) );
  AO22X1 U3566 ( .IN1(n3359), .IN2(n3360), .IN3(n3796), .IN4(n3358), .Q(
        \i_m4stg_frac/a1cout[64] ) );
  AO22X1 U3567 ( .IN1(n3797), .IN2(n3798), .IN3(n3799), .IN4(n3800), .Q(n3358)
         );
  OR2X1 U3568 ( .IN1(n3797), .IN2(n3798), .Q(n3800) );
  OR2X1 U3569 ( .IN1(n3360), .IN2(n3359), .Q(n3796) );
  INVX0 U3570 ( .INP(n3801), .ZN(n3360) );
  MUX21X1 U3571 ( .IN1(n3802), .IN2(n3803), .S(n3804), .Q(n3801) );
  INVX0 U3572 ( .INP(n3805), .ZN(n3804) );
  XNOR2X1 U3573 ( .IN1(n3778), .IN2(n3775), .Q(n3359) );
  AOI21X1 U3574 ( .IN1(n3806), .IN2(n3807), .IN3(n3808), .QN(n3775) );
  XNOR3X1 U3575 ( .IN1(n3776), .IN2(n3768), .IN3(n3809), .Q(n3778) );
  XNOR2X1 U3576 ( .IN1(n3810), .IN2(n3769), .Q(n3809) );
  AO22X1 U3577 ( .IN1(n3790), .IN2(n3649), .IN3(n3811), .IN4(n3812), .Q(n3769)
         );
  NAND2X0 U3578 ( .IN1(n3772), .IN2(n3773), .QN(n3810) );
  XOR2X1 U3579 ( .IN1(n3789), .IN2(n3788), .Q(n3768) );
  AND2X1 U3580 ( .IN1(n3813), .IN2(n3814), .Q(n3788) );
  MUX21X1 U3581 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1516 ), .Q(n3814) );
  MUX21X1 U3582 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1517 ), .Q(n3813) );
  AND2X1 U3583 ( .IN1(n3815), .IN2(n3816), .Q(n3789) );
  MUX21X1 U3584 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1519 ), .Q(n3816) );
  MUX21X1 U3585 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1518 ), .Q(n3815) );
  XNOR3X1 U3586 ( .IN1(n3794), .IN2(n3666), .IN3(n3795), .Q(n3776) );
  XOR2X1 U3587 ( .IN1(n3787), .IN2(n3785), .Q(n3795) );
  AO21X1 U3588 ( .IN1(n3819), .IN2(n3820), .IN3(n3821), .Q(n3785) );
  XOR2X1 U3589 ( .IN1(n3822), .IN2(n3657), .Q(n3666) );
  NOR2X0 U3590 ( .IN1(n3791), .IN2(n3646), .QN(n3657) );
  NOR2X0 U3591 ( .IN1(n3823), .IN2(n3629), .QN(n3646) );
  NOR2X0 U3592 ( .IN1(n3649), .IN2(n3638), .QN(n3791) );
  AO22X1 U3593 ( .IN1(n3824), .IN2(n3825), .IN3(n3826), .IN4(n3362), .Q(
        \i_m4stg_frac/a1cout[63] ) );
  AO22X1 U3594 ( .IN1(n3827), .IN2(n3828), .IN3(n3829), .IN4(n3830), .Q(n3362)
         );
  OR2X1 U3595 ( .IN1(n3827), .IN2(n3828), .Q(n3830) );
  NAND2X0 U3596 ( .IN1(n3363), .IN2(n3361), .QN(n3826) );
  INVX0 U3597 ( .INP(n3824), .ZN(n3361) );
  INVX0 U3598 ( .INP(n3363), .ZN(n3825) );
  MUX21X1 U3599 ( .IN1(n3831), .IN2(n3832), .S(n3833), .Q(n3363) );
  INVX0 U3600 ( .INP(n3834), .ZN(n3833) );
  XOR2X1 U3601 ( .IN1(n3805), .IN2(n3803), .Q(n3824) );
  AOI21X1 U3602 ( .IN1(n3835), .IN2(n3807), .IN3(n3808), .QN(n3803) );
  XNOR3X1 U3603 ( .IN1(n3798), .IN2(n3799), .IN3(n3836), .Q(n3805) );
  XNOR2X1 U3604 ( .IN1(n3802), .IN2(n3797), .Q(n3836) );
  XOR2X1 U3605 ( .IN1(n3772), .IN2(n3773), .Q(n3797) );
  NAND2X0 U3606 ( .IN1(n3837), .IN2(n3838), .QN(n3773) );
  MUX21X1 U3607 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1515 ), .Q(n3838) );
  MUX21X1 U3608 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1516 ), .Q(n3837) );
  NAND2X0 U3609 ( .IN1(n3839), .IN2(n3840), .QN(n3772) );
  MUX21X1 U3610 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1518 ), .Q(n3840) );
  MUX21X1 U3611 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1517 ), .Q(n3839) );
  XNOR2X1 U3612 ( .IN1(n3806), .IN2(n3841), .Q(n3802) );
  XOR2X1 U3613 ( .IN1(n3842), .IN2(n3811), .Q(n3806) );
  OAI21X1 U3614 ( .IN1(n3629), .IN2(n949), .IN3(n3843), .QN(n3811) );
  MUX21X1 U3615 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1519 ), .Q(n3843) );
  INVX0 U3616 ( .INP(n3638), .ZN(n3629) );
  OA21X1 U3617 ( .IN1(n907), .IN2(\i_m4stg_frac/n660 ), .IN3(n3626), .Q(n3638)
         );
  OA21X1 U3618 ( .IN1(n934), .IN2(\i_m4stg_frac/n1530 ), .IN3(n1143), .Q(n3626) );
  NOR2X0 U3619 ( .IN1(n3846), .IN2(n3847), .QN(n3799) );
  AO22X1 U3620 ( .IN1(n3790), .IN2(n3649), .IN3(n3848), .IN4(n3812), .Q(n3798)
         );
  INVX0 U3621 ( .INP(n3823), .ZN(n3649) );
  AO22X1 U3622 ( .IN1(n3849), .IN2(n3850), .IN3(n3851), .IN4(n3365), .Q(
        \i_m4stg_frac/a1cout[62] ) );
  AO22X1 U3623 ( .IN1(n3852), .IN2(n3853), .IN3(n3854), .IN4(n3855), .Q(n3365)
         );
  OR2X1 U3624 ( .IN1(n3852), .IN2(n3853), .Q(n3855) );
  NAND2X0 U3625 ( .IN1(n3366), .IN2(n3364), .QN(n3851) );
  INVX0 U3626 ( .INP(n3849), .ZN(n3364) );
  INVX0 U3627 ( .INP(n3366), .ZN(n3850) );
  MUX21X1 U3628 ( .IN1(n3856), .IN2(n3857), .S(n3858), .Q(n3366) );
  INVX0 U3629 ( .INP(n3859), .ZN(n3858) );
  XOR2X1 U3630 ( .IN1(n3834), .IN2(n3832), .Q(n3849) );
  AOI21X1 U3631 ( .IN1(n3860), .IN2(n3807), .IN3(n3808), .QN(n3832) );
  XNOR3X1 U3632 ( .IN1(n3828), .IN2(n3829), .IN3(n3861), .Q(n3834) );
  XNOR2X1 U3633 ( .IN1(n3831), .IN2(n3827), .Q(n3861) );
  XOR2X1 U3634 ( .IN1(n3847), .IN2(n3846), .Q(n3827) );
  AND2X1 U3635 ( .IN1(n3862), .IN2(n3863), .Q(n3846) );
  MUX21X1 U3636 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1514 ), .Q(n3863) );
  MUX21X1 U3637 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1515 ), .Q(n3862) );
  AND2X1 U3638 ( .IN1(n3864), .IN2(n3865), .Q(n3847) );
  MUX21X1 U3639 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1517 ), .Q(n3865) );
  MUX21X1 U3640 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1516 ), .Q(n3864) );
  XNOR2X1 U3641 ( .IN1(n3835), .IN2(n3841), .Q(n3831) );
  XOR2X1 U3642 ( .IN1(n3848), .IN2(n3842), .Q(n3835) );
  OA21X1 U3643 ( .IN1(n3822), .IN2(n3823), .IN3(n3812), .Q(n3842) );
  NAND2X0 U3644 ( .IN1(n3822), .IN2(n3823), .QN(n3812) );
  NAND2X0 U3645 ( .IN1(n3866), .IN2(n3867), .QN(n3848) );
  MUX21X1 U3646 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1518 ), .Q(n3867) );
  MUX21X1 U3647 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1519 ), .Q(n3866) );
  NOR2X0 U3648 ( .IN1(n3870), .IN2(n3871), .QN(n3829) );
  AO22X1 U3649 ( .IN1(n3872), .IN2(n3873), .IN3(n3790), .IN4(n3874), .Q(n3828)
         );
  OR2X1 U3650 ( .IN1(n3873), .IN2(n3872), .Q(n3874) );
  AO22X1 U3651 ( .IN1(n3368), .IN2(n3369), .IN3(n3875), .IN4(n3367), .Q(
        \i_m4stg_frac/a1cout[61] ) );
  AO22X1 U3652 ( .IN1(n3876), .IN2(n3877), .IN3(n3878), .IN4(n3879), .Q(n3367)
         );
  OR2X1 U3653 ( .IN1(n3876), .IN2(n3877), .Q(n3879) );
  OR2X1 U3654 ( .IN1(n3369), .IN2(n3368), .Q(n3875) );
  INVX0 U3655 ( .INP(n3880), .ZN(n3369) );
  MUX21X1 U3656 ( .IN1(n3881), .IN2(n3882), .S(n3883), .Q(n3880) );
  INVX0 U3657 ( .INP(n3884), .ZN(n3883) );
  XNOR2X1 U3658 ( .IN1(n3859), .IN2(n3856), .Q(n3368) );
  AOI21X1 U3659 ( .IN1(n3885), .IN2(n3807), .IN3(n3808), .QN(n3856) );
  XOR3X1 U3660 ( .IN1(n3886), .IN2(n3852), .IN3(n3857), .Q(n3859) );
  XNOR2X1 U3661 ( .IN1(n3860), .IN2(n3841), .Q(n3857) );
  XOR3X1 U3662 ( .IN1(n3872), .IN2(n3790), .IN3(n3873), .Q(n3860) );
  NAND2X0 U3663 ( .IN1(n3887), .IN2(n3888), .QN(n3873) );
  MUX21X1 U3664 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1517 ), .Q(n3888) );
  MUX21X1 U3665 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1518 ), .Q(n3887) );
  OAI21X1 U3666 ( .IN1(n3823), .IN2(n914), .IN3(n3889), .QN(n3872) );
  MUX21X1 U3667 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1519 ), .Q(n3889) );
  NAND2X0 U3668 ( .IN1(n3892), .IN2(n1116), .QN(n3823) );
  XOR2X1 U3669 ( .IN1(\i_m4stg_frac/n663 ), .IN2(n907), .Q(n3892) );
  XOR2X1 U3670 ( .IN1(n3871), .IN2(n3870), .Q(n3852) );
  AND2X1 U3671 ( .IN1(n3893), .IN2(n3894), .Q(n3870) );
  MUX21X1 U3672 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1513 ), .Q(n3894) );
  MUX21X1 U3673 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1514 ), .Q(n3893) );
  AND2X1 U3674 ( .IN1(n3895), .IN2(n3896), .Q(n3871) );
  MUX21X1 U3675 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1516 ), .Q(n3896) );
  MUX21X1 U3676 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1515 ), .Q(n3895) );
  XNOR2X1 U3677 ( .IN1(n3853), .IN2(n3854), .Q(n3886) );
  NOR2X0 U3678 ( .IN1(n3897), .IN2(n3898), .QN(n3854) );
  AO22X1 U3679 ( .IN1(n3790), .IN2(n3899), .IN3(n3900), .IN4(n3901), .Q(n3853)
         );
  OR2X1 U3680 ( .IN1(n3899), .IN2(n3790), .Q(n3900) );
  INVX0 U3681 ( .INP(n3822), .ZN(n3790) );
  AO22X1 U3682 ( .IN1(n3371), .IN2(n3372), .IN3(n3902), .IN4(n3370), .Q(
        \i_m4stg_frac/a1cout[60] ) );
  AO22X1 U3683 ( .IN1(n3903), .IN2(n3904), .IN3(n3905), .IN4(n3906), .Q(n3370)
         );
  OR2X1 U3684 ( .IN1(n3903), .IN2(n3904), .Q(n3906) );
  AND2X1 U3685 ( .IN1(n3907), .IN2(n3908), .Q(n3905) );
  OR2X1 U3686 ( .IN1(n3372), .IN2(n3371), .Q(n3902) );
  INVX0 U3687 ( .INP(n3909), .ZN(n3372) );
  MUX21X1 U3688 ( .IN1(n3910), .IN2(n3911), .S(n3912), .Q(n3909) );
  INVX0 U3689 ( .INP(n3913), .ZN(n3912) );
  XNOR2X1 U3690 ( .IN1(n3884), .IN2(n3881), .Q(n3371) );
  AOI21X1 U3691 ( .IN1(n3914), .IN2(n3807), .IN3(n3808), .QN(n3881) );
  INVX0 U3692 ( .INP(n3915), .ZN(n3807) );
  XOR3X1 U3693 ( .IN1(n3916), .IN2(n3876), .IN3(n3882), .Q(n3884) );
  XNOR2X1 U3694 ( .IN1(n3885), .IN2(n3841), .Q(n3882) );
  XNOR3X1 U3695 ( .IN1(n3901), .IN2(n3899), .IN3(n3822), .Q(n3885) );
  NAND2X0 U3696 ( .IN1(n3669), .IN2(n1168), .QN(n3822) );
  NAND2X0 U3697 ( .IN1(n3917), .IN2(n3918), .QN(n3899) );
  MUX21X1 U3698 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1518 ), .Q(n3918) );
  MUX21X1 U3699 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1519 ), .Q(n3917) );
  NAND2X0 U3700 ( .IN1(n3919), .IN2(n3920), .QN(n3901) );
  MUX21X1 U3701 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1516 ), .Q(n3920) );
  MUX21X1 U3702 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1517 ), .Q(n3919) );
  XOR2X1 U3703 ( .IN1(n3898), .IN2(n3897), .Q(n3876) );
  AND2X1 U3704 ( .IN1(n3921), .IN2(n3922), .Q(n3897) );
  MUX21X1 U3705 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1512 ), .Q(n3922) );
  MUX21X1 U3706 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1513 ), .Q(n3921) );
  AND2X1 U3707 ( .IN1(n3923), .IN2(n3924), .Q(n3898) );
  MUX21X1 U3708 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1515 ), .Q(n3924) );
  MUX21X1 U3709 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1514 ), .Q(n3923) );
  XNOR2X1 U3710 ( .IN1(n3877), .IN2(n3878), .Q(n3916) );
  NOR2X0 U3711 ( .IN1(n3925), .IN2(n3926), .QN(n3878) );
  AO22X1 U3712 ( .IN1(n3927), .IN2(n3928), .IN3(n3929), .IN4(n3930), .Q(n3877)
         );
  OR2X1 U3713 ( .IN1(n3927), .IN2(n3928), .Q(n3929) );
  NOR2X0 U3714 ( .IN1(n3374), .IN2(n3373), .QN(\i_m4stg_frac/a1cout[5] ) );
  XOR3X1 U3715 ( .IN1(n3687), .IN2(n3691), .IN3(n3689), .Q(n3373) );
  XOR3X1 U3716 ( .IN1(n3686), .IN2(n3684), .IN3(n3683), .Q(n3689) );
  NAND2X0 U3717 ( .IN1(n3931), .IN2(n3932), .QN(n3683) );
  MUX21X1 U3718 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1469 ), .Q(n3932) );
  MUX21X1 U3719 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1470 ), .Q(n3931) );
  NAND2X0 U3720 ( .IN1(n3933), .IN2(n3934), .QN(n3684) );
  MUX21X1 U3721 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1472 ), .Q(n3934) );
  MUX21X1 U3722 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1471 ), .Q(n3933) );
  NAND2X0 U3723 ( .IN1(n3935), .IN2(n3936), .QN(n3686) );
  MUX21X1 U3724 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1467 ), .Q(n3936) );
  MUX21X1 U3725 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1468 ), .Q(n3935) );
  INVX0 U3726 ( .INP(n3688), .ZN(n3691) );
  AO22X1 U3727 ( .IN1(n3937), .IN2(n3938), .IN3(n3939), .IN4(n3940), .Q(n3688)
         );
  OR2X1 U3728 ( .IN1(n3938), .IN2(n3937), .Q(n3939) );
  INVX0 U3729 ( .INP(n3941), .ZN(n3937) );
  AOI22X1 U3730 ( .IN1(n3942), .IN2(n3943), .IN3(n3944), .IN4(n3945), .QN(
        n3374) );
  NAND2X0 U3731 ( .IN1(n3946), .IN2(n3593), .QN(n3945) );
  AO22X1 U3732 ( .IN1(n3947), .IN2(n3948), .IN3(n3949), .IN4(n3376), .Q(
        \i_m4stg_frac/a1cout[59] ) );
  AO22X1 U3733 ( .IN1(n3950), .IN2(n3951), .IN3(n3952), .IN4(n3953), .Q(n3376)
         );
  OR2X1 U3734 ( .IN1(n3950), .IN2(n3951), .Q(n3953) );
  AND2X1 U3735 ( .IN1(n3954), .IN2(n3955), .Q(n3952) );
  NAND2X0 U3736 ( .IN1(n3377), .IN2(n3375), .QN(n3949) );
  INVX0 U3737 ( .INP(n3947), .ZN(n3375) );
  INVX0 U3738 ( .INP(n3377), .ZN(n3948) );
  MUX21X1 U3739 ( .IN1(n3956), .IN2(n3957), .S(n3958), .Q(n3377) );
  INVX0 U3740 ( .INP(n3959), .ZN(n3958) );
  XOR2X1 U3741 ( .IN1(n3913), .IN2(n3911), .Q(n3947) );
  AOI22X1 U3742 ( .IN1(n3960), .IN2(n3961), .IN3(n3962), .IN4(n3963), .QN(
        n3911) );
  OR2X1 U3743 ( .IN1(n3961), .IN2(n3960), .Q(n3963) );
  XNOR3X1 U3744 ( .IN1(n3964), .IN2(n3903), .IN3(n3910), .Q(n3913) );
  XNOR2X1 U3745 ( .IN1(n3914), .IN2(n3841), .Q(n3910) );
  NOR2X0 U3746 ( .IN1(n3915), .IN2(n3808), .QN(n3841) );
  AND2X1 U3747 ( .IN1(n3960), .IN2(n3794), .Q(n3808) );
  NOR2X0 U3748 ( .IN1(n3794), .IN2(n3960), .QN(n3915) );
  AO21X1 U3749 ( .IN1(n3965), .IN2(n3764), .IN3(n3786), .Q(n3794) );
  XOR3X1 U3750 ( .IN1(n3930), .IN2(n3928), .IN3(n3927), .Q(n3914) );
  NAND2X0 U3751 ( .IN1(n3966), .IN2(n3967), .QN(n3927) );
  MUX21X1 U3752 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1518 ), .Q(n3967) );
  MUX21X1 U3753 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1517 ), .Q(n3966) );
  AO21X1 U3754 ( .IN1(n3669), .IN2(n3606), .IN3(n3968), .Q(n3928) );
  INVX0 U3755 ( .INP(n3969), .ZN(n3968) );
  MUX21X1 U3756 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1519 ), .Q(n3969) );
  XOR2X1 U3757 ( .IN1(n912), .IN2(\i_m4stg_frac/n1530 ), .Q(n3669) );
  NAND2X0 U3758 ( .IN1(n3970), .IN2(n3971), .QN(n3930) );
  MUX21X1 U3759 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1515 ), .Q(n3971) );
  MUX21X1 U3760 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1516 ), .Q(n3970) );
  XOR2X1 U3761 ( .IN1(n3926), .IN2(n3925), .Q(n3903) );
  AND2X1 U3762 ( .IN1(n3972), .IN2(n3973), .Q(n3925) );
  MUX21X1 U3763 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1511 ), .Q(n3973) );
  MUX21X1 U3764 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1512 ), .Q(n3972) );
  AND2X1 U3765 ( .IN1(n3974), .IN2(n3975), .Q(n3926) );
  MUX21X1 U3766 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1514 ), .Q(n3975) );
  MUX21X1 U3767 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1513 ), .Q(n3974) );
  XOR2X1 U3768 ( .IN1(n3904), .IN2(n3976), .Q(n3964) );
  NAND2X0 U3769 ( .IN1(n3907), .IN2(n3908), .QN(n3976) );
  AO22X1 U3770 ( .IN1(n3977), .IN2(n3978), .IN3(n3979), .IN4(n3980), .Q(n3904)
         );
  OR2X1 U3771 ( .IN1(n3978), .IN2(n3977), .Q(n3979) );
  AO22X1 U3772 ( .IN1(n3379), .IN2(n3380), .IN3(n3981), .IN4(n3378), .Q(
        \i_m4stg_frac/a1cout[58] ) );
  AO22X1 U3773 ( .IN1(n3982), .IN2(n3983), .IN3(n3984), .IN4(n3985), .Q(n3378)
         );
  OR2X1 U3774 ( .IN1(n3982), .IN2(n3983), .Q(n3985) );
  AND2X1 U3775 ( .IN1(n3986), .IN2(n3987), .Q(n3984) );
  OR2X1 U3776 ( .IN1(n3380), .IN2(n3379), .Q(n3981) );
  INVX0 U3777 ( .INP(n3988), .ZN(n3380) );
  MUX21X1 U3778 ( .IN1(n3989), .IN2(n3990), .S(n3991), .Q(n3988) );
  INVX0 U3779 ( .INP(n3992), .ZN(n3991) );
  XNOR2X1 U3780 ( .IN1(n3959), .IN2(n3956), .Q(n3379) );
  AOI22X1 U3781 ( .IN1(n3993), .IN2(n3994), .IN3(n3995), .IN4(n3996), .QN(
        n3956) );
  OR2X1 U3782 ( .IN1(n3994), .IN2(n3993), .Q(n3996) );
  XOR3X1 U3783 ( .IN1(n3997), .IN2(n3950), .IN3(n3957), .Q(n3959) );
  XNOR3X1 U3784 ( .IN1(n3961), .IN2(n3960), .IN3(n3962), .Q(n3957) );
  XOR3X1 U3785 ( .IN1(n3977), .IN2(n3978), .IN3(n3980), .Q(n3962) );
  NAND2X0 U3786 ( .IN1(n3998), .IN2(n3999), .QN(n3980) );
  MUX21X1 U3787 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1514 ), .Q(n3999) );
  MUX21X1 U3788 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1515 ), .Q(n3998) );
  NAND2X0 U3789 ( .IN1(n4000), .IN2(n4001), .QN(n3978) );
  MUX21X1 U3790 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1518 ), .Q(n4001) );
  MUX21X1 U3791 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1519 ), .Q(n4000) );
  NAND2X0 U3792 ( .IN1(n4002), .IN2(n4003), .QN(n3977) );
  MUX21X1 U3793 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1516 ), .Q(n4003) );
  MUX21X1 U3794 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1517 ), .Q(n4002) );
  XOR2X1 U3795 ( .IN1(n4004), .IN2(n3787), .Q(n3960) );
  NAND2X0 U3796 ( .IN1(n3764), .IN2(n3760), .QN(n3787) );
  INVX0 U3797 ( .INP(n3786), .ZN(n3760) );
  NOR2X0 U3798 ( .IN1(n4005), .IN2(n3720), .QN(n3786) );
  NAND2X0 U3799 ( .IN1(n4005), .IN2(n3720), .QN(n3764) );
  AO22X1 U3800 ( .IN1(n3965), .IN2(n3762), .IN3(n4006), .IN4(n4007), .Q(n3961)
         );
  XOR2X1 U3801 ( .IN1(n3907), .IN2(n3908), .Q(n3950) );
  NAND2X0 U3802 ( .IN1(n4008), .IN2(n4009), .QN(n3908) );
  MUX21X1 U3803 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1510 ), .Q(n4009) );
  MUX21X1 U3804 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1511 ), .Q(n4008) );
  NAND2X0 U3805 ( .IN1(n4010), .IN2(n4011), .QN(n3907) );
  MUX21X1 U3806 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1513 ), .Q(n4011) );
  MUX21X1 U3807 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1512 ), .Q(n4010) );
  XOR2X1 U3808 ( .IN1(n3951), .IN2(n4012), .Q(n3997) );
  NAND2X0 U3809 ( .IN1(n3954), .IN2(n3955), .QN(n4012) );
  AO22X1 U3810 ( .IN1(n4013), .IN2(n4014), .IN3(n4015), .IN4(n4016), .Q(n3951)
         );
  OR2X1 U3811 ( .IN1(n4013), .IN2(n4014), .Q(n4015) );
  AO22X1 U3812 ( .IN1(n4017), .IN2(n4018), .IN3(n4019), .IN4(n3382), .Q(
        \i_m4stg_frac/a1cout[57] ) );
  AO22X1 U3813 ( .IN1(n4020), .IN2(n4021), .IN3(n4022), .IN4(n4023), .Q(n3382)
         );
  OR2X1 U3814 ( .IN1(n4020), .IN2(n4021), .Q(n4023) );
  AND2X1 U3815 ( .IN1(n4024), .IN2(n4025), .Q(n4022) );
  NAND2X0 U3816 ( .IN1(n3383), .IN2(n3381), .QN(n4019) );
  INVX0 U3817 ( .INP(n4017), .ZN(n3381) );
  INVX0 U3818 ( .INP(n3383), .ZN(n4018) );
  MUX21X1 U3819 ( .IN1(n4026), .IN2(n4027), .S(n4028), .Q(n3383) );
  INVX0 U3820 ( .INP(n4029), .ZN(n4028) );
  XOR2X1 U3821 ( .IN1(n3992), .IN2(n3990), .Q(n4017) );
  AOI22X1 U3822 ( .IN1(n4030), .IN2(n4031), .IN3(n4032), .IN4(n4033), .QN(
        n3990) );
  OR2X1 U3823 ( .IN1(n4031), .IN2(n4030), .Q(n4033) );
  XNOR3X1 U3824 ( .IN1(n4034), .IN2(n3982), .IN3(n3989), .Q(n3992) );
  XNOR3X1 U3825 ( .IN1(n3994), .IN2(n3993), .IN3(n3995), .Q(n3989) );
  XOR3X1 U3826 ( .IN1(n4013), .IN2(n4014), .IN3(n4016), .Q(n3995) );
  NAND2X0 U3827 ( .IN1(n4035), .IN2(n4036), .QN(n4016) );
  MUX21X1 U3828 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1513 ), .Q(n4036) );
  MUX21X1 U3829 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1514 ), .Q(n4035) );
  NAND2X0 U3830 ( .IN1(n4037), .IN2(n4038), .QN(n4014) );
  MUX21X1 U3831 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1518 ), .Q(n4038) );
  MUX21X1 U3832 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1517 ), .Q(n4037) );
  NAND2X0 U3833 ( .IN1(n4039), .IN2(n4040), .QN(n4013) );
  MUX21X1 U3834 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1515 ), .Q(n4040) );
  MUX21X1 U3835 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1516 ), .Q(n4039) );
  XOR2X1 U3836 ( .IN1(n4041), .IN2(n4006), .Q(n3993) );
  OAI21X1 U3837 ( .IN1(n3720), .IN2(n948), .IN3(n4042), .QN(n4006) );
  MUX21X1 U3838 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1519 ), .Q(n4042) );
  OAI21X1 U3839 ( .IN1(n907), .IN2(\i_m4stg_frac/n669 ), .IN3(n3723), .QN(
        n3720) );
  OA21X1 U3840 ( .IN1(n937), .IN2(\i_m4stg_frac/n1530 ), .IN3(n1142), .Q(n3723) );
  AO22X1 U3841 ( .IN1(n3965), .IN2(n3762), .IN3(n4043), .IN4(n4007), .Q(n3994)
         );
  INVX0 U3842 ( .INP(n4005), .ZN(n3762) );
  XOR2X1 U3843 ( .IN1(n3954), .IN2(n3955), .Q(n3982) );
  NAND2X0 U3844 ( .IN1(n4044), .IN2(n4045), .QN(n3955) );
  MUX21X1 U3845 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1509 ), .Q(n4045) );
  MUX21X1 U3846 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1510 ), .Q(n4044) );
  NAND2X0 U3847 ( .IN1(n4046), .IN2(n4047), .QN(n3954) );
  MUX21X1 U3848 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1512 ), .Q(n4047) );
  MUX21X1 U3849 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1511 ), .Q(n4046) );
  XOR2X1 U3850 ( .IN1(n3983), .IN2(n4048), .Q(n4034) );
  NAND2X0 U3851 ( .IN1(n3986), .IN2(n3987), .QN(n4048) );
  AO22X1 U3852 ( .IN1(n4049), .IN2(n4050), .IN3(n4051), .IN4(n4052), .Q(n3983)
         );
  OR2X1 U3853 ( .IN1(n4050), .IN2(n4049), .Q(n4051) );
  AO22X1 U3854 ( .IN1(n3385), .IN2(n3386), .IN3(n4053), .IN4(n3384), .Q(
        \i_m4stg_frac/a1cout[56] ) );
  AO22X1 U3855 ( .IN1(n4054), .IN2(n4055), .IN3(n4056), .IN4(n4057), .Q(n3384)
         );
  OR2X1 U3856 ( .IN1(n4054), .IN2(n4055), .Q(n4057) );
  AND2X1 U3857 ( .IN1(n4058), .IN2(n4059), .Q(n4056) );
  OR2X1 U3858 ( .IN1(n3386), .IN2(n3385), .Q(n4053) );
  INVX0 U3859 ( .INP(n4060), .ZN(n3386) );
  MUX21X1 U3860 ( .IN1(n4061), .IN2(n4062), .S(n4063), .Q(n4060) );
  INVX0 U3861 ( .INP(n4064), .ZN(n4063) );
  XOR2X1 U3862 ( .IN1(n4029), .IN2(n4027), .Q(n3385) );
  AOI22X1 U3863 ( .IN1(n4065), .IN2(n4066), .IN3(n4067), .IN4(n4068), .QN(
        n4027) );
  OR2X1 U3864 ( .IN1(n4066), .IN2(n4065), .Q(n4068) );
  XNOR3X1 U3865 ( .IN1(n4069), .IN2(n4020), .IN3(n4026), .Q(n4029) );
  XNOR3X1 U3866 ( .IN1(n4031), .IN2(n4030), .IN3(n4032), .Q(n4026) );
  XOR3X1 U3867 ( .IN1(n4049), .IN2(n4050), .IN3(n4052), .Q(n4032) );
  NAND2X0 U3868 ( .IN1(n4070), .IN2(n4071), .QN(n4052) );
  MUX21X1 U3869 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1512 ), .Q(n4071) );
  MUX21X1 U3870 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1513 ), .Q(n4070) );
  NAND2X0 U3871 ( .IN1(n4072), .IN2(n4073), .QN(n4050) );
  MUX21X1 U3872 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1517 ), .Q(n4073) );
  MUX21X1 U3873 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1516 ), .Q(n4072) );
  NAND2X0 U3874 ( .IN1(n4074), .IN2(n4075), .QN(n4049) );
  MUX21X1 U3875 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1514 ), .Q(n4075) );
  MUX21X1 U3876 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1515 ), .Q(n4074) );
  XOR2X1 U3877 ( .IN1(n4043), .IN2(n4041), .Q(n4030) );
  OA21X1 U3878 ( .IN1(n4004), .IN2(n4005), .IN3(n4007), .Q(n4041) );
  NAND2X0 U3879 ( .IN1(n4004), .IN2(n4005), .QN(n4007) );
  NAND2X0 U3880 ( .IN1(n4076), .IN2(n4077), .QN(n4043) );
  MUX21X1 U3881 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1518 ), .Q(n4077) );
  MUX21X1 U3882 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1519 ), .Q(n4076) );
  AO22X1 U3883 ( .IN1(n4078), .IN2(n4079), .IN3(n3965), .IN4(n4080), .Q(n4031)
         );
  OR2X1 U3884 ( .IN1(n4079), .IN2(n4078), .Q(n4080) );
  XOR2X1 U3885 ( .IN1(n3986), .IN2(n3987), .Q(n4020) );
  NAND2X0 U3886 ( .IN1(n4081), .IN2(n4082), .QN(n3987) );
  MUX21X1 U3887 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1508 ), .Q(n4082) );
  MUX21X1 U3888 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1509 ), .Q(n4081) );
  NAND2X0 U3889 ( .IN1(n4083), .IN2(n4084), .QN(n3986) );
  MUX21X1 U3890 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1511 ), .Q(n4084) );
  MUX21X1 U3891 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1510 ), .Q(n4083) );
  XOR2X1 U3892 ( .IN1(n4021), .IN2(n4085), .Q(n4069) );
  NAND2X0 U3893 ( .IN1(n4024), .IN2(n4025), .QN(n4085) );
  AO22X1 U3894 ( .IN1(n4086), .IN2(n4087), .IN3(n4088), .IN4(n4089), .Q(n4021)
         );
  OR2X1 U3895 ( .IN1(n4087), .IN2(n4086), .Q(n4088) );
  AO22X1 U3896 ( .IN1(n3388), .IN2(n3389), .IN3(n4090), .IN4(n3387), .Q(
        \i_m4stg_frac/a1cout[55] ) );
  AO22X1 U3897 ( .IN1(n4091), .IN2(n4092), .IN3(n4093), .IN4(n4094), .Q(n3387)
         );
  OR2X1 U3898 ( .IN1(n4091), .IN2(n4092), .Q(n4094) );
  AND2X1 U3899 ( .IN1(n4095), .IN2(n4096), .Q(n4093) );
  OR2X1 U3900 ( .IN1(n3389), .IN2(n3388), .Q(n4090) );
  INVX0 U3901 ( .INP(n4097), .ZN(n3389) );
  MUX21X1 U3902 ( .IN1(n4098), .IN2(n4099), .S(n4100), .Q(n4097) );
  INVX0 U3903 ( .INP(n4101), .ZN(n4100) );
  XNOR2X1 U3904 ( .IN1(n4064), .IN2(n4061), .Q(n3388) );
  OA22X1 U3905 ( .IN1(n4102), .IN2(n4103), .IN3(n4104), .IN4(n4105), .Q(n4061)
         );
  AND2X1 U3906 ( .IN1(n4103), .IN2(n4102), .Q(n4105) );
  XOR3X1 U3907 ( .IN1(n4106), .IN2(n4054), .IN3(n4062), .Q(n4064) );
  XNOR3X1 U3908 ( .IN1(n4066), .IN2(n4065), .IN3(n4067), .Q(n4062) );
  XOR3X1 U3909 ( .IN1(n4086), .IN2(n4087), .IN3(n4089), .Q(n4067) );
  NAND2X0 U3910 ( .IN1(n4107), .IN2(n4108), .QN(n4089) );
  MUX21X1 U3911 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1511 ), .Q(n4108) );
  MUX21X1 U3912 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1512 ), .Q(n4107) );
  NAND2X0 U3913 ( .IN1(n4109), .IN2(n4110), .QN(n4087) );
  MUX21X1 U3914 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1516 ), .Q(n4110) );
  MUX21X1 U3915 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1515 ), .Q(n4109) );
  NAND2X0 U3916 ( .IN1(n4111), .IN2(n4112), .QN(n4086) );
  MUX21X1 U3917 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1513 ), .Q(n4112) );
  MUX21X1 U3918 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1514 ), .Q(n4111) );
  XOR3X1 U3919 ( .IN1(n4078), .IN2(n3965), .IN3(n4079), .Q(n4065) );
  NAND2X0 U3920 ( .IN1(n4113), .IN2(n4114), .QN(n4079) );
  MUX21X1 U3921 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1517 ), .Q(n4114) );
  MUX21X1 U3922 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1518 ), .Q(n4113) );
  OAI21X1 U3923 ( .IN1(n4005), .IN2(n924), .IN3(n4115), .QN(n4078) );
  MUX21X1 U3924 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1519 ), .Q(n4115) );
  NAND2X0 U3925 ( .IN1(n4116), .IN2(n1117), .QN(n4005) );
  XOR2X1 U3926 ( .IN1(\i_m4stg_frac/n672 ), .IN2(n907), .Q(n4116) );
  AO22X1 U3927 ( .IN1(n3965), .IN2(n4117), .IN3(n4118), .IN4(n4119), .Q(n4066)
         );
  OR2X1 U3928 ( .IN1(n4117), .IN2(n3965), .Q(n4118) );
  XOR2X1 U3929 ( .IN1(n4024), .IN2(n4025), .Q(n4054) );
  NAND2X0 U3930 ( .IN1(n4120), .IN2(n4121), .QN(n4025) );
  MUX21X1 U3931 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1507 ), .Q(n4121) );
  MUX21X1 U3932 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1508 ), .Q(n4120) );
  NAND2X0 U3933 ( .IN1(n4122), .IN2(n4123), .QN(n4024) );
  MUX21X1 U3934 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1510 ), .Q(n4123) );
  MUX21X1 U3935 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1509 ), .Q(n4122) );
  XOR2X1 U3936 ( .IN1(n4055), .IN2(n4124), .Q(n4106) );
  NAND2X0 U3937 ( .IN1(n4058), .IN2(n4059), .QN(n4124) );
  AO22X1 U3938 ( .IN1(n4125), .IN2(n4126), .IN3(n4127), .IN4(n4128), .Q(n4055)
         );
  OR2X1 U3939 ( .IN1(n4125), .IN2(n4126), .Q(n4127) );
  AO22X1 U3940 ( .IN1(n3391), .IN2(n3392), .IN3(n4129), .IN4(n3390), .Q(
        \i_m4stg_frac/a1cout[54] ) );
  AO22X1 U3941 ( .IN1(n4130), .IN2(n4131), .IN3(n4132), .IN4(n4133), .Q(n3390)
         );
  OR2X1 U3942 ( .IN1(n4130), .IN2(n4131), .Q(n4133) );
  AND2X1 U3943 ( .IN1(n4134), .IN2(n4135), .Q(n4132) );
  OR2X1 U3944 ( .IN1(n3392), .IN2(n3391), .Q(n4129) );
  INVX0 U3945 ( .INP(n4136), .ZN(n3392) );
  MUX21X1 U3946 ( .IN1(n4137), .IN2(n4138), .S(n4139), .Q(n4136) );
  INVX0 U3947 ( .INP(n4140), .ZN(n4139) );
  XNOR2X1 U3948 ( .IN1(n4101), .IN2(n4098), .Q(n3391) );
  OA22X1 U3949 ( .IN1(n4141), .IN2(n4142), .IN3(n4143), .IN4(n4144), .Q(n4098)
         );
  AND2X1 U3950 ( .IN1(n4142), .IN2(n4141), .Q(n4144) );
  XOR3X1 U3951 ( .IN1(n4145), .IN2(n4091), .IN3(n4099), .Q(n4101) );
  XOR3X1 U3952 ( .IN1(n4104), .IN2(n4103), .IN3(n4102), .Q(n4099) );
  XNOR3X1 U3953 ( .IN1(n4119), .IN2(n4117), .IN3(n3965), .Q(n4102) );
  NAND2X0 U3954 ( .IN1(n4146), .IN2(n4147), .QN(n4117) );
  MUX21X1 U3955 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1518 ), .Q(n4147) );
  MUX21X1 U3956 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1519 ), .Q(n4146) );
  NAND2X0 U3957 ( .IN1(n4148), .IN2(n4149), .QN(n4119) );
  MUX21X1 U3958 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1516 ), .Q(n4149) );
  MUX21X1 U3959 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1517 ), .Q(n4148) );
  AOI22X1 U3960 ( .IN1(n4150), .IN2(n4151), .IN3(n4152), .IN4(n4153), .QN(
        n4103) );
  OR2X1 U3961 ( .IN1(n4151), .IN2(n4150), .Q(n4152) );
  XNOR3X1 U3962 ( .IN1(n4125), .IN2(n4126), .IN3(n4128), .Q(n4104) );
  NAND2X0 U3963 ( .IN1(n4154), .IN2(n4155), .QN(n4128) );
  MUX21X1 U3964 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1510 ), .Q(n4155) );
  MUX21X1 U3965 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1511 ), .Q(n4154) );
  NAND2X0 U3966 ( .IN1(n4156), .IN2(n4157), .QN(n4126) );
  MUX21X1 U3967 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1515 ), .Q(n4157) );
  MUX21X1 U3968 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1514 ), .Q(n4156) );
  NAND2X0 U3969 ( .IN1(n4158), .IN2(n4159), .QN(n4125) );
  MUX21X1 U3970 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1512 ), .Q(n4159) );
  MUX21X1 U3971 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1513 ), .Q(n4158) );
  XOR2X1 U3972 ( .IN1(n4058), .IN2(n4059), .Q(n4091) );
  NAND2X0 U3973 ( .IN1(n4160), .IN2(n4161), .QN(n4059) );
  MUX21X1 U3974 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1506 ), .Q(n4161) );
  MUX21X1 U3975 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1507 ), .Q(n4160) );
  NAND2X0 U3976 ( .IN1(n4162), .IN2(n4163), .QN(n4058) );
  MUX21X1 U3977 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1509 ), .Q(n4163) );
  MUX21X1 U3978 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1508 ), .Q(n4162) );
  XOR2X1 U3979 ( .IN1(n4092), .IN2(n4164), .Q(n4145) );
  NAND2X0 U3980 ( .IN1(n4095), .IN2(n4096), .QN(n4164) );
  AO22X1 U3981 ( .IN1(n4165), .IN2(n4166), .IN3(n4167), .IN4(n4168), .Q(n4092)
         );
  OR2X1 U3982 ( .IN1(n4165), .IN2(n4166), .Q(n4167) );
  AO22X1 U3983 ( .IN1(n4169), .IN2(n4170), .IN3(n4171), .IN4(n3394), .Q(
        \i_m4stg_frac/a1cout[53] ) );
  AO22X1 U3984 ( .IN1(n4172), .IN2(n4173), .IN3(n4174), .IN4(n4175), .Q(n3394)
         );
  OR2X1 U3985 ( .IN1(n4172), .IN2(n4173), .Q(n4175) );
  AND2X1 U3986 ( .IN1(n4176), .IN2(n4177), .Q(n4174) );
  NAND2X0 U3987 ( .IN1(n3395), .IN2(n3393), .QN(n4171) );
  INVX0 U3988 ( .INP(n4169), .ZN(n3393) );
  INVX0 U3989 ( .INP(n3395), .ZN(n4170) );
  MUX21X1 U3990 ( .IN1(n4178), .IN2(n4179), .S(n4180), .Q(n3395) );
  INVX0 U3991 ( .INP(n4181), .ZN(n4180) );
  XOR2X1 U3992 ( .IN1(n4140), .IN2(n4138), .Q(n4169) );
  OA22X1 U3993 ( .IN1(n4182), .IN2(n4183), .IN3(n4184), .IN4(n4185), .Q(n4138)
         );
  AND2X1 U3994 ( .IN1(n4183), .IN2(n4182), .Q(n4185) );
  XNOR3X1 U3995 ( .IN1(n4186), .IN2(n4130), .IN3(n4137), .Q(n4140) );
  XOR3X1 U3996 ( .IN1(n4143), .IN2(n4142), .IN3(n4141), .Q(n4137) );
  XNOR3X1 U3997 ( .IN1(n4150), .IN2(n4151), .IN3(n4153), .Q(n4141) );
  NAND2X0 U3998 ( .IN1(n4187), .IN2(n4188), .QN(n4153) );
  MUX21X1 U3999 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1515 ), .Q(n4188) );
  MUX21X1 U4000 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1516 ), .Q(n4187) );
  AO21X1 U4001 ( .IN1(n3965), .IN2(\i_m4stg_frac/n677 ), .IN3(n4189), .Q(n4151) );
  INVX0 U4002 ( .INP(n4190), .ZN(n4189) );
  MUX21X1 U4003 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1519 ), .Q(n4190) );
  INVX0 U4004 ( .INP(n4004), .ZN(n3965) );
  NAND2X0 U4005 ( .IN1(n3819), .IN2(n1134), .QN(n4004) );
  XOR2X1 U4006 ( .IN1(n1040), .IN2(\i_m4stg_frac/n1530 ), .Q(n3819) );
  NAND2X0 U4007 ( .IN1(n4191), .IN2(n4192), .QN(n4150) );
  MUX21X1 U4008 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1518 ), .Q(n4192) );
  MUX21X1 U4009 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1517 ), .Q(n4191) );
  AOI22X1 U4010 ( .IN1(n4193), .IN2(n4194), .IN3(n4195), .IN4(n4196), .QN(
        n4142) );
  OR2X1 U4011 ( .IN1(n4194), .IN2(n4193), .Q(n4195) );
  XNOR3X1 U4012 ( .IN1(n4165), .IN2(n4166), .IN3(n4168), .Q(n4143) );
  NAND2X0 U4013 ( .IN1(n4197), .IN2(n4198), .QN(n4168) );
  MUX21X1 U4014 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1509 ), .Q(n4198) );
  MUX21X1 U4015 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1510 ), .Q(n4197) );
  NAND2X0 U4016 ( .IN1(n4199), .IN2(n4200), .QN(n4166) );
  MUX21X1 U4017 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1514 ), .Q(n4200) );
  MUX21X1 U4018 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1513 ), .Q(n4199) );
  NAND2X0 U4019 ( .IN1(n4201), .IN2(n4202), .QN(n4165) );
  MUX21X1 U4020 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1511 ), .Q(n4202) );
  MUX21X1 U4021 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1512 ), .Q(n4201) );
  XOR2X1 U4022 ( .IN1(n4095), .IN2(n4096), .Q(n4130) );
  NAND2X0 U4023 ( .IN1(n4203), .IN2(n4204), .QN(n4096) );
  MUX21X1 U4024 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1505 ), .Q(n4204) );
  MUX21X1 U4025 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1506 ), .Q(n4203) );
  NAND2X0 U4026 ( .IN1(n4205), .IN2(n4206), .QN(n4095) );
  MUX21X1 U4027 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1508 ), .Q(n4206) );
  MUX21X1 U4028 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1507 ), .Q(n4205) );
  XOR2X1 U4029 ( .IN1(n4131), .IN2(n4207), .Q(n4186) );
  NAND2X0 U4030 ( .IN1(n4134), .IN2(n4135), .QN(n4207) );
  AO22X1 U4031 ( .IN1(n4208), .IN2(n4209), .IN3(n4210), .IN4(n4211), .Q(n4131)
         );
  OR2X1 U4032 ( .IN1(n4209), .IN2(n4208), .Q(n4210) );
  AO22X1 U4033 ( .IN1(n4212), .IN2(n4213), .IN3(n4214), .IN4(n3397), .Q(
        \i_m4stg_frac/a1cout[52] ) );
  AO22X1 U4034 ( .IN1(n4215), .IN2(n4216), .IN3(n4217), .IN4(n4218), .Q(n3397)
         );
  OR2X1 U4035 ( .IN1(n4215), .IN2(n4216), .Q(n4218) );
  AND2X1 U4036 ( .IN1(n4219), .IN2(n4220), .Q(n4217) );
  NAND2X0 U4037 ( .IN1(n3398), .IN2(n3396), .QN(n4214) );
  INVX0 U4038 ( .INP(n4212), .ZN(n3396) );
  INVX0 U4039 ( .INP(n3398), .ZN(n4213) );
  MUX21X1 U4040 ( .IN1(n4221), .IN2(n4222), .S(n4223), .Q(n3398) );
  INVX0 U4041 ( .INP(n4224), .ZN(n4223) );
  XOR2X1 U4042 ( .IN1(n4181), .IN2(n4179), .Q(n4212) );
  OA22X1 U4043 ( .IN1(n4225), .IN2(n4226), .IN3(n4227), .IN4(n4228), .Q(n4179)
         );
  AND2X1 U4044 ( .IN1(n4226), .IN2(n4225), .Q(n4228) );
  XNOR3X1 U4045 ( .IN1(n4229), .IN2(n4172), .IN3(n4178), .Q(n4181) );
  XOR3X1 U4046 ( .IN1(n4184), .IN2(n4183), .IN3(n4182), .Q(n4178) );
  XNOR3X1 U4047 ( .IN1(n4196), .IN2(n4194), .IN3(n4193), .Q(n4182) );
  NAND2X0 U4048 ( .IN1(n4230), .IN2(n4231), .QN(n4193) );
  MUX21X1 U4049 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1516 ), .Q(n4231) );
  MUX21X1 U4050 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1517 ), .Q(n4230) );
  NAND2X0 U4051 ( .IN1(n4232), .IN2(n4233), .QN(n4194) );
  MUX21X1 U4052 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1518 ), .Q(n4233) );
  MUX21X1 U4053 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1519 ), .Q(n4232) );
  NAND2X0 U4054 ( .IN1(n4234), .IN2(n4235), .QN(n4196) );
  MUX21X1 U4055 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1514 ), .Q(n4235) );
  MUX21X1 U4056 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1515 ), .Q(n4234) );
  AOI22X1 U4057 ( .IN1(n4236), .IN2(n4237), .IN3(n4238), .IN4(n4239), .QN(
        n4183) );
  OR2X1 U4058 ( .IN1(n4237), .IN2(n4236), .Q(n4238) );
  XNOR3X1 U4059 ( .IN1(n4208), .IN2(n4209), .IN3(n4211), .Q(n4184) );
  NAND2X0 U4060 ( .IN1(n4240), .IN2(n4241), .QN(n4211) );
  MUX21X1 U4061 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1508 ), .Q(n4241) );
  MUX21X1 U4062 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1509 ), .Q(n4240) );
  NAND2X0 U4063 ( .IN1(n4242), .IN2(n4243), .QN(n4209) );
  MUX21X1 U4064 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1513 ), .Q(n4243) );
  MUX21X1 U4065 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1512 ), .Q(n4242) );
  NAND2X0 U4066 ( .IN1(n4244), .IN2(n4245), .QN(n4208) );
  MUX21X1 U4067 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1510 ), .Q(n4245) );
  MUX21X1 U4068 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1511 ), .Q(n4244) );
  XOR2X1 U4069 ( .IN1(n4134), .IN2(n4135), .Q(n4172) );
  NAND2X0 U4070 ( .IN1(n4246), .IN2(n4247), .QN(n4135) );
  MUX21X1 U4071 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1504 ), .Q(n4247) );
  MUX21X1 U4072 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1505 ), .Q(n4246) );
  NAND2X0 U4073 ( .IN1(n4248), .IN2(n4249), .QN(n4134) );
  MUX21X1 U4074 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1507 ), .Q(n4249) );
  MUX21X1 U4075 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1506 ), .Q(n4248) );
  XOR2X1 U4076 ( .IN1(n4173), .IN2(n4250), .Q(n4229) );
  NAND2X0 U4077 ( .IN1(n4176), .IN2(n4177), .QN(n4250) );
  AO22X1 U4078 ( .IN1(n4251), .IN2(n4252), .IN3(n4253), .IN4(n4254), .Q(n4173)
         );
  OR2X1 U4079 ( .IN1(n4252), .IN2(n4251), .Q(n4253) );
  AO22X1 U4080 ( .IN1(n4255), .IN2(n4256), .IN3(n4257), .IN4(n3400), .Q(
        \i_m4stg_frac/a1cout[51] ) );
  AO22X1 U4081 ( .IN1(n4258), .IN2(n4259), .IN3(n4260), .IN4(n4261), .Q(n3400)
         );
  OR2X1 U4082 ( .IN1(n4258), .IN2(n4259), .Q(n4261) );
  AND2X1 U4083 ( .IN1(n4262), .IN2(n4263), .Q(n4260) );
  NAND2X0 U4084 ( .IN1(n3401), .IN2(n3399), .QN(n4257) );
  INVX0 U4085 ( .INP(n4255), .ZN(n3399) );
  INVX0 U4086 ( .INP(n3401), .ZN(n4256) );
  MUX21X1 U4087 ( .IN1(n4264), .IN2(n4265), .S(n4266), .Q(n3401) );
  INVX0 U4088 ( .INP(n4267), .ZN(n4266) );
  XOR2X1 U4089 ( .IN1(n4224), .IN2(n4222), .Q(n4255) );
  OA22X1 U4090 ( .IN1(n4268), .IN2(n4269), .IN3(n4270), .IN4(n4271), .Q(n4222)
         );
  AND2X1 U4091 ( .IN1(n4269), .IN2(n4268), .Q(n4271) );
  XNOR3X1 U4092 ( .IN1(n4272), .IN2(n4215), .IN3(n4221), .Q(n4224) );
  XOR3X1 U4093 ( .IN1(n4227), .IN2(n4226), .IN3(n4225), .Q(n4221) );
  XNOR3X1 U4094 ( .IN1(n4239), .IN2(n4237), .IN3(n4236), .Q(n4225) );
  NAND2X0 U4095 ( .IN1(n4273), .IN2(n4274), .QN(n4236) );
  MUX21X1 U4096 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1515 ), .Q(n4274) );
  MUX21X1 U4097 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1516 ), .Q(n4273) );
  NAND2X0 U4098 ( .IN1(n4275), .IN2(n4276), .QN(n4237) );
  MUX21X1 U4099 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1518 ), .Q(n4276) );
  MUX21X1 U4100 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1517 ), .Q(n4275) );
  NAND2X0 U4101 ( .IN1(n4277), .IN2(n4278), .QN(n4239) );
  MUX21X1 U4102 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1513 ), .Q(n4278) );
  MUX21X1 U4103 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1514 ), .Q(n4277) );
  AOI22X1 U4104 ( .IN1(n4279), .IN2(n4280), .IN3(n4281), .IN4(n4282), .QN(
        n4226) );
  OR2X1 U4105 ( .IN1(n4280), .IN2(n4279), .Q(n4281) );
  XNOR3X1 U4106 ( .IN1(n4251), .IN2(n4252), .IN3(n4254), .Q(n4227) );
  NAND2X0 U4107 ( .IN1(n4283), .IN2(n4284), .QN(n4254) );
  MUX21X1 U4108 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1507 ), .Q(n4284) );
  MUX21X1 U4109 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1508 ), .Q(n4283) );
  NAND2X0 U4110 ( .IN1(n4285), .IN2(n4286), .QN(n4252) );
  MUX21X1 U4111 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1512 ), .Q(n4286) );
  MUX21X1 U4112 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1511 ), .Q(n4285) );
  NAND2X0 U4113 ( .IN1(n4287), .IN2(n4288), .QN(n4251) );
  MUX21X1 U4114 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1509 ), .Q(n4288) );
  MUX21X1 U4115 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1510 ), .Q(n4287) );
  XOR2X1 U4116 ( .IN1(n4176), .IN2(n4177), .Q(n4215) );
  NAND2X0 U4117 ( .IN1(n4289), .IN2(n4290), .QN(n4177) );
  MUX21X1 U4118 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1503 ), .Q(n4290) );
  MUX21X1 U4119 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1504 ), .Q(n4289) );
  NAND2X0 U4120 ( .IN1(n4291), .IN2(n4292), .QN(n4176) );
  MUX21X1 U4121 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1506 ), .Q(n4292) );
  MUX21X1 U4122 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1505 ), .Q(n4291) );
  XOR2X1 U4123 ( .IN1(n4216), .IN2(n4293), .Q(n4272) );
  NAND2X0 U4124 ( .IN1(n4219), .IN2(n4220), .QN(n4293) );
  AO22X1 U4125 ( .IN1(n4294), .IN2(n4295), .IN3(n4296), .IN4(n4297), .Q(n4216)
         );
  OR2X1 U4126 ( .IN1(n4295), .IN2(n4294), .Q(n4296) );
  AO22X1 U4127 ( .IN1(n4298), .IN2(n4299), .IN3(n4300), .IN4(n3403), .Q(
        \i_m4stg_frac/a1cout[50] ) );
  AO22X1 U4128 ( .IN1(n4301), .IN2(n4302), .IN3(n4303), .IN4(n4304), .Q(n3403)
         );
  OR2X1 U4129 ( .IN1(n4301), .IN2(n4302), .Q(n4304) );
  AND2X1 U4130 ( .IN1(n4305), .IN2(n4306), .Q(n4303) );
  NAND2X0 U4131 ( .IN1(n3404), .IN2(n3402), .QN(n4300) );
  INVX0 U4132 ( .INP(n4298), .ZN(n3402) );
  INVX0 U4133 ( .INP(n3404), .ZN(n4299) );
  MUX21X1 U4134 ( .IN1(n4307), .IN2(n4308), .S(n4309), .Q(n3404) );
  INVX0 U4135 ( .INP(n4310), .ZN(n4309) );
  XOR2X1 U4136 ( .IN1(n4267), .IN2(n4265), .Q(n4298) );
  OA22X1 U4137 ( .IN1(n4311), .IN2(n4312), .IN3(n4313), .IN4(n4314), .Q(n4265)
         );
  AND2X1 U4138 ( .IN1(n4312), .IN2(n4311), .Q(n4314) );
  XNOR3X1 U4139 ( .IN1(n4315), .IN2(n4258), .IN3(n4264), .Q(n4267) );
  XOR3X1 U4140 ( .IN1(n4270), .IN2(n4269), .IN3(n4268), .Q(n4264) );
  XNOR3X1 U4141 ( .IN1(n4282), .IN2(n4280), .IN3(n4279), .Q(n4268) );
  NAND2X0 U4142 ( .IN1(n4316), .IN2(n4317), .QN(n4279) );
  MUX21X1 U4143 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1514 ), .Q(n4317) );
  MUX21X1 U4144 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1515 ), .Q(n4316) );
  NAND2X0 U4145 ( .IN1(n4318), .IN2(n4319), .QN(n4280) );
  MUX21X1 U4146 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1517 ), .Q(n4319) );
  MUX21X1 U4147 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1516 ), .Q(n4318) );
  NAND2X0 U4148 ( .IN1(n4320), .IN2(n4321), .QN(n4282) );
  MUX21X1 U4149 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1512 ), .Q(n4321) );
  MUX21X1 U4150 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1513 ), .Q(n4320) );
  AOI22X1 U4151 ( .IN1(n4322), .IN2(n4323), .IN3(n4324), .IN4(n4325), .QN(
        n4269) );
  OR2X1 U4152 ( .IN1(n4323), .IN2(n4322), .Q(n4324) );
  XNOR3X1 U4153 ( .IN1(n4294), .IN2(n4295), .IN3(n4297), .Q(n4270) );
  NAND2X0 U4154 ( .IN1(n4326), .IN2(n4327), .QN(n4297) );
  MUX21X1 U4155 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1506 ), .Q(n4327) );
  MUX21X1 U4156 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1507 ), .Q(n4326) );
  NAND2X0 U4157 ( .IN1(n4328), .IN2(n4329), .QN(n4295) );
  MUX21X1 U4158 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1511 ), .Q(n4329) );
  MUX21X1 U4159 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1510 ), .Q(n4328) );
  NAND2X0 U4160 ( .IN1(n4330), .IN2(n4331), .QN(n4294) );
  MUX21X1 U4161 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1508 ), .Q(n4331) );
  MUX21X1 U4162 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1509 ), .Q(n4330) );
  XOR2X1 U4163 ( .IN1(n4219), .IN2(n4220), .Q(n4258) );
  NAND2X0 U4164 ( .IN1(n4332), .IN2(n4333), .QN(n4220) );
  MUX21X1 U4165 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1502 ), .Q(n4333) );
  MUX21X1 U4166 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1503 ), .Q(n4332) );
  NAND2X0 U4167 ( .IN1(n4334), .IN2(n4335), .QN(n4219) );
  MUX21X1 U4168 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1505 ), .Q(n4335) );
  MUX21X1 U4169 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1504 ), .Q(n4334) );
  XOR2X1 U4170 ( .IN1(n4259), .IN2(n4336), .Q(n4315) );
  NAND2X0 U4171 ( .IN1(n4262), .IN2(n4263), .QN(n4336) );
  AO22X1 U4172 ( .IN1(n4337), .IN2(n4338), .IN3(n4339), .IN4(n4340), .Q(n4259)
         );
  OR2X1 U4173 ( .IN1(n4338), .IN2(n4337), .Q(n4339) );
  NOR2X0 U4174 ( .IN1(n3405), .IN2(n3406), .QN(\i_m4stg_frac/a1cout[4] ) );
  XNOR3X1 U4175 ( .IN1(n3593), .IN2(n3946), .IN3(n3944), .Q(n3406) );
  XNOR3X1 U4176 ( .IN1(n3940), .IN2(n3938), .IN3(n3941), .Q(n3944) );
  MUX21X1 U4177 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1467 ), .Q(n3941) );
  NAND2X0 U4178 ( .IN1(n4341), .IN2(n4342), .QN(n3938) );
  MUX21X1 U4179 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1471 ), .Q(n4342) );
  MUX21X1 U4180 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1470 ), .Q(n4341) );
  NAND2X0 U4181 ( .IN1(n4343), .IN2(n4344), .QN(n3940) );
  MUX21X1 U4182 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1468 ), .Q(n4344) );
  MUX21X1 U4183 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1469 ), .Q(n4343) );
  INVX0 U4184 ( .INP(n3943), .ZN(n3946) );
  AO22X1 U4185 ( .IN1(n4345), .IN2(n4346), .IN3(n4347), .IN4(n4348), .Q(n3943)
         );
  OR2X1 U4186 ( .IN1(n4346), .IN2(n4345), .Q(n4348) );
  INVX0 U4187 ( .INP(n3581), .ZN(n4347) );
  AOI22X1 U4188 ( .IN1(n4349), .IN2(n4350), .IN3(n4351), .IN4(n3437), .QN(
        n3405) );
  AO22X1 U4189 ( .IN1(n4352), .IN2(n4353), .IN3(n4354), .IN4(n4355), .Q(n3437)
         );
  INVX0 U4190 ( .INP(n3580), .ZN(n4355) );
  NOR2X0 U4191 ( .IN1(n4356), .IN2(n1034), .QN(n4354) );
  NAND2X0 U4192 ( .IN1(n4356), .IN2(\i_m4stg_frac/n1467 ), .QN(n4353) );
  INVX0 U4193 ( .INP(n3579), .ZN(n4352) );
  NAND2X0 U4194 ( .IN1(n3439), .IN2(n3438), .QN(n4351) );
  INVX0 U4195 ( .INP(n3439), .ZN(n4350) );
  XOR3X1 U4196 ( .IN1(n3581), .IN2(n4346), .IN3(n4345), .Q(n3439) );
  NAND2X0 U4197 ( .IN1(n4357), .IN2(n4358), .QN(n4345) );
  MUX21X1 U4198 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1470 ), .Q(n4358) );
  MUX21X1 U4199 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1469 ), .Q(n4357) );
  NAND2X0 U4200 ( .IN1(n4359), .IN2(n4360), .QN(n4346) );
  MUX21X1 U4201 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1467 ), .Q(n4360) );
  MUX21X1 U4202 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1468 ), .Q(n4359) );
  INVX0 U4203 ( .INP(n3438), .ZN(n4349) );
  NAND2X0 U4204 ( .IN1(n3470), .IN2(n3471), .QN(n3438) );
  XOR2X1 U4205 ( .IN1(n4361), .IN2(n4356), .Q(n3471) );
  AOI21X1 U4206 ( .IN1(n4362), .IN2(n3820), .IN3(n4363), .QN(n4356) );
  MUX21X1 U4207 ( .IN1(n3821), .IN2(n4364), .S(\i_m4stg_frac/n1469 ), .Q(n4363) );
  INVX0 U4208 ( .INP(n3586), .ZN(n4364) );
  INVX0 U4209 ( .INP(n3585), .ZN(n3821) );
  NAND3X0 U4210 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(n1117), .IN3(
        \i_m4stg_frac/n674 ), .QN(n4361) );
  INVX0 U4211 ( .INP(n3504), .ZN(n3470) );
  NAND3X0 U4212 ( .IN1(n3505), .IN2(n3503), .IN3(n3506), .QN(n3504) );
  NAND2X0 U4213 ( .IN1(n4365), .IN2(n4366), .QN(n3503) );
  NAND3X0 U4214 ( .IN1(\i_m4stg_frac/n677 ), .IN2(n1134), .IN3(n4362), .QN(
        n4366) );
  XOR2X1 U4215 ( .IN1(n1040), .IN2(\i_m4stg_frac/n1468 ), .Q(n4362) );
  MUX21X1 U4216 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1467 ), .Q(n4365) );
  NAND2X0 U4217 ( .IN1(\i_m4stg_frac/n677 ), .IN2(\i_m4stg_frac/n1467 ), .QN(
        n3505) );
  AO22X1 U4218 ( .IN1(n4367), .IN2(n4368), .IN3(n4369), .IN4(n3408), .Q(
        \i_m4stg_frac/a1cout[49] ) );
  AO22X1 U4219 ( .IN1(n4370), .IN2(n4371), .IN3(n4372), .IN4(n4373), .Q(n3408)
         );
  OR2X1 U4220 ( .IN1(n4370), .IN2(n4371), .Q(n4373) );
  AND2X1 U4221 ( .IN1(n4374), .IN2(n4375), .Q(n4372) );
  NAND2X0 U4222 ( .IN1(n3409), .IN2(n3407), .QN(n4369) );
  INVX0 U4223 ( .INP(n4367), .ZN(n3407) );
  INVX0 U4224 ( .INP(n3409), .ZN(n4368) );
  MUX21X1 U4225 ( .IN1(n4376), .IN2(n4377), .S(n4378), .Q(n3409) );
  INVX0 U4226 ( .INP(n4379), .ZN(n4378) );
  XOR2X1 U4227 ( .IN1(n4310), .IN2(n4308), .Q(n4367) );
  OA22X1 U4228 ( .IN1(n4380), .IN2(n4381), .IN3(n4382), .IN4(n4383), .Q(n4308)
         );
  AND2X1 U4229 ( .IN1(n4381), .IN2(n4380), .Q(n4383) );
  XNOR3X1 U4230 ( .IN1(n4384), .IN2(n4301), .IN3(n4307), .Q(n4310) );
  XOR3X1 U4231 ( .IN1(n4313), .IN2(n4312), .IN3(n4311), .Q(n4307) );
  XNOR3X1 U4232 ( .IN1(n4325), .IN2(n4323), .IN3(n4322), .Q(n4311) );
  NAND2X0 U4233 ( .IN1(n4385), .IN2(n4386), .QN(n4322) );
  MUX21X1 U4234 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1513 ), .Q(n4386) );
  MUX21X1 U4235 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1514 ), .Q(n4385) );
  NAND2X0 U4236 ( .IN1(n4387), .IN2(n4388), .QN(n4323) );
  MUX21X1 U4237 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1516 ), .Q(n4388) );
  MUX21X1 U4238 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1515 ), .Q(n4387) );
  NAND2X0 U4239 ( .IN1(n4389), .IN2(n4390), .QN(n4325) );
  MUX21X1 U4240 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1511 ), .Q(n4390) );
  MUX21X1 U4241 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1512 ), .Q(n4389) );
  AOI22X1 U4242 ( .IN1(n4391), .IN2(n4392), .IN3(n4393), .IN4(n4394), .QN(
        n4312) );
  OR2X1 U4243 ( .IN1(n4392), .IN2(n4391), .Q(n4393) );
  XNOR3X1 U4244 ( .IN1(n4337), .IN2(n4338), .IN3(n4340), .Q(n4313) );
  NAND2X0 U4245 ( .IN1(n4395), .IN2(n4396), .QN(n4340) );
  MUX21X1 U4246 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1505 ), .Q(n4396) );
  MUX21X1 U4247 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1506 ), .Q(n4395) );
  NAND2X0 U4248 ( .IN1(n4397), .IN2(n4398), .QN(n4338) );
  MUX21X1 U4249 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1510 ), .Q(n4398) );
  MUX21X1 U4250 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1509 ), .Q(n4397) );
  NAND2X0 U4251 ( .IN1(n4399), .IN2(n4400), .QN(n4337) );
  MUX21X1 U4252 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1507 ), .Q(n4400) );
  MUX21X1 U4253 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1508 ), .Q(n4399) );
  XOR2X1 U4254 ( .IN1(n4262), .IN2(n4263), .Q(n4301) );
  NAND2X0 U4255 ( .IN1(n4401), .IN2(n4402), .QN(n4263) );
  MUX21X1 U4256 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1501 ), .Q(n4402) );
  MUX21X1 U4257 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1502 ), .Q(n4401) );
  NAND2X0 U4258 ( .IN1(n4403), .IN2(n4404), .QN(n4262) );
  MUX21X1 U4259 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1504 ), .Q(n4404) );
  MUX21X1 U4260 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1503 ), .Q(n4403) );
  XOR2X1 U4261 ( .IN1(n4302), .IN2(n4405), .Q(n4384) );
  NAND2X0 U4262 ( .IN1(n4305), .IN2(n4306), .QN(n4405) );
  AO22X1 U4263 ( .IN1(n4406), .IN2(n4407), .IN3(n4408), .IN4(n4409), .Q(n4302)
         );
  OR2X1 U4264 ( .IN1(n4407), .IN2(n4406), .Q(n4408) );
  AO22X1 U4265 ( .IN1(n4410), .IN2(n4411), .IN3(n4412), .IN4(n3411), .Q(
        \i_m4stg_frac/a1cout[48] ) );
  AO22X1 U4266 ( .IN1(n4413), .IN2(n4414), .IN3(n4415), .IN4(n4416), .Q(n3411)
         );
  OR2X1 U4267 ( .IN1(n4413), .IN2(n4414), .Q(n4416) );
  AND2X1 U4268 ( .IN1(n4417), .IN2(n4418), .Q(n4415) );
  NAND2X0 U4269 ( .IN1(n3412), .IN2(n3410), .QN(n4412) );
  INVX0 U4270 ( .INP(n4410), .ZN(n3410) );
  INVX0 U4271 ( .INP(n3412), .ZN(n4411) );
  MUX21X1 U4272 ( .IN1(n4419), .IN2(n4420), .S(n4421), .Q(n3412) );
  INVX0 U4273 ( .INP(n4422), .ZN(n4421) );
  XOR2X1 U4274 ( .IN1(n4379), .IN2(n4377), .Q(n4410) );
  OA22X1 U4275 ( .IN1(n4423), .IN2(n4424), .IN3(n4425), .IN4(n4426), .Q(n4377)
         );
  AND2X1 U4276 ( .IN1(n4424), .IN2(n4423), .Q(n4426) );
  XNOR3X1 U4277 ( .IN1(n4427), .IN2(n4370), .IN3(n4376), .Q(n4379) );
  XOR3X1 U4278 ( .IN1(n4382), .IN2(n4381), .IN3(n4380), .Q(n4376) );
  XNOR3X1 U4279 ( .IN1(n4394), .IN2(n4392), .IN3(n4391), .Q(n4380) );
  NAND2X0 U4280 ( .IN1(n4428), .IN2(n4429), .QN(n4391) );
  MUX21X1 U4281 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1512 ), .Q(n4429) );
  MUX21X1 U4282 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1513 ), .Q(n4428) );
  NAND2X0 U4283 ( .IN1(n4430), .IN2(n4431), .QN(n4392) );
  MUX21X1 U4284 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1515 ), .Q(n4431) );
  MUX21X1 U4285 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1514 ), .Q(n4430) );
  NAND2X0 U4286 ( .IN1(n4432), .IN2(n4433), .QN(n4394) );
  MUX21X1 U4287 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1510 ), .Q(n4433) );
  MUX21X1 U4288 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1511 ), .Q(n4432) );
  AOI22X1 U4289 ( .IN1(n4434), .IN2(n4435), .IN3(n4436), .IN4(n4437), .QN(
        n4381) );
  OR2X1 U4290 ( .IN1(n4435), .IN2(n4434), .Q(n4436) );
  XNOR3X1 U4291 ( .IN1(n4406), .IN2(n4407), .IN3(n4409), .Q(n4382) );
  NAND2X0 U4292 ( .IN1(n4438), .IN2(n4439), .QN(n4409) );
  MUX21X1 U4293 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1504 ), .Q(n4439) );
  MUX21X1 U4294 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1505 ), .Q(n4438) );
  NAND2X0 U4295 ( .IN1(n4440), .IN2(n4441), .QN(n4407) );
  MUX21X1 U4296 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1509 ), .Q(n4441) );
  MUX21X1 U4297 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1508 ), .Q(n4440) );
  NAND2X0 U4298 ( .IN1(n4442), .IN2(n4443), .QN(n4406) );
  MUX21X1 U4299 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1506 ), .Q(n4443) );
  MUX21X1 U4300 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1507 ), .Q(n4442) );
  XOR2X1 U4301 ( .IN1(n4305), .IN2(n4306), .Q(n4370) );
  NAND2X0 U4302 ( .IN1(n4444), .IN2(n4445), .QN(n4306) );
  MUX21X1 U4303 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1500 ), .Q(n4445) );
  MUX21X1 U4304 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1501 ), .Q(n4444) );
  NAND2X0 U4305 ( .IN1(n4446), .IN2(n4447), .QN(n4305) );
  MUX21X1 U4306 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1503 ), .Q(n4447) );
  MUX21X1 U4307 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1502 ), .Q(n4446) );
  XOR2X1 U4308 ( .IN1(n4371), .IN2(n4448), .Q(n4427) );
  NAND2X0 U4309 ( .IN1(n4374), .IN2(n4375), .QN(n4448) );
  AO22X1 U4310 ( .IN1(n4449), .IN2(n4450), .IN3(n4451), .IN4(n4452), .Q(n4371)
         );
  OR2X1 U4311 ( .IN1(n4450), .IN2(n4449), .Q(n4451) );
  AO22X1 U4312 ( .IN1(n4453), .IN2(n4454), .IN3(n4455), .IN4(n3414), .Q(
        \i_m4stg_frac/a1cout[47] ) );
  AO22X1 U4313 ( .IN1(n4456), .IN2(n4457), .IN3(n4458), .IN4(n4459), .Q(n3414)
         );
  OR2X1 U4314 ( .IN1(n4456), .IN2(n4457), .Q(n4459) );
  AND2X1 U4315 ( .IN1(n4460), .IN2(n4461), .Q(n4458) );
  NAND2X0 U4316 ( .IN1(n3415), .IN2(n3413), .QN(n4455) );
  INVX0 U4317 ( .INP(n4453), .ZN(n3413) );
  INVX0 U4318 ( .INP(n3415), .ZN(n4454) );
  MUX21X1 U4319 ( .IN1(n4462), .IN2(n4463), .S(n4464), .Q(n3415) );
  INVX0 U4320 ( .INP(n4465), .ZN(n4464) );
  XOR2X1 U4321 ( .IN1(n4422), .IN2(n4420), .Q(n4453) );
  OA22X1 U4322 ( .IN1(n4466), .IN2(n4467), .IN3(n4468), .IN4(n4469), .Q(n4420)
         );
  AND2X1 U4323 ( .IN1(n4467), .IN2(n4466), .Q(n4469) );
  XNOR3X1 U4324 ( .IN1(n4470), .IN2(n4413), .IN3(n4419), .Q(n4422) );
  XOR3X1 U4325 ( .IN1(n4425), .IN2(n4424), .IN3(n4423), .Q(n4419) );
  XNOR3X1 U4326 ( .IN1(n4437), .IN2(n4435), .IN3(n4434), .Q(n4423) );
  NAND2X0 U4327 ( .IN1(n4471), .IN2(n4472), .QN(n4434) );
  MUX21X1 U4328 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1511 ), .Q(n4472) );
  MUX21X1 U4329 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1512 ), .Q(n4471) );
  NAND2X0 U4330 ( .IN1(n4473), .IN2(n4474), .QN(n4435) );
  MUX21X1 U4331 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1514 ), .Q(n4474) );
  MUX21X1 U4332 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1513 ), .Q(n4473) );
  NAND2X0 U4333 ( .IN1(n4475), .IN2(n4476), .QN(n4437) );
  MUX21X1 U4334 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1509 ), .Q(n4476) );
  MUX21X1 U4335 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1510 ), .Q(n4475) );
  AOI22X1 U4336 ( .IN1(n4477), .IN2(n4478), .IN3(n4479), .IN4(n4480), .QN(
        n4424) );
  OR2X1 U4337 ( .IN1(n4478), .IN2(n4477), .Q(n4479) );
  XNOR3X1 U4338 ( .IN1(n4449), .IN2(n4450), .IN3(n4452), .Q(n4425) );
  NAND2X0 U4339 ( .IN1(n4481), .IN2(n4482), .QN(n4452) );
  MUX21X1 U4340 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1503 ), .Q(n4482) );
  MUX21X1 U4341 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1504 ), .Q(n4481) );
  NAND2X0 U4342 ( .IN1(n4483), .IN2(n4484), .QN(n4450) );
  MUX21X1 U4343 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1508 ), .Q(n4484) );
  MUX21X1 U4344 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1507 ), .Q(n4483) );
  NAND2X0 U4345 ( .IN1(n4485), .IN2(n4486), .QN(n4449) );
  MUX21X1 U4346 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1505 ), .Q(n4486) );
  MUX21X1 U4347 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1506 ), .Q(n4485) );
  XOR2X1 U4348 ( .IN1(n4374), .IN2(n4375), .Q(n4413) );
  NAND2X0 U4349 ( .IN1(n4487), .IN2(n4488), .QN(n4375) );
  MUX21X1 U4350 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1499 ), .Q(n4488) );
  MUX21X1 U4351 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1500 ), .Q(n4487) );
  NAND2X0 U4352 ( .IN1(n4489), .IN2(n4490), .QN(n4374) );
  MUX21X1 U4353 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1502 ), .Q(n4490) );
  MUX21X1 U4354 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1501 ), .Q(n4489) );
  XOR2X1 U4355 ( .IN1(n4414), .IN2(n4491), .Q(n4470) );
  NAND2X0 U4356 ( .IN1(n4417), .IN2(n4418), .QN(n4491) );
  AO22X1 U4357 ( .IN1(n4492), .IN2(n4493), .IN3(n4494), .IN4(n4495), .Q(n4414)
         );
  OR2X1 U4358 ( .IN1(n4493), .IN2(n4492), .Q(n4494) );
  AO22X1 U4359 ( .IN1(n4496), .IN2(n4497), .IN3(n4498), .IN4(n3417), .Q(
        \i_m4stg_frac/a1cout[46] ) );
  AO22X1 U4360 ( .IN1(n4499), .IN2(n4500), .IN3(n4501), .IN4(n4502), .Q(n3417)
         );
  OR2X1 U4361 ( .IN1(n4499), .IN2(n4500), .Q(n4502) );
  AND2X1 U4362 ( .IN1(n4503), .IN2(n4504), .Q(n4501) );
  NAND2X0 U4363 ( .IN1(n3418), .IN2(n3416), .QN(n4498) );
  INVX0 U4364 ( .INP(n4496), .ZN(n3416) );
  INVX0 U4365 ( .INP(n3418), .ZN(n4497) );
  MUX21X1 U4366 ( .IN1(n4505), .IN2(n4506), .S(n4507), .Q(n3418) );
  INVX0 U4367 ( .INP(n4508), .ZN(n4507) );
  XOR2X1 U4368 ( .IN1(n4465), .IN2(n4463), .Q(n4496) );
  OA22X1 U4369 ( .IN1(n4509), .IN2(n4510), .IN3(n4511), .IN4(n4512), .Q(n4463)
         );
  AND2X1 U4370 ( .IN1(n4510), .IN2(n4509), .Q(n4512) );
  XNOR3X1 U4371 ( .IN1(n4513), .IN2(n4456), .IN3(n4462), .Q(n4465) );
  XOR3X1 U4372 ( .IN1(n4468), .IN2(n4467), .IN3(n4466), .Q(n4462) );
  XNOR3X1 U4373 ( .IN1(n4480), .IN2(n4478), .IN3(n4477), .Q(n4466) );
  NAND2X0 U4374 ( .IN1(n4514), .IN2(n4515), .QN(n4477) );
  MUX21X1 U4375 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1510 ), .Q(n4515) );
  MUX21X1 U4376 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1511 ), .Q(n4514) );
  NAND2X0 U4377 ( .IN1(n4516), .IN2(n4517), .QN(n4478) );
  MUX21X1 U4378 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1513 ), .Q(n4517) );
  MUX21X1 U4379 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1512 ), .Q(n4516) );
  NAND2X0 U4380 ( .IN1(n4518), .IN2(n4519), .QN(n4480) );
  MUX21X1 U4381 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1508 ), .Q(n4519) );
  MUX21X1 U4382 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1509 ), .Q(n4518) );
  AOI22X1 U4383 ( .IN1(n4520), .IN2(n4521), .IN3(n4522), .IN4(n4523), .QN(
        n4467) );
  OR2X1 U4384 ( .IN1(n4521), .IN2(n4520), .Q(n4522) );
  XNOR3X1 U4385 ( .IN1(n4492), .IN2(n4493), .IN3(n4495), .Q(n4468) );
  NAND2X0 U4386 ( .IN1(n4524), .IN2(n4525), .QN(n4495) );
  MUX21X1 U4387 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1502 ), .Q(n4525) );
  MUX21X1 U4388 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1503 ), .Q(n4524) );
  NAND2X0 U4389 ( .IN1(n4526), .IN2(n4527), .QN(n4493) );
  MUX21X1 U4390 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1507 ), .Q(n4527) );
  MUX21X1 U4391 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1506 ), .Q(n4526) );
  NAND2X0 U4392 ( .IN1(n4528), .IN2(n4529), .QN(n4492) );
  MUX21X1 U4393 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1504 ), .Q(n4529) );
  MUX21X1 U4394 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1505 ), .Q(n4528) );
  XOR2X1 U4395 ( .IN1(n4417), .IN2(n4418), .Q(n4456) );
  NAND2X0 U4396 ( .IN1(n4530), .IN2(n4531), .QN(n4418) );
  MUX21X1 U4397 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1498 ), .Q(n4531) );
  MUX21X1 U4398 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1499 ), .Q(n4530) );
  NAND2X0 U4399 ( .IN1(n4532), .IN2(n4533), .QN(n4417) );
  MUX21X1 U4400 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1501 ), .Q(n4533) );
  MUX21X1 U4401 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1500 ), .Q(n4532) );
  XOR2X1 U4402 ( .IN1(n4457), .IN2(n4534), .Q(n4513) );
  NAND2X0 U4403 ( .IN1(n4460), .IN2(n4461), .QN(n4534) );
  AO22X1 U4404 ( .IN1(n4535), .IN2(n4536), .IN3(n4537), .IN4(n4538), .Q(n4457)
         );
  OR2X1 U4405 ( .IN1(n4536), .IN2(n4535), .Q(n4537) );
  AO22X1 U4406 ( .IN1(n4539), .IN2(n4540), .IN3(n4541), .IN4(n3420), .Q(
        \i_m4stg_frac/a1cout[45] ) );
  AO22X1 U4407 ( .IN1(n4542), .IN2(n4543), .IN3(n4544), .IN4(n4545), .Q(n3420)
         );
  OR2X1 U4408 ( .IN1(n4542), .IN2(n4543), .Q(n4545) );
  AND2X1 U4409 ( .IN1(n4546), .IN2(n4547), .Q(n4544) );
  NAND2X0 U4410 ( .IN1(n3421), .IN2(n3419), .QN(n4541) );
  INVX0 U4411 ( .INP(n4539), .ZN(n3419) );
  INVX0 U4412 ( .INP(n3421), .ZN(n4540) );
  MUX21X1 U4413 ( .IN1(n4548), .IN2(n4549), .S(n4550), .Q(n3421) );
  INVX0 U4414 ( .INP(n4551), .ZN(n4550) );
  XOR2X1 U4415 ( .IN1(n4508), .IN2(n4506), .Q(n4539) );
  OA22X1 U4416 ( .IN1(n4552), .IN2(n4553), .IN3(n4554), .IN4(n4555), .Q(n4506)
         );
  AND2X1 U4417 ( .IN1(n4553), .IN2(n4552), .Q(n4555) );
  XNOR3X1 U4418 ( .IN1(n4556), .IN2(n4499), .IN3(n4505), .Q(n4508) );
  XOR3X1 U4419 ( .IN1(n4511), .IN2(n4510), .IN3(n4509), .Q(n4505) );
  XNOR3X1 U4420 ( .IN1(n4523), .IN2(n4521), .IN3(n4520), .Q(n4509) );
  NAND2X0 U4421 ( .IN1(n4557), .IN2(n4558), .QN(n4520) );
  MUX21X1 U4422 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1509 ), .Q(n4558) );
  MUX21X1 U4423 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1510 ), .Q(n4557) );
  NAND2X0 U4424 ( .IN1(n4559), .IN2(n4560), .QN(n4521) );
  MUX21X1 U4425 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1512 ), .Q(n4560) );
  MUX21X1 U4426 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1511 ), .Q(n4559) );
  NAND2X0 U4427 ( .IN1(n4561), .IN2(n4562), .QN(n4523) );
  MUX21X1 U4428 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1507 ), .Q(n4562) );
  MUX21X1 U4429 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1508 ), .Q(n4561) );
  AOI22X1 U4430 ( .IN1(n4563), .IN2(n4564), .IN3(n4565), .IN4(n4566), .QN(
        n4510) );
  OR2X1 U4431 ( .IN1(n4564), .IN2(n4563), .Q(n4565) );
  XNOR3X1 U4432 ( .IN1(n4535), .IN2(n4536), .IN3(n4538), .Q(n4511) );
  NAND2X0 U4433 ( .IN1(n4567), .IN2(n4568), .QN(n4538) );
  MUX21X1 U4434 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1501 ), .Q(n4568) );
  MUX21X1 U4435 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1502 ), .Q(n4567) );
  NAND2X0 U4436 ( .IN1(n4569), .IN2(n4570), .QN(n4536) );
  MUX21X1 U4437 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1506 ), .Q(n4570) );
  MUX21X1 U4438 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1505 ), .Q(n4569) );
  NAND2X0 U4439 ( .IN1(n4571), .IN2(n4572), .QN(n4535) );
  MUX21X1 U4440 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1503 ), .Q(n4572) );
  MUX21X1 U4441 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1504 ), .Q(n4571) );
  XOR2X1 U4442 ( .IN1(n4460), .IN2(n4461), .Q(n4499) );
  NAND2X0 U4443 ( .IN1(n4573), .IN2(n4574), .QN(n4461) );
  MUX21X1 U4444 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1497 ), .Q(n4574) );
  MUX21X1 U4445 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1498 ), .Q(n4573) );
  NAND2X0 U4446 ( .IN1(n4575), .IN2(n4576), .QN(n4460) );
  MUX21X1 U4447 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1500 ), .Q(n4576) );
  MUX21X1 U4448 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1499 ), .Q(n4575) );
  XOR2X1 U4449 ( .IN1(n4500), .IN2(n4577), .Q(n4556) );
  NAND2X0 U4450 ( .IN1(n4503), .IN2(n4504), .QN(n4577) );
  AO22X1 U4451 ( .IN1(n4578), .IN2(n4579), .IN3(n4580), .IN4(n4581), .Q(n4500)
         );
  OR2X1 U4452 ( .IN1(n4579), .IN2(n4578), .Q(n4580) );
  AO22X1 U4453 ( .IN1(n4582), .IN2(n4583), .IN3(n4584), .IN4(n3423), .Q(
        \i_m4stg_frac/a1cout[44] ) );
  AO22X1 U4454 ( .IN1(n4585), .IN2(n4586), .IN3(n4587), .IN4(n4588), .Q(n3423)
         );
  OR2X1 U4455 ( .IN1(n4585), .IN2(n4586), .Q(n4588) );
  AND2X1 U4456 ( .IN1(n4589), .IN2(n4590), .Q(n4587) );
  NAND2X0 U4457 ( .IN1(n3424), .IN2(n3422), .QN(n4584) );
  INVX0 U4458 ( .INP(n4582), .ZN(n3422) );
  INVX0 U4459 ( .INP(n3424), .ZN(n4583) );
  MUX21X1 U4460 ( .IN1(n4591), .IN2(n4592), .S(n4593), .Q(n3424) );
  INVX0 U4461 ( .INP(n4594), .ZN(n4593) );
  XOR2X1 U4462 ( .IN1(n4551), .IN2(n4549), .Q(n4582) );
  OA22X1 U4463 ( .IN1(n4595), .IN2(n4596), .IN3(n4597), .IN4(n4598), .Q(n4549)
         );
  AND2X1 U4464 ( .IN1(n4596), .IN2(n4595), .Q(n4598) );
  XNOR3X1 U4465 ( .IN1(n4599), .IN2(n4542), .IN3(n4548), .Q(n4551) );
  XOR3X1 U4466 ( .IN1(n4554), .IN2(n4553), .IN3(n4552), .Q(n4548) );
  XNOR3X1 U4467 ( .IN1(n4566), .IN2(n4564), .IN3(n4563), .Q(n4552) );
  NAND2X0 U4468 ( .IN1(n4600), .IN2(n4601), .QN(n4563) );
  MUX21X1 U4469 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1508 ), .Q(n4601) );
  MUX21X1 U4470 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1509 ), .Q(n4600) );
  NAND2X0 U4471 ( .IN1(n4602), .IN2(n4603), .QN(n4564) );
  MUX21X1 U4472 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1511 ), .Q(n4603) );
  MUX21X1 U4473 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1510 ), .Q(n4602) );
  NAND2X0 U4474 ( .IN1(n4604), .IN2(n4605), .QN(n4566) );
  MUX21X1 U4475 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1506 ), .Q(n4605) );
  MUX21X1 U4476 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1507 ), .Q(n4604) );
  AOI22X1 U4477 ( .IN1(n4606), .IN2(n4607), .IN3(n4608), .IN4(n4609), .QN(
        n4553) );
  OR2X1 U4478 ( .IN1(n4607), .IN2(n4606), .Q(n4608) );
  XNOR3X1 U4479 ( .IN1(n4578), .IN2(n4579), .IN3(n4581), .Q(n4554) );
  NAND2X0 U4480 ( .IN1(n4610), .IN2(n4611), .QN(n4581) );
  MUX21X1 U4481 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1500 ), .Q(n4611) );
  MUX21X1 U4482 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1501 ), .Q(n4610) );
  NAND2X0 U4483 ( .IN1(n4612), .IN2(n4613), .QN(n4579) );
  MUX21X1 U4484 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1505 ), .Q(n4613) );
  MUX21X1 U4485 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1504 ), .Q(n4612) );
  NAND2X0 U4486 ( .IN1(n4614), .IN2(n4615), .QN(n4578) );
  MUX21X1 U4487 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1502 ), .Q(n4615) );
  MUX21X1 U4488 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1503 ), .Q(n4614) );
  XOR2X1 U4489 ( .IN1(n4503), .IN2(n4504), .Q(n4542) );
  NAND2X0 U4490 ( .IN1(n4616), .IN2(n4617), .QN(n4504) );
  MUX21X1 U4491 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1496 ), .Q(n4617) );
  MUX21X1 U4492 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1497 ), .Q(n4616) );
  NAND2X0 U4493 ( .IN1(n4618), .IN2(n4619), .QN(n4503) );
  MUX21X1 U4494 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1499 ), .Q(n4619) );
  MUX21X1 U4495 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1498 ), .Q(n4618) );
  XOR2X1 U4496 ( .IN1(n4543), .IN2(n4620), .Q(n4599) );
  NAND2X0 U4497 ( .IN1(n4546), .IN2(n4547), .QN(n4620) );
  AO22X1 U4498 ( .IN1(n4621), .IN2(n4622), .IN3(n4623), .IN4(n4624), .Q(n4543)
         );
  OR2X1 U4499 ( .IN1(n4622), .IN2(n4621), .Q(n4623) );
  AO22X1 U4500 ( .IN1(n4625), .IN2(n4626), .IN3(n4627), .IN4(n3426), .Q(
        \i_m4stg_frac/a1cout[43] ) );
  AO22X1 U4501 ( .IN1(n4628), .IN2(n4629), .IN3(n4630), .IN4(n4631), .Q(n3426)
         );
  OR2X1 U4502 ( .IN1(n4628), .IN2(n4629), .Q(n4631) );
  AND2X1 U4503 ( .IN1(n4632), .IN2(n4633), .Q(n4630) );
  NAND2X0 U4504 ( .IN1(n3427), .IN2(n3425), .QN(n4627) );
  INVX0 U4505 ( .INP(n4625), .ZN(n3425) );
  INVX0 U4506 ( .INP(n3427), .ZN(n4626) );
  MUX21X1 U4507 ( .IN1(n4634), .IN2(n4635), .S(n4636), .Q(n3427) );
  INVX0 U4508 ( .INP(n4637), .ZN(n4636) );
  XOR2X1 U4509 ( .IN1(n4594), .IN2(n4592), .Q(n4625) );
  OA22X1 U4510 ( .IN1(n4638), .IN2(n4639), .IN3(n4640), .IN4(n4641), .Q(n4592)
         );
  AND2X1 U4511 ( .IN1(n4639), .IN2(n4638), .Q(n4641) );
  XNOR3X1 U4512 ( .IN1(n4642), .IN2(n4585), .IN3(n4591), .Q(n4594) );
  XOR3X1 U4513 ( .IN1(n4597), .IN2(n4596), .IN3(n4595), .Q(n4591) );
  XNOR3X1 U4514 ( .IN1(n4609), .IN2(n4607), .IN3(n4606), .Q(n4595) );
  NAND2X0 U4515 ( .IN1(n4643), .IN2(n4644), .QN(n4606) );
  MUX21X1 U4516 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1507 ), .Q(n4644) );
  MUX21X1 U4517 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1508 ), .Q(n4643) );
  NAND2X0 U4518 ( .IN1(n4645), .IN2(n4646), .QN(n4607) );
  MUX21X1 U4519 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1510 ), .Q(n4646) );
  MUX21X1 U4520 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1509 ), .Q(n4645) );
  NAND2X0 U4521 ( .IN1(n4647), .IN2(n4648), .QN(n4609) );
  MUX21X1 U4522 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1505 ), .Q(n4648) );
  MUX21X1 U4523 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1506 ), .Q(n4647) );
  AOI22X1 U4524 ( .IN1(n4649), .IN2(n4650), .IN3(n4651), .IN4(n4652), .QN(
        n4596) );
  OR2X1 U4525 ( .IN1(n4650), .IN2(n4649), .Q(n4651) );
  XNOR3X1 U4526 ( .IN1(n4621), .IN2(n4622), .IN3(n4624), .Q(n4597) );
  NAND2X0 U4527 ( .IN1(n4653), .IN2(n4654), .QN(n4624) );
  MUX21X1 U4528 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1499 ), .Q(n4654) );
  MUX21X1 U4529 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1500 ), .Q(n4653) );
  NAND2X0 U4530 ( .IN1(n4655), .IN2(n4656), .QN(n4622) );
  MUX21X1 U4531 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1504 ), .Q(n4656) );
  MUX21X1 U4532 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1503 ), .Q(n4655) );
  NAND2X0 U4533 ( .IN1(n4657), .IN2(n4658), .QN(n4621) );
  MUX21X1 U4534 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1501 ), .Q(n4658) );
  MUX21X1 U4535 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1502 ), .Q(n4657) );
  XOR2X1 U4536 ( .IN1(n4546), .IN2(n4547), .Q(n4585) );
  NAND2X0 U4537 ( .IN1(n4659), .IN2(n4660), .QN(n4547) );
  MUX21X1 U4538 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1495 ), .Q(n4660) );
  MUX21X1 U4539 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1496 ), .Q(n4659) );
  NAND2X0 U4540 ( .IN1(n4661), .IN2(n4662), .QN(n4546) );
  MUX21X1 U4541 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1498 ), .Q(n4662) );
  MUX21X1 U4542 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1497 ), .Q(n4661) );
  XOR2X1 U4543 ( .IN1(n4586), .IN2(n4663), .Q(n4642) );
  NAND2X0 U4544 ( .IN1(n4589), .IN2(n4590), .QN(n4663) );
  AO22X1 U4545 ( .IN1(n4664), .IN2(n4665), .IN3(n4666), .IN4(n4667), .Q(n4586)
         );
  OR2X1 U4546 ( .IN1(n4665), .IN2(n4664), .Q(n4666) );
  AO22X1 U4547 ( .IN1(n4668), .IN2(n4669), .IN3(n4670), .IN4(n3429), .Q(
        \i_m4stg_frac/a1cout[42] ) );
  AO22X1 U4548 ( .IN1(n4671), .IN2(n4672), .IN3(n4673), .IN4(n4674), .Q(n3429)
         );
  OR2X1 U4549 ( .IN1(n4671), .IN2(n4672), .Q(n4674) );
  AND2X1 U4550 ( .IN1(n4675), .IN2(n4676), .Q(n4673) );
  NAND2X0 U4551 ( .IN1(n3430), .IN2(n3428), .QN(n4670) );
  INVX0 U4552 ( .INP(n4668), .ZN(n3428) );
  INVX0 U4553 ( .INP(n3430), .ZN(n4669) );
  MUX21X1 U4554 ( .IN1(n4677), .IN2(n4678), .S(n4679), .Q(n3430) );
  INVX0 U4555 ( .INP(n4680), .ZN(n4679) );
  XOR2X1 U4556 ( .IN1(n4637), .IN2(n4635), .Q(n4668) );
  OA22X1 U4557 ( .IN1(n4681), .IN2(n4682), .IN3(n4683), .IN4(n4684), .Q(n4635)
         );
  AND2X1 U4558 ( .IN1(n4682), .IN2(n4681), .Q(n4684) );
  XNOR3X1 U4559 ( .IN1(n4685), .IN2(n4628), .IN3(n4634), .Q(n4637) );
  XOR3X1 U4560 ( .IN1(n4640), .IN2(n4639), .IN3(n4638), .Q(n4634) );
  XNOR3X1 U4561 ( .IN1(n4652), .IN2(n4650), .IN3(n4649), .Q(n4638) );
  NAND2X0 U4562 ( .IN1(n4686), .IN2(n4687), .QN(n4649) );
  MUX21X1 U4563 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1506 ), .Q(n4687) );
  MUX21X1 U4564 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1507 ), .Q(n4686) );
  NAND2X0 U4565 ( .IN1(n4688), .IN2(n4689), .QN(n4650) );
  MUX21X1 U4566 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1509 ), .Q(n4689) );
  MUX21X1 U4567 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1508 ), .Q(n4688) );
  NAND2X0 U4568 ( .IN1(n4690), .IN2(n4691), .QN(n4652) );
  MUX21X1 U4569 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1504 ), .Q(n4691) );
  MUX21X1 U4570 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1505 ), .Q(n4690) );
  AOI22X1 U4571 ( .IN1(n4692), .IN2(n4693), .IN3(n4694), .IN4(n4695), .QN(
        n4639) );
  OR2X1 U4572 ( .IN1(n4693), .IN2(n4692), .Q(n4694) );
  XNOR3X1 U4573 ( .IN1(n4664), .IN2(n4665), .IN3(n4667), .Q(n4640) );
  NAND2X0 U4574 ( .IN1(n4696), .IN2(n4697), .QN(n4667) );
  MUX21X1 U4575 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1498 ), .Q(n4697) );
  MUX21X1 U4576 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1499 ), .Q(n4696) );
  NAND2X0 U4577 ( .IN1(n4698), .IN2(n4699), .QN(n4665) );
  MUX21X1 U4578 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1503 ), .Q(n4699) );
  MUX21X1 U4579 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1502 ), .Q(n4698) );
  NAND2X0 U4580 ( .IN1(n4700), .IN2(n4701), .QN(n4664) );
  MUX21X1 U4581 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1500 ), .Q(n4701) );
  MUX21X1 U4582 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1501 ), .Q(n4700) );
  XOR2X1 U4583 ( .IN1(n4589), .IN2(n4590), .Q(n4628) );
  NAND2X0 U4584 ( .IN1(n4702), .IN2(n4703), .QN(n4590) );
  MUX21X1 U4585 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1494 ), .Q(n4703) );
  MUX21X1 U4586 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1495 ), .Q(n4702) );
  NAND2X0 U4587 ( .IN1(n4704), .IN2(n4705), .QN(n4589) );
  MUX21X1 U4588 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1497 ), .Q(n4705) );
  MUX21X1 U4589 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1496 ), .Q(n4704) );
  XOR2X1 U4590 ( .IN1(n4629), .IN2(n4706), .Q(n4685) );
  NAND2X0 U4591 ( .IN1(n4632), .IN2(n4633), .QN(n4706) );
  AO22X1 U4592 ( .IN1(n4707), .IN2(n4708), .IN3(n4709), .IN4(n4710), .Q(n4629)
         );
  OR2X1 U4593 ( .IN1(n4708), .IN2(n4707), .Q(n4709) );
  AO22X1 U4594 ( .IN1(n4711), .IN2(n4712), .IN3(n4713), .IN4(n3432), .Q(
        \i_m4stg_frac/a1cout[41] ) );
  AO22X1 U4595 ( .IN1(n4714), .IN2(n4715), .IN3(n4716), .IN4(n4717), .Q(n3432)
         );
  OR2X1 U4596 ( .IN1(n4714), .IN2(n4715), .Q(n4717) );
  AND2X1 U4597 ( .IN1(n4718), .IN2(n4719), .Q(n4716) );
  NAND2X0 U4598 ( .IN1(n3433), .IN2(n3431), .QN(n4713) );
  INVX0 U4599 ( .INP(n4711), .ZN(n3431) );
  INVX0 U4600 ( .INP(n3433), .ZN(n4712) );
  MUX21X1 U4601 ( .IN1(n4720), .IN2(n4721), .S(n4722), .Q(n3433) );
  INVX0 U4602 ( .INP(n4723), .ZN(n4722) );
  XOR2X1 U4603 ( .IN1(n4680), .IN2(n4678), .Q(n4711) );
  OA22X1 U4604 ( .IN1(n4724), .IN2(n4725), .IN3(n4726), .IN4(n4727), .Q(n4678)
         );
  AND2X1 U4605 ( .IN1(n4725), .IN2(n4724), .Q(n4727) );
  XNOR3X1 U4606 ( .IN1(n4728), .IN2(n4671), .IN3(n4677), .Q(n4680) );
  XOR3X1 U4607 ( .IN1(n4683), .IN2(n4682), .IN3(n4681), .Q(n4677) );
  XNOR3X1 U4608 ( .IN1(n4695), .IN2(n4693), .IN3(n4692), .Q(n4681) );
  NAND2X0 U4609 ( .IN1(n4729), .IN2(n4730), .QN(n4692) );
  MUX21X1 U4610 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1505 ), .Q(n4730) );
  MUX21X1 U4611 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1506 ), .Q(n4729) );
  NAND2X0 U4612 ( .IN1(n4731), .IN2(n4732), .QN(n4693) );
  MUX21X1 U4613 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1508 ), .Q(n4732) );
  MUX21X1 U4614 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1507 ), .Q(n4731) );
  NAND2X0 U4615 ( .IN1(n4733), .IN2(n4734), .QN(n4695) );
  MUX21X1 U4616 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1503 ), .Q(n4734) );
  MUX21X1 U4617 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1504 ), .Q(n4733) );
  AOI22X1 U4618 ( .IN1(n4735), .IN2(n4736), .IN3(n4737), .IN4(n4738), .QN(
        n4682) );
  OR2X1 U4619 ( .IN1(n4736), .IN2(n4735), .Q(n4737) );
  XNOR3X1 U4620 ( .IN1(n4707), .IN2(n4708), .IN3(n4710), .Q(n4683) );
  NAND2X0 U4621 ( .IN1(n4739), .IN2(n4740), .QN(n4710) );
  MUX21X1 U4622 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1497 ), .Q(n4740) );
  MUX21X1 U4623 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1498 ), .Q(n4739) );
  NAND2X0 U4624 ( .IN1(n4741), .IN2(n4742), .QN(n4708) );
  MUX21X1 U4625 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1502 ), .Q(n4742) );
  MUX21X1 U4626 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1501 ), .Q(n4741) );
  NAND2X0 U4627 ( .IN1(n4743), .IN2(n4744), .QN(n4707) );
  MUX21X1 U4628 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1499 ), .Q(n4744) );
  MUX21X1 U4629 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1500 ), .Q(n4743) );
  XOR2X1 U4630 ( .IN1(n4632), .IN2(n4633), .Q(n4671) );
  NAND2X0 U4631 ( .IN1(n4745), .IN2(n4746), .QN(n4633) );
  MUX21X1 U4632 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1493 ), .Q(n4746) );
  MUX21X1 U4633 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1494 ), .Q(n4745) );
  NAND2X0 U4634 ( .IN1(n4747), .IN2(n4748), .QN(n4632) );
  MUX21X1 U4635 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1496 ), .Q(n4748) );
  MUX21X1 U4636 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1495 ), .Q(n4747) );
  XOR2X1 U4637 ( .IN1(n4672), .IN2(n4749), .Q(n4728) );
  NAND2X0 U4638 ( .IN1(n4675), .IN2(n4676), .QN(n4749) );
  AO22X1 U4639 ( .IN1(n4750), .IN2(n4751), .IN3(n4752), .IN4(n4753), .Q(n4672)
         );
  OR2X1 U4640 ( .IN1(n4751), .IN2(n4750), .Q(n4752) );
  AO22X1 U4641 ( .IN1(n4754), .IN2(n4755), .IN3(n4756), .IN4(n3435), .Q(
        \i_m4stg_frac/a1cout[40] ) );
  AO22X1 U4642 ( .IN1(n4757), .IN2(n4758), .IN3(n4759), .IN4(n4760), .Q(n3435)
         );
  OR2X1 U4643 ( .IN1(n4757), .IN2(n4758), .Q(n4760) );
  AND2X1 U4644 ( .IN1(n4761), .IN2(n4762), .Q(n4759) );
  NAND2X0 U4645 ( .IN1(n3436), .IN2(n3434), .QN(n4756) );
  INVX0 U4646 ( .INP(n4754), .ZN(n3434) );
  INVX0 U4647 ( .INP(n3436), .ZN(n4755) );
  MUX21X1 U4648 ( .IN1(n4763), .IN2(n4764), .S(n4765), .Q(n3436) );
  INVX0 U4649 ( .INP(n4766), .ZN(n4765) );
  XOR2X1 U4650 ( .IN1(n4723), .IN2(n4721), .Q(n4754) );
  OA22X1 U4651 ( .IN1(n4767), .IN2(n4768), .IN3(n4769), .IN4(n4770), .Q(n4721)
         );
  AND2X1 U4652 ( .IN1(n4768), .IN2(n4767), .Q(n4770) );
  XNOR3X1 U4653 ( .IN1(n4771), .IN2(n4714), .IN3(n4720), .Q(n4723) );
  XOR3X1 U4654 ( .IN1(n4726), .IN2(n4725), .IN3(n4724), .Q(n4720) );
  XNOR3X1 U4655 ( .IN1(n4738), .IN2(n4736), .IN3(n4735), .Q(n4724) );
  NAND2X0 U4656 ( .IN1(n4772), .IN2(n4773), .QN(n4735) );
  MUX21X1 U4657 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1504 ), .Q(n4773) );
  MUX21X1 U4658 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1505 ), .Q(n4772) );
  NAND2X0 U4659 ( .IN1(n4774), .IN2(n4775), .QN(n4736) );
  MUX21X1 U4660 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1507 ), .Q(n4775) );
  MUX21X1 U4661 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1506 ), .Q(n4774) );
  NAND2X0 U4662 ( .IN1(n4776), .IN2(n4777), .QN(n4738) );
  MUX21X1 U4663 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1502 ), .Q(n4777) );
  MUX21X1 U4664 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1503 ), .Q(n4776) );
  AOI22X1 U4665 ( .IN1(n4778), .IN2(n4779), .IN3(n4780), .IN4(n4781), .QN(
        n4725) );
  OR2X1 U4666 ( .IN1(n4779), .IN2(n4778), .Q(n4780) );
  XNOR3X1 U4667 ( .IN1(n4750), .IN2(n4751), .IN3(n4753), .Q(n4726) );
  NAND2X0 U4668 ( .IN1(n4782), .IN2(n4783), .QN(n4753) );
  MUX21X1 U4669 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1496 ), .Q(n4783) );
  MUX21X1 U4670 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1497 ), .Q(n4782) );
  NAND2X0 U4671 ( .IN1(n4784), .IN2(n4785), .QN(n4751) );
  MUX21X1 U4672 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1501 ), .Q(n4785) );
  MUX21X1 U4673 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1500 ), .Q(n4784) );
  NAND2X0 U4674 ( .IN1(n4786), .IN2(n4787), .QN(n4750) );
  MUX21X1 U4675 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1498 ), .Q(n4787) );
  MUX21X1 U4676 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1499 ), .Q(n4786) );
  XOR2X1 U4677 ( .IN1(n4675), .IN2(n4676), .Q(n4714) );
  NAND2X0 U4678 ( .IN1(n4788), .IN2(n4789), .QN(n4676) );
  MUX21X1 U4679 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1492 ), .Q(n4789) );
  MUX21X1 U4680 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1493 ), .Q(n4788) );
  NAND2X0 U4681 ( .IN1(n4790), .IN2(n4791), .QN(n4675) );
  MUX21X1 U4682 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1495 ), .Q(n4791) );
  MUX21X1 U4683 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1494 ), .Q(n4790) );
  XOR2X1 U4684 ( .IN1(n4715), .IN2(n4792), .Q(n4771) );
  NAND2X0 U4685 ( .IN1(n4718), .IN2(n4719), .QN(n4792) );
  AO22X1 U4686 ( .IN1(n4793), .IN2(n4794), .IN3(n4795), .IN4(n4796), .Q(n4715)
         );
  OR2X1 U4687 ( .IN1(n4794), .IN2(n4793), .Q(n4795) );
  AO22X1 U4688 ( .IN1(n4797), .IN2(n4798), .IN3(n4799), .IN4(n3441), .Q(
        \i_m4stg_frac/a1cout[39] ) );
  AO22X1 U4689 ( .IN1(n4800), .IN2(n4801), .IN3(n4802), .IN4(n4803), .Q(n3441)
         );
  OR2X1 U4690 ( .IN1(n4800), .IN2(n4801), .Q(n4803) );
  AND2X1 U4691 ( .IN1(n4804), .IN2(n4805), .Q(n4802) );
  NAND2X0 U4692 ( .IN1(n3442), .IN2(n3440), .QN(n4799) );
  INVX0 U4693 ( .INP(n4797), .ZN(n3440) );
  INVX0 U4694 ( .INP(n3442), .ZN(n4798) );
  MUX21X1 U4695 ( .IN1(n4806), .IN2(n4807), .S(n4808), .Q(n3442) );
  INVX0 U4696 ( .INP(n4809), .ZN(n4808) );
  XOR2X1 U4697 ( .IN1(n4766), .IN2(n4764), .Q(n4797) );
  OA22X1 U4698 ( .IN1(n4810), .IN2(n4811), .IN3(n4812), .IN4(n4813), .Q(n4764)
         );
  AND2X1 U4699 ( .IN1(n4811), .IN2(n4810), .Q(n4813) );
  XNOR3X1 U4700 ( .IN1(n4814), .IN2(n4757), .IN3(n4763), .Q(n4766) );
  XOR3X1 U4701 ( .IN1(n4769), .IN2(n4768), .IN3(n4767), .Q(n4763) );
  XNOR3X1 U4702 ( .IN1(n4781), .IN2(n4779), .IN3(n4778), .Q(n4767) );
  NAND2X0 U4703 ( .IN1(n4815), .IN2(n4816), .QN(n4778) );
  MUX21X1 U4704 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1503 ), .Q(n4816) );
  MUX21X1 U4705 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1504 ), .Q(n4815) );
  NAND2X0 U4706 ( .IN1(n4817), .IN2(n4818), .QN(n4779) );
  MUX21X1 U4707 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1506 ), .Q(n4818) );
  MUX21X1 U4708 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1505 ), .Q(n4817) );
  NAND2X0 U4709 ( .IN1(n4819), .IN2(n4820), .QN(n4781) );
  MUX21X1 U4710 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1501 ), .Q(n4820) );
  MUX21X1 U4711 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1502 ), .Q(n4819) );
  AOI22X1 U4712 ( .IN1(n4821), .IN2(n4822), .IN3(n4823), .IN4(n4824), .QN(
        n4768) );
  OR2X1 U4713 ( .IN1(n4822), .IN2(n4821), .Q(n4823) );
  XNOR3X1 U4714 ( .IN1(n4793), .IN2(n4794), .IN3(n4796), .Q(n4769) );
  NAND2X0 U4715 ( .IN1(n4825), .IN2(n4826), .QN(n4796) );
  MUX21X1 U4716 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1495 ), .Q(n4826) );
  MUX21X1 U4717 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1496 ), .Q(n4825) );
  NAND2X0 U4718 ( .IN1(n4827), .IN2(n4828), .QN(n4794) );
  MUX21X1 U4719 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1500 ), .Q(n4828) );
  MUX21X1 U4720 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1499 ), .Q(n4827) );
  NAND2X0 U4721 ( .IN1(n4829), .IN2(n4830), .QN(n4793) );
  MUX21X1 U4722 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1497 ), .Q(n4830) );
  MUX21X1 U4723 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1498 ), .Q(n4829) );
  XOR2X1 U4724 ( .IN1(n4718), .IN2(n4719), .Q(n4757) );
  NAND2X0 U4725 ( .IN1(n4831), .IN2(n4832), .QN(n4719) );
  MUX21X1 U4726 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1491 ), .Q(n4832) );
  MUX21X1 U4727 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1492 ), .Q(n4831) );
  NAND2X0 U4728 ( .IN1(n4833), .IN2(n4834), .QN(n4718) );
  MUX21X1 U4729 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1494 ), .Q(n4834) );
  MUX21X1 U4730 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1493 ), .Q(n4833) );
  XOR2X1 U4731 ( .IN1(n4758), .IN2(n4835), .Q(n4814) );
  NAND2X0 U4732 ( .IN1(n4761), .IN2(n4762), .QN(n4835) );
  AO22X1 U4733 ( .IN1(n4836), .IN2(n4837), .IN3(n4838), .IN4(n4839), .Q(n4758)
         );
  OR2X1 U4734 ( .IN1(n4837), .IN2(n4836), .Q(n4838) );
  AO22X1 U4735 ( .IN1(n4840), .IN2(n4841), .IN3(n4842), .IN4(n3444), .Q(
        \i_m4stg_frac/a1cout[38] ) );
  AO22X1 U4736 ( .IN1(n4843), .IN2(n4844), .IN3(n4845), .IN4(n4846), .Q(n3444)
         );
  OR2X1 U4737 ( .IN1(n4843), .IN2(n4844), .Q(n4846) );
  AND2X1 U4738 ( .IN1(n4847), .IN2(n4848), .Q(n4845) );
  NAND2X0 U4739 ( .IN1(n3445), .IN2(n3443), .QN(n4842) );
  INVX0 U4740 ( .INP(n4840), .ZN(n3443) );
  INVX0 U4741 ( .INP(n3445), .ZN(n4841) );
  MUX21X1 U4742 ( .IN1(n4849), .IN2(n4850), .S(n4851), .Q(n3445) );
  INVX0 U4743 ( .INP(n4852), .ZN(n4851) );
  XOR2X1 U4744 ( .IN1(n4809), .IN2(n4807), .Q(n4840) );
  OA22X1 U4745 ( .IN1(n4853), .IN2(n4854), .IN3(n4855), .IN4(n4856), .Q(n4807)
         );
  AND2X1 U4746 ( .IN1(n4854), .IN2(n4853), .Q(n4856) );
  XNOR3X1 U4747 ( .IN1(n4857), .IN2(n4800), .IN3(n4806), .Q(n4809) );
  XOR3X1 U4748 ( .IN1(n4812), .IN2(n4811), .IN3(n4810), .Q(n4806) );
  XNOR3X1 U4749 ( .IN1(n4824), .IN2(n4822), .IN3(n4821), .Q(n4810) );
  NAND2X0 U4750 ( .IN1(n4858), .IN2(n4859), .QN(n4821) );
  MUX21X1 U4751 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1502 ), .Q(n4859) );
  MUX21X1 U4752 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1503 ), .Q(n4858) );
  NAND2X0 U4753 ( .IN1(n4860), .IN2(n4861), .QN(n4822) );
  MUX21X1 U4754 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1505 ), .Q(n4861) );
  MUX21X1 U4755 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1504 ), .Q(n4860) );
  NAND2X0 U4756 ( .IN1(n4862), .IN2(n4863), .QN(n4824) );
  MUX21X1 U4757 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1500 ), .Q(n4863) );
  MUX21X1 U4758 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1501 ), .Q(n4862) );
  AOI22X1 U4759 ( .IN1(n4864), .IN2(n4865), .IN3(n4866), .IN4(n4867), .QN(
        n4811) );
  OR2X1 U4760 ( .IN1(n4865), .IN2(n4864), .Q(n4866) );
  XNOR3X1 U4761 ( .IN1(n4836), .IN2(n4837), .IN3(n4839), .Q(n4812) );
  NAND2X0 U4762 ( .IN1(n4868), .IN2(n4869), .QN(n4839) );
  MUX21X1 U4763 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1494 ), .Q(n4869) );
  MUX21X1 U4764 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1495 ), .Q(n4868) );
  NAND2X0 U4765 ( .IN1(n4870), .IN2(n4871), .QN(n4837) );
  MUX21X1 U4766 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1499 ), .Q(n4871) );
  MUX21X1 U4767 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1498 ), .Q(n4870) );
  NAND2X0 U4768 ( .IN1(n4872), .IN2(n4873), .QN(n4836) );
  MUX21X1 U4769 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1496 ), .Q(n4873) );
  MUX21X1 U4770 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1497 ), .Q(n4872) );
  XOR2X1 U4771 ( .IN1(n4761), .IN2(n4762), .Q(n4800) );
  NAND2X0 U4772 ( .IN1(n4874), .IN2(n4875), .QN(n4762) );
  MUX21X1 U4773 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1490 ), .Q(n4875) );
  MUX21X1 U4774 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1491 ), .Q(n4874) );
  NAND2X0 U4775 ( .IN1(n4876), .IN2(n4877), .QN(n4761) );
  MUX21X1 U4776 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1493 ), .Q(n4877) );
  MUX21X1 U4777 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1492 ), .Q(n4876) );
  XOR2X1 U4778 ( .IN1(n4801), .IN2(n4878), .Q(n4857) );
  NAND2X0 U4779 ( .IN1(n4804), .IN2(n4805), .QN(n4878) );
  AO22X1 U4780 ( .IN1(n4879), .IN2(n4880), .IN3(n4881), .IN4(n4882), .Q(n4801)
         );
  OR2X1 U4781 ( .IN1(n4880), .IN2(n4879), .Q(n4881) );
  AO22X1 U4782 ( .IN1(n4883), .IN2(n4884), .IN3(n4885), .IN4(n3447), .Q(
        \i_m4stg_frac/a1cout[37] ) );
  AO22X1 U4783 ( .IN1(n4886), .IN2(n4887), .IN3(n4888), .IN4(n4889), .Q(n3447)
         );
  OR2X1 U4784 ( .IN1(n4886), .IN2(n4887), .Q(n4889) );
  AND2X1 U4785 ( .IN1(n4890), .IN2(n4891), .Q(n4888) );
  NAND2X0 U4786 ( .IN1(n3448), .IN2(n3446), .QN(n4885) );
  INVX0 U4787 ( .INP(n4883), .ZN(n3446) );
  INVX0 U4788 ( .INP(n3448), .ZN(n4884) );
  MUX21X1 U4789 ( .IN1(n4892), .IN2(n4893), .S(n4894), .Q(n3448) );
  INVX0 U4790 ( .INP(n4895), .ZN(n4894) );
  XOR2X1 U4791 ( .IN1(n4852), .IN2(n4850), .Q(n4883) );
  OA22X1 U4792 ( .IN1(n4896), .IN2(n4897), .IN3(n4898), .IN4(n4899), .Q(n4850)
         );
  AND2X1 U4793 ( .IN1(n4897), .IN2(n4896), .Q(n4899) );
  XNOR3X1 U4794 ( .IN1(n4900), .IN2(n4843), .IN3(n4849), .Q(n4852) );
  XOR3X1 U4795 ( .IN1(n4855), .IN2(n4854), .IN3(n4853), .Q(n4849) );
  XNOR3X1 U4796 ( .IN1(n4867), .IN2(n4865), .IN3(n4864), .Q(n4853) );
  NAND2X0 U4797 ( .IN1(n4901), .IN2(n4902), .QN(n4864) );
  MUX21X1 U4798 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1501 ), .Q(n4902) );
  MUX21X1 U4799 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1502 ), .Q(n4901) );
  NAND2X0 U4800 ( .IN1(n4903), .IN2(n4904), .QN(n4865) );
  MUX21X1 U4801 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1504 ), .Q(n4904) );
  MUX21X1 U4802 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1503 ), .Q(n4903) );
  NAND2X0 U4803 ( .IN1(n4905), .IN2(n4906), .QN(n4867) );
  MUX21X1 U4804 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1499 ), .Q(n4906) );
  MUX21X1 U4805 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1500 ), .Q(n4905) );
  AOI22X1 U4806 ( .IN1(n4907), .IN2(n4908), .IN3(n4909), .IN4(n4910), .QN(
        n4854) );
  OR2X1 U4807 ( .IN1(n4908), .IN2(n4907), .Q(n4909) );
  XNOR3X1 U4808 ( .IN1(n4879), .IN2(n4880), .IN3(n4882), .Q(n4855) );
  NAND2X0 U4809 ( .IN1(n4911), .IN2(n4912), .QN(n4882) );
  MUX21X1 U4810 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1493 ), .Q(n4912) );
  MUX21X1 U4811 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1494 ), .Q(n4911) );
  NAND2X0 U4812 ( .IN1(n4913), .IN2(n4914), .QN(n4880) );
  MUX21X1 U4813 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1498 ), .Q(n4914) );
  MUX21X1 U4814 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1497 ), .Q(n4913) );
  NAND2X0 U4815 ( .IN1(n4915), .IN2(n4916), .QN(n4879) );
  MUX21X1 U4816 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1495 ), .Q(n4916) );
  MUX21X1 U4817 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1496 ), .Q(n4915) );
  XOR2X1 U4818 ( .IN1(n4804), .IN2(n4805), .Q(n4843) );
  NAND2X0 U4819 ( .IN1(n4917), .IN2(n4918), .QN(n4805) );
  MUX21X1 U4820 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1489 ), .Q(n4918) );
  MUX21X1 U4821 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1490 ), .Q(n4917) );
  NAND2X0 U4822 ( .IN1(n4919), .IN2(n4920), .QN(n4804) );
  MUX21X1 U4823 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1492 ), .Q(n4920) );
  MUX21X1 U4824 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1491 ), .Q(n4919) );
  XOR2X1 U4825 ( .IN1(n4844), .IN2(n4921), .Q(n4900) );
  NAND2X0 U4826 ( .IN1(n4847), .IN2(n4848), .QN(n4921) );
  AO22X1 U4827 ( .IN1(n4922), .IN2(n4923), .IN3(n4924), .IN4(n4925), .Q(n4844)
         );
  OR2X1 U4828 ( .IN1(n4923), .IN2(n4922), .Q(n4924) );
  AO22X1 U4829 ( .IN1(n4926), .IN2(n4927), .IN3(n4928), .IN4(n3450), .Q(
        \i_m4stg_frac/a1cout[36] ) );
  AO22X1 U4830 ( .IN1(n4929), .IN2(n4930), .IN3(n4931), .IN4(n4932), .Q(n3450)
         );
  OR2X1 U4831 ( .IN1(n4929), .IN2(n4930), .Q(n4932) );
  AND2X1 U4832 ( .IN1(n4933), .IN2(n4934), .Q(n4931) );
  NAND2X0 U4833 ( .IN1(n3451), .IN2(n3449), .QN(n4928) );
  INVX0 U4834 ( .INP(n4926), .ZN(n3449) );
  INVX0 U4835 ( .INP(n3451), .ZN(n4927) );
  MUX21X1 U4836 ( .IN1(n4935), .IN2(n4936), .S(n4937), .Q(n3451) );
  INVX0 U4837 ( .INP(n4938), .ZN(n4937) );
  XOR2X1 U4838 ( .IN1(n4895), .IN2(n4893), .Q(n4926) );
  OA22X1 U4839 ( .IN1(n4939), .IN2(n4940), .IN3(n4941), .IN4(n4942), .Q(n4893)
         );
  AND2X1 U4840 ( .IN1(n4940), .IN2(n4939), .Q(n4942) );
  XNOR3X1 U4841 ( .IN1(n4943), .IN2(n4886), .IN3(n4892), .Q(n4895) );
  XOR3X1 U4842 ( .IN1(n4898), .IN2(n4897), .IN3(n4896), .Q(n4892) );
  XNOR3X1 U4843 ( .IN1(n4910), .IN2(n4908), .IN3(n4907), .Q(n4896) );
  NAND2X0 U4844 ( .IN1(n4944), .IN2(n4945), .QN(n4907) );
  MUX21X1 U4845 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1500 ), .Q(n4945) );
  MUX21X1 U4846 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1501 ), .Q(n4944) );
  NAND2X0 U4847 ( .IN1(n4946), .IN2(n4947), .QN(n4908) );
  MUX21X1 U4848 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1503 ), .Q(n4947) );
  MUX21X1 U4849 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1502 ), .Q(n4946) );
  NAND2X0 U4850 ( .IN1(n4948), .IN2(n4949), .QN(n4910) );
  MUX21X1 U4851 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1498 ), .Q(n4949) );
  MUX21X1 U4852 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1499 ), .Q(n4948) );
  AOI22X1 U4853 ( .IN1(n4950), .IN2(n4951), .IN3(n4952), .IN4(n4953), .QN(
        n4897) );
  OR2X1 U4854 ( .IN1(n4951), .IN2(n4950), .Q(n4952) );
  XNOR3X1 U4855 ( .IN1(n4922), .IN2(n4923), .IN3(n4925), .Q(n4898) );
  NAND2X0 U4856 ( .IN1(n4954), .IN2(n4955), .QN(n4925) );
  MUX21X1 U4857 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1492 ), .Q(n4955) );
  MUX21X1 U4858 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1493 ), .Q(n4954) );
  NAND2X0 U4859 ( .IN1(n4956), .IN2(n4957), .QN(n4923) );
  MUX21X1 U4860 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1497 ), .Q(n4957) );
  MUX21X1 U4861 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1496 ), .Q(n4956) );
  NAND2X0 U4862 ( .IN1(n4958), .IN2(n4959), .QN(n4922) );
  MUX21X1 U4863 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1494 ), .Q(n4959) );
  MUX21X1 U4864 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1495 ), .Q(n4958) );
  XOR2X1 U4865 ( .IN1(n4847), .IN2(n4848), .Q(n4886) );
  NAND2X0 U4866 ( .IN1(n4960), .IN2(n4961), .QN(n4848) );
  MUX21X1 U4867 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1488 ), .Q(n4961) );
  MUX21X1 U4868 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1489 ), .Q(n4960) );
  NAND2X0 U4869 ( .IN1(n4962), .IN2(n4963), .QN(n4847) );
  MUX21X1 U4870 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1491 ), .Q(n4963) );
  MUX21X1 U4871 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1490 ), .Q(n4962) );
  XOR2X1 U4872 ( .IN1(n4887), .IN2(n4964), .Q(n4943) );
  NAND2X0 U4873 ( .IN1(n4890), .IN2(n4891), .QN(n4964) );
  AO22X1 U4874 ( .IN1(n4965), .IN2(n4966), .IN3(n4967), .IN4(n4968), .Q(n4887)
         );
  OR2X1 U4875 ( .IN1(n4966), .IN2(n4965), .Q(n4967) );
  AO22X1 U4876 ( .IN1(n4969), .IN2(n4970), .IN3(n4971), .IN4(n3453), .Q(
        \i_m4stg_frac/a1cout[35] ) );
  AO22X1 U4877 ( .IN1(n4972), .IN2(n4973), .IN3(n4974), .IN4(n4975), .Q(n3453)
         );
  OR2X1 U4878 ( .IN1(n4972), .IN2(n4973), .Q(n4975) );
  AND2X1 U4879 ( .IN1(n4976), .IN2(n4977), .Q(n4974) );
  NAND2X0 U4880 ( .IN1(n3454), .IN2(n3452), .QN(n4971) );
  INVX0 U4881 ( .INP(n4969), .ZN(n3452) );
  INVX0 U4882 ( .INP(n3454), .ZN(n4970) );
  MUX21X1 U4883 ( .IN1(n4978), .IN2(n4979), .S(n4980), .Q(n3454) );
  INVX0 U4884 ( .INP(n4981), .ZN(n4980) );
  XOR2X1 U4885 ( .IN1(n4938), .IN2(n4936), .Q(n4969) );
  OA22X1 U4886 ( .IN1(n4982), .IN2(n4983), .IN3(n4984), .IN4(n4985), .Q(n4936)
         );
  AND2X1 U4887 ( .IN1(n4983), .IN2(n4982), .Q(n4985) );
  XNOR3X1 U4888 ( .IN1(n4986), .IN2(n4929), .IN3(n4935), .Q(n4938) );
  XOR3X1 U4889 ( .IN1(n4941), .IN2(n4940), .IN3(n4939), .Q(n4935) );
  XNOR3X1 U4890 ( .IN1(n4953), .IN2(n4951), .IN3(n4950), .Q(n4939) );
  NAND2X0 U4891 ( .IN1(n4987), .IN2(n4988), .QN(n4950) );
  MUX21X1 U4892 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1499 ), .Q(n4988) );
  MUX21X1 U4893 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1500 ), .Q(n4987) );
  NAND2X0 U4894 ( .IN1(n4989), .IN2(n4990), .QN(n4951) );
  MUX21X1 U4895 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1502 ), .Q(n4990) );
  MUX21X1 U4896 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1501 ), .Q(n4989) );
  NAND2X0 U4897 ( .IN1(n4991), .IN2(n4992), .QN(n4953) );
  MUX21X1 U4898 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1497 ), .Q(n4992) );
  MUX21X1 U4899 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1498 ), .Q(n4991) );
  AOI22X1 U4900 ( .IN1(n4993), .IN2(n4994), .IN3(n4995), .IN4(n4996), .QN(
        n4940) );
  OR2X1 U4901 ( .IN1(n4994), .IN2(n4993), .Q(n4995) );
  XNOR3X1 U4902 ( .IN1(n4965), .IN2(n4966), .IN3(n4968), .Q(n4941) );
  NAND2X0 U4903 ( .IN1(n4997), .IN2(n4998), .QN(n4968) );
  MUX21X1 U4904 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1491 ), .Q(n4998) );
  MUX21X1 U4905 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1492 ), .Q(n4997) );
  NAND2X0 U4906 ( .IN1(n4999), .IN2(n5000), .QN(n4966) );
  MUX21X1 U4907 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1496 ), .Q(n5000) );
  MUX21X1 U4908 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1495 ), .Q(n4999) );
  NAND2X0 U4909 ( .IN1(n5001), .IN2(n5002), .QN(n4965) );
  MUX21X1 U4910 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1493 ), .Q(n5002) );
  MUX21X1 U4911 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1494 ), .Q(n5001) );
  XOR2X1 U4912 ( .IN1(n4890), .IN2(n4891), .Q(n4929) );
  NAND2X0 U4913 ( .IN1(n5003), .IN2(n5004), .QN(n4891) );
  MUX21X1 U4914 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1487 ), .Q(n5004) );
  MUX21X1 U4915 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1488 ), .Q(n5003) );
  NAND2X0 U4916 ( .IN1(n5005), .IN2(n5006), .QN(n4890) );
  MUX21X1 U4917 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1490 ), .Q(n5006) );
  MUX21X1 U4918 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1489 ), .Q(n5005) );
  XOR2X1 U4919 ( .IN1(n4930), .IN2(n5007), .Q(n4986) );
  NAND2X0 U4920 ( .IN1(n4933), .IN2(n4934), .QN(n5007) );
  AO22X1 U4921 ( .IN1(n5008), .IN2(n5009), .IN3(n5010), .IN4(n5011), .Q(n4930)
         );
  OR2X1 U4922 ( .IN1(n5009), .IN2(n5008), .Q(n5010) );
  AO22X1 U4923 ( .IN1(n5012), .IN2(n5013), .IN3(n5014), .IN4(n3456), .Q(
        \i_m4stg_frac/a1cout[34] ) );
  AO22X1 U4924 ( .IN1(n5015), .IN2(n5016), .IN3(n5017), .IN4(n5018), .Q(n3456)
         );
  OR2X1 U4925 ( .IN1(n5015), .IN2(n5016), .Q(n5018) );
  AND2X1 U4926 ( .IN1(n5019), .IN2(n5020), .Q(n5017) );
  NAND2X0 U4927 ( .IN1(n3457), .IN2(n3455), .QN(n5014) );
  INVX0 U4928 ( .INP(n5012), .ZN(n3455) );
  INVX0 U4929 ( .INP(n3457), .ZN(n5013) );
  MUX21X1 U4930 ( .IN1(n5021), .IN2(n5022), .S(n5023), .Q(n3457) );
  INVX0 U4931 ( .INP(n5024), .ZN(n5023) );
  XOR2X1 U4932 ( .IN1(n4981), .IN2(n4979), .Q(n5012) );
  OA22X1 U4933 ( .IN1(n5025), .IN2(n5026), .IN3(n5027), .IN4(n5028), .Q(n4979)
         );
  AND2X1 U4934 ( .IN1(n5026), .IN2(n5025), .Q(n5028) );
  XNOR3X1 U4935 ( .IN1(n5029), .IN2(n4972), .IN3(n4978), .Q(n4981) );
  XOR3X1 U4936 ( .IN1(n4984), .IN2(n4983), .IN3(n4982), .Q(n4978) );
  XNOR3X1 U4937 ( .IN1(n4996), .IN2(n4994), .IN3(n4993), .Q(n4982) );
  NAND2X0 U4938 ( .IN1(n5030), .IN2(n5031), .QN(n4993) );
  MUX21X1 U4939 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1498 ), .Q(n5031) );
  MUX21X1 U4940 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1499 ), .Q(n5030) );
  NAND2X0 U4941 ( .IN1(n5032), .IN2(n5033), .QN(n4994) );
  MUX21X1 U4942 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1501 ), .Q(n5033) );
  MUX21X1 U4943 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1500 ), .Q(n5032) );
  NAND2X0 U4944 ( .IN1(n5034), .IN2(n5035), .QN(n4996) );
  MUX21X1 U4945 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1496 ), .Q(n5035) );
  MUX21X1 U4946 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1497 ), .Q(n5034) );
  AOI22X1 U4947 ( .IN1(n5036), .IN2(n5037), .IN3(n5038), .IN4(n5039), .QN(
        n4983) );
  OR2X1 U4948 ( .IN1(n5037), .IN2(n5036), .Q(n5038) );
  XNOR3X1 U4949 ( .IN1(n5008), .IN2(n5009), .IN3(n5011), .Q(n4984) );
  NAND2X0 U4950 ( .IN1(n5040), .IN2(n5041), .QN(n5011) );
  MUX21X1 U4951 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1490 ), .Q(n5041) );
  MUX21X1 U4952 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1491 ), .Q(n5040) );
  NAND2X0 U4953 ( .IN1(n5042), .IN2(n5043), .QN(n5009) );
  MUX21X1 U4954 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1495 ), .Q(n5043) );
  MUX21X1 U4955 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1494 ), .Q(n5042) );
  NAND2X0 U4956 ( .IN1(n5044), .IN2(n5045), .QN(n5008) );
  MUX21X1 U4957 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1492 ), .Q(n5045) );
  MUX21X1 U4958 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1493 ), .Q(n5044) );
  XOR2X1 U4959 ( .IN1(n4933), .IN2(n4934), .Q(n4972) );
  NAND2X0 U4960 ( .IN1(n5046), .IN2(n5047), .QN(n4934) );
  MUX21X1 U4961 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1486 ), .Q(n5047) );
  MUX21X1 U4962 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1487 ), .Q(n5046) );
  NAND2X0 U4963 ( .IN1(n5048), .IN2(n5049), .QN(n4933) );
  MUX21X1 U4964 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1489 ), .Q(n5049) );
  MUX21X1 U4965 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1488 ), .Q(n5048) );
  XOR2X1 U4966 ( .IN1(n4973), .IN2(n5050), .Q(n5029) );
  NAND2X0 U4967 ( .IN1(n4976), .IN2(n4977), .QN(n5050) );
  AO22X1 U4968 ( .IN1(n5051), .IN2(n5052), .IN3(n5053), .IN4(n5054), .Q(n4973)
         );
  OR2X1 U4969 ( .IN1(n5052), .IN2(n5051), .Q(n5053) );
  AO22X1 U4970 ( .IN1(n5055), .IN2(n5056), .IN3(n5057), .IN4(n3459), .Q(
        \i_m4stg_frac/a1cout[33] ) );
  AO22X1 U4971 ( .IN1(n5058), .IN2(n5059), .IN3(n5060), .IN4(n5061), .Q(n3459)
         );
  OR2X1 U4972 ( .IN1(n5058), .IN2(n5059), .Q(n5061) );
  AND2X1 U4973 ( .IN1(n5062), .IN2(n5063), .Q(n5060) );
  NAND2X0 U4974 ( .IN1(n3460), .IN2(n3458), .QN(n5057) );
  INVX0 U4975 ( .INP(n5055), .ZN(n3458) );
  INVX0 U4976 ( .INP(n3460), .ZN(n5056) );
  MUX21X1 U4977 ( .IN1(n5064), .IN2(n5065), .S(n5066), .Q(n3460) );
  INVX0 U4978 ( .INP(n5067), .ZN(n5066) );
  XOR2X1 U4979 ( .IN1(n5024), .IN2(n5022), .Q(n5055) );
  OA22X1 U4980 ( .IN1(n5068), .IN2(n5069), .IN3(n5070), .IN4(n5071), .Q(n5022)
         );
  AND2X1 U4981 ( .IN1(n5069), .IN2(n5068), .Q(n5071) );
  XNOR3X1 U4982 ( .IN1(n5072), .IN2(n5015), .IN3(n5021), .Q(n5024) );
  XOR3X1 U4983 ( .IN1(n5027), .IN2(n5026), .IN3(n5025), .Q(n5021) );
  XNOR3X1 U4984 ( .IN1(n5039), .IN2(n5037), .IN3(n5036), .Q(n5025) );
  NAND2X0 U4985 ( .IN1(n5073), .IN2(n5074), .QN(n5036) );
  MUX21X1 U4986 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1497 ), .Q(n5074) );
  MUX21X1 U4987 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1498 ), .Q(n5073) );
  NAND2X0 U4988 ( .IN1(n5075), .IN2(n5076), .QN(n5037) );
  MUX21X1 U4989 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1500 ), .Q(n5076) );
  MUX21X1 U4990 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1499 ), .Q(n5075) );
  NAND2X0 U4991 ( .IN1(n5077), .IN2(n5078), .QN(n5039) );
  MUX21X1 U4992 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1495 ), .Q(n5078) );
  MUX21X1 U4993 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1496 ), .Q(n5077) );
  AOI22X1 U4994 ( .IN1(n5079), .IN2(n5080), .IN3(n5081), .IN4(n5082), .QN(
        n5026) );
  OR2X1 U4995 ( .IN1(n5080), .IN2(n5079), .Q(n5081) );
  XNOR3X1 U4996 ( .IN1(n5051), .IN2(n5052), .IN3(n5054), .Q(n5027) );
  NAND2X0 U4997 ( .IN1(n5083), .IN2(n5084), .QN(n5054) );
  MUX21X1 U4998 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1489 ), .Q(n5084) );
  MUX21X1 U4999 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1490 ), .Q(n5083) );
  NAND2X0 U5000 ( .IN1(n5085), .IN2(n5086), .QN(n5052) );
  MUX21X1 U5001 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1494 ), .Q(n5086) );
  MUX21X1 U5002 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1493 ), .Q(n5085) );
  NAND2X0 U5003 ( .IN1(n5087), .IN2(n5088), .QN(n5051) );
  MUX21X1 U5004 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1491 ), .Q(n5088) );
  MUX21X1 U5005 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1492 ), .Q(n5087) );
  XOR2X1 U5006 ( .IN1(n4976), .IN2(n4977), .Q(n5015) );
  NAND2X0 U5007 ( .IN1(n5089), .IN2(n5090), .QN(n4977) );
  MUX21X1 U5008 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1485 ), .Q(n5090) );
  MUX21X1 U5009 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1486 ), .Q(n5089) );
  NAND2X0 U5010 ( .IN1(n5091), .IN2(n5092), .QN(n4976) );
  MUX21X1 U5011 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1488 ), .Q(n5092) );
  MUX21X1 U5012 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1487 ), .Q(n5091) );
  XOR2X1 U5013 ( .IN1(n5016), .IN2(n5093), .Q(n5072) );
  NAND2X0 U5014 ( .IN1(n5019), .IN2(n5020), .QN(n5093) );
  AO22X1 U5015 ( .IN1(n5094), .IN2(n5095), .IN3(n5096), .IN4(n5097), .Q(n5016)
         );
  OR2X1 U5016 ( .IN1(n5095), .IN2(n5094), .Q(n5096) );
  AO22X1 U5017 ( .IN1(n5098), .IN2(n5099), .IN3(n5100), .IN4(n3462), .Q(
        \i_m4stg_frac/a1cout[32] ) );
  AO22X1 U5018 ( .IN1(n5101), .IN2(n5102), .IN3(n5103), .IN4(n5104), .Q(n3462)
         );
  OR2X1 U5019 ( .IN1(n5101), .IN2(n5102), .Q(n5104) );
  AND2X1 U5020 ( .IN1(n5105), .IN2(n5106), .Q(n5103) );
  NAND2X0 U5021 ( .IN1(n3463), .IN2(n3461), .QN(n5100) );
  INVX0 U5022 ( .INP(n5098), .ZN(n3461) );
  INVX0 U5023 ( .INP(n3463), .ZN(n5099) );
  MUX21X1 U5024 ( .IN1(n5107), .IN2(n5108), .S(n5109), .Q(n3463) );
  INVX0 U5025 ( .INP(n5110), .ZN(n5109) );
  XOR2X1 U5026 ( .IN1(n5067), .IN2(n5065), .Q(n5098) );
  OA22X1 U5027 ( .IN1(n5111), .IN2(n5112), .IN3(n5113), .IN4(n5114), .Q(n5065)
         );
  AND2X1 U5028 ( .IN1(n5112), .IN2(n5111), .Q(n5114) );
  XNOR3X1 U5029 ( .IN1(n5115), .IN2(n5058), .IN3(n5064), .Q(n5067) );
  XOR3X1 U5030 ( .IN1(n5070), .IN2(n5069), .IN3(n5068), .Q(n5064) );
  XNOR3X1 U5031 ( .IN1(n5082), .IN2(n5080), .IN3(n5079), .Q(n5068) );
  NAND2X0 U5032 ( .IN1(n5116), .IN2(n5117), .QN(n5079) );
  MUX21X1 U5033 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1496 ), .Q(n5117) );
  MUX21X1 U5034 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1497 ), .Q(n5116) );
  NAND2X0 U5035 ( .IN1(n5118), .IN2(n5119), .QN(n5080) );
  MUX21X1 U5036 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1499 ), .Q(n5119) );
  MUX21X1 U5037 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1498 ), .Q(n5118) );
  NAND2X0 U5038 ( .IN1(n5120), .IN2(n5121), .QN(n5082) );
  MUX21X1 U5039 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1494 ), .Q(n5121) );
  MUX21X1 U5040 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1495 ), .Q(n5120) );
  AOI22X1 U5041 ( .IN1(n5122), .IN2(n5123), .IN3(n5124), .IN4(n5125), .QN(
        n5069) );
  OR2X1 U5042 ( .IN1(n5123), .IN2(n5122), .Q(n5124) );
  XNOR3X1 U5043 ( .IN1(n5094), .IN2(n5095), .IN3(n5097), .Q(n5070) );
  NAND2X0 U5044 ( .IN1(n5126), .IN2(n5127), .QN(n5097) );
  MUX21X1 U5045 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1488 ), .Q(n5127) );
  MUX21X1 U5046 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1489 ), .Q(n5126) );
  NAND2X0 U5047 ( .IN1(n5128), .IN2(n5129), .QN(n5095) );
  MUX21X1 U5048 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1493 ), .Q(n5129) );
  MUX21X1 U5049 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1492 ), .Q(n5128) );
  NAND2X0 U5050 ( .IN1(n5130), .IN2(n5131), .QN(n5094) );
  MUX21X1 U5051 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1490 ), .Q(n5131) );
  MUX21X1 U5052 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1491 ), .Q(n5130) );
  XOR2X1 U5053 ( .IN1(n5019), .IN2(n5020), .Q(n5058) );
  NAND2X0 U5054 ( .IN1(n5132), .IN2(n5133), .QN(n5020) );
  MUX21X1 U5055 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1484 ), .Q(n5133) );
  MUX21X1 U5056 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1485 ), .Q(n5132) );
  NAND2X0 U5057 ( .IN1(n5134), .IN2(n5135), .QN(n5019) );
  MUX21X1 U5058 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1487 ), .Q(n5135) );
  MUX21X1 U5059 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1486 ), .Q(n5134) );
  XOR2X1 U5060 ( .IN1(n5059), .IN2(n5136), .Q(n5115) );
  NAND2X0 U5061 ( .IN1(n5062), .IN2(n5063), .QN(n5136) );
  AO22X1 U5062 ( .IN1(n5137), .IN2(n5138), .IN3(n5139), .IN4(n5140), .Q(n5059)
         );
  OR2X1 U5063 ( .IN1(n5138), .IN2(n5137), .Q(n5139) );
  AO22X1 U5064 ( .IN1(n5141), .IN2(n5142), .IN3(n5143), .IN4(n3465), .Q(
        \i_m4stg_frac/a1cout[31] ) );
  AO22X1 U5065 ( .IN1(n5144), .IN2(n5145), .IN3(n5146), .IN4(n5147), .Q(n3465)
         );
  OR2X1 U5066 ( .IN1(n5144), .IN2(n5145), .Q(n5147) );
  AND2X1 U5067 ( .IN1(n5148), .IN2(n5149), .Q(n5146) );
  NAND2X0 U5068 ( .IN1(n3466), .IN2(n3464), .QN(n5143) );
  INVX0 U5069 ( .INP(n5141), .ZN(n3464) );
  INVX0 U5070 ( .INP(n3466), .ZN(n5142) );
  MUX21X1 U5071 ( .IN1(n5150), .IN2(n5151), .S(n5152), .Q(n3466) );
  INVX0 U5072 ( .INP(n5153), .ZN(n5152) );
  XOR2X1 U5073 ( .IN1(n5110), .IN2(n5108), .Q(n5141) );
  OA22X1 U5074 ( .IN1(n5154), .IN2(n5155), .IN3(n5156), .IN4(n5157), .Q(n5108)
         );
  AND2X1 U5075 ( .IN1(n5155), .IN2(n5154), .Q(n5157) );
  XNOR3X1 U5076 ( .IN1(n5158), .IN2(n5101), .IN3(n5107), .Q(n5110) );
  XOR3X1 U5077 ( .IN1(n5113), .IN2(n5112), .IN3(n5111), .Q(n5107) );
  XNOR3X1 U5078 ( .IN1(n5125), .IN2(n5123), .IN3(n5122), .Q(n5111) );
  NAND2X0 U5079 ( .IN1(n5159), .IN2(n5160), .QN(n5122) );
  MUX21X1 U5080 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1495 ), .Q(n5160) );
  MUX21X1 U5081 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1496 ), .Q(n5159) );
  NAND2X0 U5082 ( .IN1(n5161), .IN2(n5162), .QN(n5123) );
  MUX21X1 U5083 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1498 ), .Q(n5162) );
  MUX21X1 U5084 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1497 ), .Q(n5161) );
  NAND2X0 U5085 ( .IN1(n5163), .IN2(n5164), .QN(n5125) );
  MUX21X1 U5086 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1493 ), .Q(n5164) );
  MUX21X1 U5087 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1494 ), .Q(n5163) );
  AOI22X1 U5088 ( .IN1(n5165), .IN2(n5166), .IN3(n5167), .IN4(n5168), .QN(
        n5112) );
  OR2X1 U5089 ( .IN1(n5166), .IN2(n5165), .Q(n5167) );
  XNOR3X1 U5090 ( .IN1(n5137), .IN2(n5138), .IN3(n5140), .Q(n5113) );
  NAND2X0 U5091 ( .IN1(n5169), .IN2(n5170), .QN(n5140) );
  MUX21X1 U5092 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1487 ), .Q(n5170) );
  MUX21X1 U5093 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1488 ), .Q(n5169) );
  NAND2X0 U5094 ( .IN1(n5171), .IN2(n5172), .QN(n5138) );
  MUX21X1 U5095 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1492 ), .Q(n5172) );
  MUX21X1 U5096 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1491 ), .Q(n5171) );
  NAND2X0 U5097 ( .IN1(n5173), .IN2(n5174), .QN(n5137) );
  MUX21X1 U5098 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1489 ), .Q(n5174) );
  MUX21X1 U5099 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1490 ), .Q(n5173) );
  XOR2X1 U5100 ( .IN1(n5062), .IN2(n5063), .Q(n5101) );
  NAND2X0 U5101 ( .IN1(n5175), .IN2(n5176), .QN(n5063) );
  MUX21X1 U5102 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1483 ), .Q(n5176) );
  MUX21X1 U5103 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1484 ), .Q(n5175) );
  NAND2X0 U5104 ( .IN1(n5177), .IN2(n5178), .QN(n5062) );
  MUX21X1 U5105 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1486 ), .Q(n5178) );
  MUX21X1 U5106 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1485 ), .Q(n5177) );
  XOR2X1 U5107 ( .IN1(n5102), .IN2(n5179), .Q(n5158) );
  NAND2X0 U5108 ( .IN1(n5105), .IN2(n5106), .QN(n5179) );
  AO22X1 U5109 ( .IN1(n5180), .IN2(n5181), .IN3(n5182), .IN4(n5183), .Q(n5102)
         );
  OR2X1 U5110 ( .IN1(n5181), .IN2(n5180), .Q(n5182) );
  AO22X1 U5111 ( .IN1(n5184), .IN2(n5185), .IN3(n5186), .IN4(n3468), .Q(
        \i_m4stg_frac/a1cout[30] ) );
  AO22X1 U5112 ( .IN1(n5187), .IN2(n5188), .IN3(n5189), .IN4(n5190), .Q(n3468)
         );
  OR2X1 U5113 ( .IN1(n5187), .IN2(n5188), .Q(n5190) );
  AND2X1 U5114 ( .IN1(n5191), .IN2(n5192), .Q(n5189) );
  NAND2X0 U5115 ( .IN1(n3469), .IN2(n3467), .QN(n5186) );
  INVX0 U5116 ( .INP(n5184), .ZN(n3467) );
  INVX0 U5117 ( .INP(n3469), .ZN(n5185) );
  MUX21X1 U5118 ( .IN1(n5193), .IN2(n5194), .S(n5195), .Q(n3469) );
  INVX0 U5119 ( .INP(n5196), .ZN(n5195) );
  XOR2X1 U5120 ( .IN1(n5153), .IN2(n5151), .Q(n5184) );
  OA22X1 U5121 ( .IN1(n5197), .IN2(n5198), .IN3(n5199), .IN4(n5200), .Q(n5151)
         );
  AND2X1 U5122 ( .IN1(n5198), .IN2(n5197), .Q(n5200) );
  XNOR3X1 U5123 ( .IN1(n5201), .IN2(n5144), .IN3(n5150), .Q(n5153) );
  XOR3X1 U5124 ( .IN1(n5156), .IN2(n5155), .IN3(n5154), .Q(n5150) );
  XNOR3X1 U5125 ( .IN1(n5168), .IN2(n5166), .IN3(n5165), .Q(n5154) );
  NAND2X0 U5126 ( .IN1(n5202), .IN2(n5203), .QN(n5165) );
  MUX21X1 U5127 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1494 ), .Q(n5203) );
  MUX21X1 U5128 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1495 ), .Q(n5202) );
  NAND2X0 U5129 ( .IN1(n5204), .IN2(n5205), .QN(n5166) );
  MUX21X1 U5130 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1497 ), .Q(n5205) );
  MUX21X1 U5131 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1496 ), .Q(n5204) );
  NAND2X0 U5132 ( .IN1(n5206), .IN2(n5207), .QN(n5168) );
  MUX21X1 U5133 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1492 ), .Q(n5207) );
  MUX21X1 U5134 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1493 ), .Q(n5206) );
  AOI22X1 U5135 ( .IN1(n5208), .IN2(n5209), .IN3(n5210), .IN4(n5211), .QN(
        n5155) );
  OR2X1 U5136 ( .IN1(n5209), .IN2(n5208), .Q(n5210) );
  XNOR3X1 U5137 ( .IN1(n5180), .IN2(n5181), .IN3(n5183), .Q(n5156) );
  NAND2X0 U5138 ( .IN1(n5212), .IN2(n5213), .QN(n5183) );
  MUX21X1 U5139 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1486 ), .Q(n5213) );
  MUX21X1 U5140 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1487 ), .Q(n5212) );
  NAND2X0 U5141 ( .IN1(n5214), .IN2(n5215), .QN(n5181) );
  MUX21X1 U5142 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1491 ), .Q(n5215) );
  MUX21X1 U5143 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1490 ), .Q(n5214) );
  NAND2X0 U5144 ( .IN1(n5216), .IN2(n5217), .QN(n5180) );
  MUX21X1 U5145 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1488 ), .Q(n5217) );
  MUX21X1 U5146 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1489 ), .Q(n5216) );
  XOR2X1 U5147 ( .IN1(n5105), .IN2(n5106), .Q(n5144) );
  NAND2X0 U5148 ( .IN1(n5218), .IN2(n5219), .QN(n5106) );
  MUX21X1 U5149 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1482 ), .Q(n5219) );
  MUX21X1 U5150 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1483 ), .Q(n5218) );
  NAND2X0 U5151 ( .IN1(n5220), .IN2(n5221), .QN(n5105) );
  MUX21X1 U5152 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1485 ), .Q(n5221) );
  MUX21X1 U5153 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1484 ), .Q(n5220) );
  XOR2X1 U5154 ( .IN1(n5145), .IN2(n5222), .Q(n5201) );
  NAND2X0 U5155 ( .IN1(n5148), .IN2(n5149), .QN(n5222) );
  AO22X1 U5156 ( .IN1(n5223), .IN2(n5224), .IN3(n5225), .IN4(n5226), .Q(n5145)
         );
  OR2X1 U5157 ( .IN1(n5224), .IN2(n5223), .Q(n5225) );
  AO22X1 U5158 ( .IN1(n5227), .IN2(n5228), .IN3(n5229), .IN4(n3473), .Q(
        \i_m4stg_frac/a1cout[29] ) );
  AO22X1 U5159 ( .IN1(n5230), .IN2(n5231), .IN3(n5232), .IN4(n5233), .Q(n3473)
         );
  OR2X1 U5160 ( .IN1(n5230), .IN2(n5231), .Q(n5233) );
  AND2X1 U5161 ( .IN1(n5234), .IN2(n5235), .Q(n5232) );
  NAND2X0 U5162 ( .IN1(n3474), .IN2(n3472), .QN(n5229) );
  INVX0 U5163 ( .INP(n5227), .ZN(n3472) );
  INVX0 U5164 ( .INP(n3474), .ZN(n5228) );
  MUX21X1 U5165 ( .IN1(n5236), .IN2(n5237), .S(n5238), .Q(n3474) );
  INVX0 U5166 ( .INP(n5239), .ZN(n5238) );
  XOR2X1 U5167 ( .IN1(n5196), .IN2(n5194), .Q(n5227) );
  OA22X1 U5168 ( .IN1(n5240), .IN2(n5241), .IN3(n5242), .IN4(n5243), .Q(n5194)
         );
  AND2X1 U5169 ( .IN1(n5241), .IN2(n5240), .Q(n5243) );
  XNOR3X1 U5170 ( .IN1(n5244), .IN2(n5187), .IN3(n5193), .Q(n5196) );
  XOR3X1 U5171 ( .IN1(n5199), .IN2(n5198), .IN3(n5197), .Q(n5193) );
  XNOR3X1 U5172 ( .IN1(n5211), .IN2(n5209), .IN3(n5208), .Q(n5197) );
  NAND2X0 U5173 ( .IN1(n5245), .IN2(n5246), .QN(n5208) );
  MUX21X1 U5174 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1493 ), .Q(n5246) );
  MUX21X1 U5175 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1494 ), .Q(n5245) );
  NAND2X0 U5176 ( .IN1(n5247), .IN2(n5248), .QN(n5209) );
  MUX21X1 U5177 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1496 ), .Q(n5248) );
  MUX21X1 U5178 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1495 ), .Q(n5247) );
  NAND2X0 U5179 ( .IN1(n5249), .IN2(n5250), .QN(n5211) );
  MUX21X1 U5180 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1491 ), .Q(n5250) );
  MUX21X1 U5181 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1492 ), .Q(n5249) );
  AOI22X1 U5182 ( .IN1(n5251), .IN2(n5252), .IN3(n5253), .IN4(n5254), .QN(
        n5198) );
  OR2X1 U5183 ( .IN1(n5252), .IN2(n5251), .Q(n5253) );
  XNOR3X1 U5184 ( .IN1(n5223), .IN2(n5224), .IN3(n5226), .Q(n5199) );
  NAND2X0 U5185 ( .IN1(n5255), .IN2(n5256), .QN(n5226) );
  MUX21X1 U5186 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1485 ), .Q(n5256) );
  MUX21X1 U5187 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1486 ), .Q(n5255) );
  NAND2X0 U5188 ( .IN1(n5257), .IN2(n5258), .QN(n5224) );
  MUX21X1 U5189 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1490 ), .Q(n5258) );
  MUX21X1 U5190 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1489 ), .Q(n5257) );
  NAND2X0 U5191 ( .IN1(n5259), .IN2(n5260), .QN(n5223) );
  MUX21X1 U5192 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1487 ), .Q(n5260) );
  MUX21X1 U5193 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1488 ), .Q(n5259) );
  XOR2X1 U5194 ( .IN1(n5148), .IN2(n5149), .Q(n5187) );
  NAND2X0 U5195 ( .IN1(n5261), .IN2(n5262), .QN(n5149) );
  MUX21X1 U5196 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1481 ), .Q(n5262) );
  MUX21X1 U5197 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1482 ), .Q(n5261) );
  NAND2X0 U5198 ( .IN1(n5263), .IN2(n5264), .QN(n5148) );
  MUX21X1 U5199 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1484 ), .Q(n5264) );
  MUX21X1 U5200 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1483 ), .Q(n5263) );
  XOR2X1 U5201 ( .IN1(n5188), .IN2(n5265), .Q(n5244) );
  NAND2X0 U5202 ( .IN1(n5191), .IN2(n5192), .QN(n5265) );
  AO22X1 U5203 ( .IN1(n5266), .IN2(n5267), .IN3(n5268), .IN4(n5269), .Q(n5188)
         );
  OR2X1 U5204 ( .IN1(n5267), .IN2(n5266), .Q(n5268) );
  AO22X1 U5205 ( .IN1(n5270), .IN2(n5271), .IN3(n5272), .IN4(n3476), .Q(
        \i_m4stg_frac/a1cout[28] ) );
  AO22X1 U5206 ( .IN1(n5273), .IN2(n5274), .IN3(n5275), .IN4(n5276), .Q(n3476)
         );
  OR2X1 U5207 ( .IN1(n5273), .IN2(n5274), .Q(n5276) );
  AND2X1 U5208 ( .IN1(n5277), .IN2(n5278), .Q(n5275) );
  NAND2X0 U5209 ( .IN1(n3477), .IN2(n3475), .QN(n5272) );
  INVX0 U5210 ( .INP(n5270), .ZN(n3475) );
  INVX0 U5211 ( .INP(n3477), .ZN(n5271) );
  MUX21X1 U5212 ( .IN1(n5279), .IN2(n5280), .S(n5281), .Q(n3477) );
  INVX0 U5213 ( .INP(n5282), .ZN(n5281) );
  XOR2X1 U5214 ( .IN1(n5239), .IN2(n5237), .Q(n5270) );
  OA22X1 U5215 ( .IN1(n5283), .IN2(n5284), .IN3(n5285), .IN4(n5286), .Q(n5237)
         );
  AND2X1 U5216 ( .IN1(n5284), .IN2(n5283), .Q(n5286) );
  XNOR3X1 U5217 ( .IN1(n5287), .IN2(n5230), .IN3(n5236), .Q(n5239) );
  XOR3X1 U5218 ( .IN1(n5242), .IN2(n5241), .IN3(n5240), .Q(n5236) );
  XNOR3X1 U5219 ( .IN1(n5254), .IN2(n5252), .IN3(n5251), .Q(n5240) );
  NAND2X0 U5220 ( .IN1(n5288), .IN2(n5289), .QN(n5251) );
  MUX21X1 U5221 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1492 ), .Q(n5289) );
  MUX21X1 U5222 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1493 ), .Q(n5288) );
  NAND2X0 U5223 ( .IN1(n5290), .IN2(n5291), .QN(n5252) );
  MUX21X1 U5224 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1495 ), .Q(n5291) );
  MUX21X1 U5225 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1494 ), .Q(n5290) );
  NAND2X0 U5226 ( .IN1(n5292), .IN2(n5293), .QN(n5254) );
  MUX21X1 U5227 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1490 ), .Q(n5293) );
  MUX21X1 U5228 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1491 ), .Q(n5292) );
  AOI22X1 U5229 ( .IN1(n5294), .IN2(n5295), .IN3(n5296), .IN4(n5297), .QN(
        n5241) );
  OR2X1 U5230 ( .IN1(n5295), .IN2(n5294), .Q(n5296) );
  XNOR3X1 U5231 ( .IN1(n5266), .IN2(n5267), .IN3(n5269), .Q(n5242) );
  NAND2X0 U5232 ( .IN1(n5298), .IN2(n5299), .QN(n5269) );
  MUX21X1 U5233 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1484 ), .Q(n5299) );
  MUX21X1 U5234 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1485 ), .Q(n5298) );
  NAND2X0 U5235 ( .IN1(n5300), .IN2(n5301), .QN(n5267) );
  MUX21X1 U5236 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1489 ), .Q(n5301) );
  MUX21X1 U5237 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1488 ), .Q(n5300) );
  NAND2X0 U5238 ( .IN1(n5302), .IN2(n5303), .QN(n5266) );
  MUX21X1 U5239 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1486 ), .Q(n5303) );
  MUX21X1 U5240 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1487 ), .Q(n5302) );
  XOR2X1 U5241 ( .IN1(n5191), .IN2(n5192), .Q(n5230) );
  NAND2X0 U5242 ( .IN1(n5304), .IN2(n5305), .QN(n5192) );
  MUX21X1 U5243 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1480 ), .Q(n5305) );
  MUX21X1 U5244 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1481 ), .Q(n5304) );
  NAND2X0 U5245 ( .IN1(n5306), .IN2(n5307), .QN(n5191) );
  MUX21X1 U5246 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1483 ), .Q(n5307) );
  MUX21X1 U5247 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1482 ), .Q(n5306) );
  XOR2X1 U5248 ( .IN1(n5231), .IN2(n5308), .Q(n5287) );
  NAND2X0 U5249 ( .IN1(n5234), .IN2(n5235), .QN(n5308) );
  AO22X1 U5250 ( .IN1(n5309), .IN2(n5310), .IN3(n5311), .IN4(n5312), .Q(n5231)
         );
  OR2X1 U5251 ( .IN1(n5310), .IN2(n5309), .Q(n5311) );
  AO22X1 U5252 ( .IN1(n5313), .IN2(n5314), .IN3(n5315), .IN4(n3479), .Q(
        \i_m4stg_frac/a1cout[27] ) );
  AO22X1 U5253 ( .IN1(n5316), .IN2(n5317), .IN3(n5318), .IN4(n5319), .Q(n3479)
         );
  OR2X1 U5254 ( .IN1(n5316), .IN2(n5317), .Q(n5319) );
  AND2X1 U5255 ( .IN1(n5320), .IN2(n5321), .Q(n5318) );
  NAND2X0 U5256 ( .IN1(n3480), .IN2(n3478), .QN(n5315) );
  INVX0 U5257 ( .INP(n5313), .ZN(n3478) );
  INVX0 U5258 ( .INP(n3480), .ZN(n5314) );
  MUX21X1 U5259 ( .IN1(n5322), .IN2(n5323), .S(n5324), .Q(n3480) );
  INVX0 U5260 ( .INP(n5325), .ZN(n5324) );
  XOR2X1 U5261 ( .IN1(n5282), .IN2(n5280), .Q(n5313) );
  OA22X1 U5262 ( .IN1(n5326), .IN2(n5327), .IN3(n5328), .IN4(n5329), .Q(n5280)
         );
  AND2X1 U5263 ( .IN1(n5327), .IN2(n5326), .Q(n5329) );
  XNOR3X1 U5264 ( .IN1(n5330), .IN2(n5273), .IN3(n5279), .Q(n5282) );
  XOR3X1 U5265 ( .IN1(n5285), .IN2(n5284), .IN3(n5283), .Q(n5279) );
  XNOR3X1 U5266 ( .IN1(n5297), .IN2(n5295), .IN3(n5294), .Q(n5283) );
  NAND2X0 U5267 ( .IN1(n5331), .IN2(n5332), .QN(n5294) );
  MUX21X1 U5268 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1491 ), .Q(n5332) );
  MUX21X1 U5269 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1492 ), .Q(n5331) );
  NAND2X0 U5270 ( .IN1(n5333), .IN2(n5334), .QN(n5295) );
  MUX21X1 U5271 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1494 ), .Q(n5334) );
  MUX21X1 U5272 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1493 ), .Q(n5333) );
  NAND2X0 U5273 ( .IN1(n5335), .IN2(n5336), .QN(n5297) );
  MUX21X1 U5274 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1489 ), .Q(n5336) );
  MUX21X1 U5275 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1490 ), .Q(n5335) );
  AOI22X1 U5276 ( .IN1(n5337), .IN2(n5338), .IN3(n5339), .IN4(n5340), .QN(
        n5284) );
  OR2X1 U5277 ( .IN1(n5338), .IN2(n5337), .Q(n5339) );
  XNOR3X1 U5278 ( .IN1(n5309), .IN2(n5310), .IN3(n5312), .Q(n5285) );
  NAND2X0 U5279 ( .IN1(n5341), .IN2(n5342), .QN(n5312) );
  MUX21X1 U5280 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1483 ), .Q(n5342) );
  MUX21X1 U5281 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1484 ), .Q(n5341) );
  NAND2X0 U5282 ( .IN1(n5343), .IN2(n5344), .QN(n5310) );
  MUX21X1 U5283 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1488 ), .Q(n5344) );
  MUX21X1 U5284 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1487 ), .Q(n5343) );
  NAND2X0 U5285 ( .IN1(n5345), .IN2(n5346), .QN(n5309) );
  MUX21X1 U5286 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1485 ), .Q(n5346) );
  MUX21X1 U5287 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1486 ), .Q(n5345) );
  XOR2X1 U5288 ( .IN1(n5234), .IN2(n5235), .Q(n5273) );
  NAND2X0 U5289 ( .IN1(n5347), .IN2(n5348), .QN(n5235) );
  MUX21X1 U5290 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1479 ), .Q(n5348) );
  MUX21X1 U5291 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1480 ), .Q(n5347) );
  NAND2X0 U5292 ( .IN1(n5349), .IN2(n5350), .QN(n5234) );
  MUX21X1 U5293 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1482 ), .Q(n5350) );
  MUX21X1 U5294 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1481 ), .Q(n5349) );
  XOR2X1 U5295 ( .IN1(n5274), .IN2(n5351), .Q(n5330) );
  NAND2X0 U5296 ( .IN1(n5277), .IN2(n5278), .QN(n5351) );
  AO22X1 U5297 ( .IN1(n5352), .IN2(n5353), .IN3(n5354), .IN4(n5355), .Q(n5274)
         );
  OR2X1 U5298 ( .IN1(n5353), .IN2(n5352), .Q(n5354) );
  AO22X1 U5299 ( .IN1(n5356), .IN2(n5357), .IN3(n5358), .IN4(n3482), .Q(
        \i_m4stg_frac/a1cout[26] ) );
  AO22X1 U5300 ( .IN1(n5359), .IN2(n5360), .IN3(n5361), .IN4(n5362), .Q(n3482)
         );
  OR2X1 U5301 ( .IN1(n5359), .IN2(n5360), .Q(n5362) );
  AND2X1 U5302 ( .IN1(n5363), .IN2(n5364), .Q(n5361) );
  NAND2X0 U5303 ( .IN1(n3483), .IN2(n3481), .QN(n5358) );
  INVX0 U5304 ( .INP(n5356), .ZN(n3481) );
  INVX0 U5305 ( .INP(n3483), .ZN(n5357) );
  MUX21X1 U5306 ( .IN1(n5365), .IN2(n5366), .S(n5367), .Q(n3483) );
  INVX0 U5307 ( .INP(n5368), .ZN(n5367) );
  XOR2X1 U5308 ( .IN1(n5325), .IN2(n5323), .Q(n5356) );
  OA22X1 U5309 ( .IN1(n5369), .IN2(n5370), .IN3(n5371), .IN4(n5372), .Q(n5323)
         );
  AND2X1 U5310 ( .IN1(n5370), .IN2(n5369), .Q(n5372) );
  XNOR3X1 U5311 ( .IN1(n5373), .IN2(n5316), .IN3(n5322), .Q(n5325) );
  XOR3X1 U5312 ( .IN1(n5328), .IN2(n5327), .IN3(n5326), .Q(n5322) );
  XNOR3X1 U5313 ( .IN1(n5340), .IN2(n5338), .IN3(n5337), .Q(n5326) );
  NAND2X0 U5314 ( .IN1(n5374), .IN2(n5375), .QN(n5337) );
  MUX21X1 U5315 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1490 ), .Q(n5375) );
  MUX21X1 U5316 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1491 ), .Q(n5374) );
  NAND2X0 U5317 ( .IN1(n5376), .IN2(n5377), .QN(n5338) );
  MUX21X1 U5318 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1493 ), .Q(n5377) );
  MUX21X1 U5319 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1492 ), .Q(n5376) );
  NAND2X0 U5320 ( .IN1(n5378), .IN2(n5379), .QN(n5340) );
  MUX21X1 U5321 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1488 ), .Q(n5379) );
  MUX21X1 U5322 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1489 ), .Q(n5378) );
  AOI22X1 U5323 ( .IN1(n5380), .IN2(n5381), .IN3(n5382), .IN4(n5383), .QN(
        n5327) );
  OR2X1 U5324 ( .IN1(n5381), .IN2(n5380), .Q(n5382) );
  XNOR3X1 U5325 ( .IN1(n5352), .IN2(n5353), .IN3(n5355), .Q(n5328) );
  NAND2X0 U5326 ( .IN1(n5384), .IN2(n5385), .QN(n5355) );
  MUX21X1 U5327 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1482 ), .Q(n5385) );
  MUX21X1 U5328 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1483 ), .Q(n5384) );
  NAND2X0 U5329 ( .IN1(n5386), .IN2(n5387), .QN(n5353) );
  MUX21X1 U5330 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1487 ), .Q(n5387) );
  MUX21X1 U5331 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1486 ), .Q(n5386) );
  NAND2X0 U5332 ( .IN1(n5388), .IN2(n5389), .QN(n5352) );
  MUX21X1 U5333 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1484 ), .Q(n5389) );
  MUX21X1 U5334 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1485 ), .Q(n5388) );
  XOR2X1 U5335 ( .IN1(n5277), .IN2(n5278), .Q(n5316) );
  NAND2X0 U5336 ( .IN1(n5390), .IN2(n5391), .QN(n5278) );
  MUX21X1 U5337 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1478 ), .Q(n5391) );
  MUX21X1 U5338 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1479 ), .Q(n5390) );
  NAND2X0 U5339 ( .IN1(n5392), .IN2(n5393), .QN(n5277) );
  MUX21X1 U5340 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1481 ), .Q(n5393) );
  MUX21X1 U5341 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1480 ), .Q(n5392) );
  XOR2X1 U5342 ( .IN1(n5317), .IN2(n5394), .Q(n5373) );
  NAND2X0 U5343 ( .IN1(n5320), .IN2(n5321), .QN(n5394) );
  AO22X1 U5344 ( .IN1(n5395), .IN2(n5396), .IN3(n5397), .IN4(n5398), .Q(n5317)
         );
  OR2X1 U5345 ( .IN1(n5396), .IN2(n5395), .Q(n5397) );
  AO22X1 U5346 ( .IN1(n5399), .IN2(n5400), .IN3(n5401), .IN4(n3485), .Q(
        \i_m4stg_frac/a1cout[25] ) );
  AO22X1 U5347 ( .IN1(n5402), .IN2(n5403), .IN3(n5404), .IN4(n5405), .Q(n3485)
         );
  OR2X1 U5348 ( .IN1(n5402), .IN2(n5403), .Q(n5405) );
  AND2X1 U5349 ( .IN1(n5406), .IN2(n5407), .Q(n5404) );
  NAND2X0 U5350 ( .IN1(n3486), .IN2(n3484), .QN(n5401) );
  INVX0 U5351 ( .INP(n5399), .ZN(n3484) );
  INVX0 U5352 ( .INP(n3486), .ZN(n5400) );
  MUX21X1 U5353 ( .IN1(n5408), .IN2(n5409), .S(n5410), .Q(n3486) );
  INVX0 U5354 ( .INP(n5411), .ZN(n5410) );
  XOR2X1 U5355 ( .IN1(n5368), .IN2(n5366), .Q(n5399) );
  OA22X1 U5356 ( .IN1(n5412), .IN2(n5413), .IN3(n5414), .IN4(n5415), .Q(n5366)
         );
  AND2X1 U5357 ( .IN1(n5413), .IN2(n5412), .Q(n5415) );
  XNOR3X1 U5358 ( .IN1(n5416), .IN2(n5359), .IN3(n5365), .Q(n5368) );
  XOR3X1 U5359 ( .IN1(n5371), .IN2(n5370), .IN3(n5369), .Q(n5365) );
  XNOR3X1 U5360 ( .IN1(n5383), .IN2(n5381), .IN3(n5380), .Q(n5369) );
  NAND2X0 U5361 ( .IN1(n5417), .IN2(n5418), .QN(n5380) );
  MUX21X1 U5362 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1489 ), .Q(n5418) );
  MUX21X1 U5363 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1490 ), .Q(n5417) );
  NAND2X0 U5364 ( .IN1(n5419), .IN2(n5420), .QN(n5381) );
  MUX21X1 U5365 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1492 ), .Q(n5420) );
  MUX21X1 U5366 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1491 ), .Q(n5419) );
  NAND2X0 U5367 ( .IN1(n5421), .IN2(n5422), .QN(n5383) );
  MUX21X1 U5368 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1487 ), .Q(n5422) );
  MUX21X1 U5369 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1488 ), .Q(n5421) );
  AOI22X1 U5370 ( .IN1(n5423), .IN2(n5424), .IN3(n5425), .IN4(n5426), .QN(
        n5370) );
  OR2X1 U5371 ( .IN1(n5424), .IN2(n5423), .Q(n5425) );
  XNOR3X1 U5372 ( .IN1(n5395), .IN2(n5396), .IN3(n5398), .Q(n5371) );
  NAND2X0 U5373 ( .IN1(n5427), .IN2(n5428), .QN(n5398) );
  MUX21X1 U5374 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1481 ), .Q(n5428) );
  MUX21X1 U5375 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1482 ), .Q(n5427) );
  NAND2X0 U5376 ( .IN1(n5429), .IN2(n5430), .QN(n5396) );
  MUX21X1 U5377 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1486 ), .Q(n5430) );
  MUX21X1 U5378 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1485 ), .Q(n5429) );
  NAND2X0 U5379 ( .IN1(n5431), .IN2(n5432), .QN(n5395) );
  MUX21X1 U5380 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1483 ), .Q(n5432) );
  MUX21X1 U5381 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1484 ), .Q(n5431) );
  XOR2X1 U5382 ( .IN1(n5320), .IN2(n5321), .Q(n5359) );
  NAND2X0 U5383 ( .IN1(n5433), .IN2(n5434), .QN(n5321) );
  MUX21X1 U5384 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1477 ), .Q(n5434) );
  MUX21X1 U5385 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1478 ), .Q(n5433) );
  NAND2X0 U5386 ( .IN1(n5435), .IN2(n5436), .QN(n5320) );
  MUX21X1 U5387 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1480 ), .Q(n5436) );
  MUX21X1 U5388 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1479 ), .Q(n5435) );
  XOR2X1 U5389 ( .IN1(n5360), .IN2(n5437), .Q(n5416) );
  NAND2X0 U5390 ( .IN1(n5363), .IN2(n5364), .QN(n5437) );
  AO22X1 U5391 ( .IN1(n5438), .IN2(n5439), .IN3(n5440), .IN4(n5441), .Q(n5360)
         );
  OR2X1 U5392 ( .IN1(n5439), .IN2(n5438), .Q(n5440) );
  AO22X1 U5393 ( .IN1(n5442), .IN2(n5443), .IN3(n5444), .IN4(n3488), .Q(
        \i_m4stg_frac/a1cout[24] ) );
  AO22X1 U5394 ( .IN1(n5445), .IN2(n5446), .IN3(n5447), .IN4(n5448), .Q(n3488)
         );
  OR2X1 U5395 ( .IN1(n5445), .IN2(n5446), .Q(n5448) );
  AND2X1 U5396 ( .IN1(n5449), .IN2(n5450), .Q(n5447) );
  NAND2X0 U5397 ( .IN1(n3489), .IN2(n3487), .QN(n5444) );
  INVX0 U5398 ( .INP(n5442), .ZN(n3487) );
  INVX0 U5399 ( .INP(n3489), .ZN(n5443) );
  MUX21X1 U5400 ( .IN1(n5451), .IN2(n5452), .S(n5453), .Q(n3489) );
  INVX0 U5401 ( .INP(n5454), .ZN(n5453) );
  XOR2X1 U5402 ( .IN1(n5411), .IN2(n5409), .Q(n5442) );
  OA22X1 U5403 ( .IN1(n5455), .IN2(n5456), .IN3(n5457), .IN4(n5458), .Q(n5409)
         );
  AND2X1 U5404 ( .IN1(n5456), .IN2(n5455), .Q(n5458) );
  XNOR3X1 U5405 ( .IN1(n5459), .IN2(n5402), .IN3(n5408), .Q(n5411) );
  XOR3X1 U5406 ( .IN1(n5414), .IN2(n5413), .IN3(n5412), .Q(n5408) );
  XNOR3X1 U5407 ( .IN1(n5426), .IN2(n5424), .IN3(n5423), .Q(n5412) );
  NAND2X0 U5408 ( .IN1(n5460), .IN2(n5461), .QN(n5423) );
  MUX21X1 U5409 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1488 ), .Q(n5461) );
  MUX21X1 U5410 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1489 ), .Q(n5460) );
  NAND2X0 U5411 ( .IN1(n5462), .IN2(n5463), .QN(n5424) );
  MUX21X1 U5412 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1491 ), .Q(n5463) );
  MUX21X1 U5413 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1490 ), .Q(n5462) );
  NAND2X0 U5414 ( .IN1(n5464), .IN2(n5465), .QN(n5426) );
  MUX21X1 U5415 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1486 ), .Q(n5465) );
  MUX21X1 U5416 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1487 ), .Q(n5464) );
  AOI22X1 U5417 ( .IN1(n5466), .IN2(n5467), .IN3(n5468), .IN4(n5469), .QN(
        n5413) );
  OR2X1 U5418 ( .IN1(n5467), .IN2(n5466), .Q(n5468) );
  XNOR3X1 U5419 ( .IN1(n5438), .IN2(n5439), .IN3(n5441), .Q(n5414) );
  NAND2X0 U5420 ( .IN1(n5470), .IN2(n5471), .QN(n5441) );
  MUX21X1 U5421 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1480 ), .Q(n5471) );
  MUX21X1 U5422 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1481 ), .Q(n5470) );
  NAND2X0 U5423 ( .IN1(n5472), .IN2(n5473), .QN(n5439) );
  MUX21X1 U5424 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1485 ), .Q(n5473) );
  MUX21X1 U5425 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1484 ), .Q(n5472) );
  NAND2X0 U5426 ( .IN1(n5474), .IN2(n5475), .QN(n5438) );
  MUX21X1 U5427 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1482 ), .Q(n5475) );
  MUX21X1 U5428 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1483 ), .Q(n5474) );
  XOR2X1 U5429 ( .IN1(n5363), .IN2(n5364), .Q(n5402) );
  NAND2X0 U5430 ( .IN1(n5476), .IN2(n5477), .QN(n5364) );
  MUX21X1 U5431 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1476 ), .Q(n5477) );
  MUX21X1 U5432 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1477 ), .Q(n5476) );
  NAND2X0 U5433 ( .IN1(n5478), .IN2(n5479), .QN(n5363) );
  MUX21X1 U5434 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1479 ), .Q(n5479) );
  MUX21X1 U5435 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1478 ), .Q(n5478) );
  XOR2X1 U5436 ( .IN1(n5403), .IN2(n5480), .Q(n5459) );
  NAND2X0 U5437 ( .IN1(n5406), .IN2(n5407), .QN(n5480) );
  AO22X1 U5438 ( .IN1(n5481), .IN2(n5482), .IN3(n5483), .IN4(n5484), .Q(n5403)
         );
  OR2X1 U5439 ( .IN1(n5482), .IN2(n5481), .Q(n5483) );
  AO22X1 U5440 ( .IN1(n5485), .IN2(n5486), .IN3(n5487), .IN4(n3491), .Q(
        \i_m4stg_frac/a1cout[23] ) );
  AO22X1 U5441 ( .IN1(n5488), .IN2(n5489), .IN3(n5490), .IN4(n5491), .Q(n3491)
         );
  OR2X1 U5442 ( .IN1(n5488), .IN2(n5489), .Q(n5491) );
  AND2X1 U5443 ( .IN1(n5492), .IN2(n5493), .Q(n5490) );
  NAND2X0 U5444 ( .IN1(n3492), .IN2(n3490), .QN(n5487) );
  INVX0 U5445 ( .INP(n5485), .ZN(n3490) );
  INVX0 U5446 ( .INP(n3492), .ZN(n5486) );
  MUX21X1 U5447 ( .IN1(n5494), .IN2(n5495), .S(n5496), .Q(n3492) );
  INVX0 U5448 ( .INP(n5497), .ZN(n5496) );
  XOR2X1 U5449 ( .IN1(n5454), .IN2(n5452), .Q(n5485) );
  OA22X1 U5450 ( .IN1(n5498), .IN2(n5499), .IN3(n5500), .IN4(n5501), .Q(n5452)
         );
  AND2X1 U5451 ( .IN1(n5499), .IN2(n5498), .Q(n5501) );
  XNOR3X1 U5452 ( .IN1(n5502), .IN2(n5445), .IN3(n5451), .Q(n5454) );
  XOR3X1 U5453 ( .IN1(n5457), .IN2(n5456), .IN3(n5455), .Q(n5451) );
  XNOR3X1 U5454 ( .IN1(n5469), .IN2(n5467), .IN3(n5466), .Q(n5455) );
  NAND2X0 U5455 ( .IN1(n5503), .IN2(n5504), .QN(n5466) );
  MUX21X1 U5456 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1487 ), .Q(n5504) );
  MUX21X1 U5457 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1488 ), .Q(n5503) );
  NAND2X0 U5458 ( .IN1(n5505), .IN2(n5506), .QN(n5467) );
  MUX21X1 U5459 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1490 ), .Q(n5506) );
  MUX21X1 U5460 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1489 ), .Q(n5505) );
  NAND2X0 U5461 ( .IN1(n5507), .IN2(n5508), .QN(n5469) );
  MUX21X1 U5462 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1485 ), .Q(n5508) );
  MUX21X1 U5463 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1486 ), .Q(n5507) );
  AOI22X1 U5464 ( .IN1(n5509), .IN2(n5510), .IN3(n5511), .IN4(n5512), .QN(
        n5456) );
  OR2X1 U5465 ( .IN1(n5510), .IN2(n5509), .Q(n5511) );
  XNOR3X1 U5466 ( .IN1(n5481), .IN2(n5482), .IN3(n5484), .Q(n5457) );
  NAND2X0 U5467 ( .IN1(n5513), .IN2(n5514), .QN(n5484) );
  MUX21X1 U5468 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1479 ), .Q(n5514) );
  MUX21X1 U5469 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1480 ), .Q(n5513) );
  NAND2X0 U5470 ( .IN1(n5515), .IN2(n5516), .QN(n5482) );
  MUX21X1 U5471 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1484 ), .Q(n5516) );
  MUX21X1 U5472 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1483 ), .Q(n5515) );
  NAND2X0 U5473 ( .IN1(n5517), .IN2(n5518), .QN(n5481) );
  MUX21X1 U5474 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1481 ), .Q(n5518) );
  MUX21X1 U5475 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1482 ), .Q(n5517) );
  XOR2X1 U5476 ( .IN1(n5406), .IN2(n5407), .Q(n5445) );
  NAND2X0 U5477 ( .IN1(n5519), .IN2(n5520), .QN(n5407) );
  MUX21X1 U5478 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1476 ), .Q(n5520) );
  MUX21X1 U5479 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1475 ), .Q(n5519) );
  NAND2X0 U5480 ( .IN1(n5521), .IN2(n5522), .QN(n5406) );
  MUX21X1 U5481 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1478 ), .Q(n5522) );
  MUX21X1 U5482 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1477 ), .Q(n5521) );
  XOR2X1 U5483 ( .IN1(n5446), .IN2(n5523), .Q(n5502) );
  NAND2X0 U5484 ( .IN1(n5449), .IN2(n5450), .QN(n5523) );
  AO22X1 U5485 ( .IN1(n5524), .IN2(n5525), .IN3(n5526), .IN4(n5527), .Q(n5446)
         );
  OR2X1 U5486 ( .IN1(n5525), .IN2(n5524), .Q(n5526) );
  AO22X1 U5487 ( .IN1(n5528), .IN2(n5529), .IN3(n5530), .IN4(n3494), .Q(
        \i_m4stg_frac/a1cout[22] ) );
  AO22X1 U5488 ( .IN1(n5531), .IN2(n5532), .IN3(n5533), .IN4(n5534), .Q(n3494)
         );
  OR2X1 U5489 ( .IN1(n5531), .IN2(n5532), .Q(n5534) );
  AND2X1 U5490 ( .IN1(n5535), .IN2(n5536), .Q(n5533) );
  NAND2X0 U5491 ( .IN1(n3495), .IN2(n3493), .QN(n5530) );
  INVX0 U5492 ( .INP(n5528), .ZN(n3493) );
  INVX0 U5493 ( .INP(n3495), .ZN(n5529) );
  MUX21X1 U5494 ( .IN1(n5537), .IN2(n5538), .S(n5539), .Q(n3495) );
  INVX0 U5495 ( .INP(n5540), .ZN(n5539) );
  XOR2X1 U5496 ( .IN1(n5497), .IN2(n5495), .Q(n5528) );
  OA22X1 U5497 ( .IN1(n5541), .IN2(n5542), .IN3(n5543), .IN4(n5544), .Q(n5495)
         );
  AND2X1 U5498 ( .IN1(n5542), .IN2(n5541), .Q(n5544) );
  XNOR3X1 U5499 ( .IN1(n5545), .IN2(n5488), .IN3(n5494), .Q(n5497) );
  XOR3X1 U5500 ( .IN1(n5500), .IN2(n5499), .IN3(n5498), .Q(n5494) );
  XNOR3X1 U5501 ( .IN1(n5512), .IN2(n5510), .IN3(n5509), .Q(n5498) );
  NAND2X0 U5502 ( .IN1(n5546), .IN2(n5547), .QN(n5509) );
  MUX21X1 U5503 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1486 ), .Q(n5547) );
  MUX21X1 U5504 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1487 ), .Q(n5546) );
  NAND2X0 U5505 ( .IN1(n5548), .IN2(n5549), .QN(n5510) );
  MUX21X1 U5506 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1489 ), .Q(n5549) );
  MUX21X1 U5507 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1488 ), .Q(n5548) );
  NAND2X0 U5508 ( .IN1(n5550), .IN2(n5551), .QN(n5512) );
  MUX21X1 U5509 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1484 ), .Q(n5551) );
  MUX21X1 U5510 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1485 ), .Q(n5550) );
  AOI22X1 U5511 ( .IN1(n5552), .IN2(n5553), .IN3(n5554), .IN4(n5555), .QN(
        n5499) );
  OR2X1 U5512 ( .IN1(n5553), .IN2(n5552), .Q(n5554) );
  XNOR3X1 U5513 ( .IN1(n5524), .IN2(n5525), .IN3(n5527), .Q(n5500) );
  NAND2X0 U5514 ( .IN1(n5556), .IN2(n5557), .QN(n5527) );
  MUX21X1 U5515 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1478 ), .Q(n5557) );
  MUX21X1 U5516 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1479 ), .Q(n5556) );
  NAND2X0 U5517 ( .IN1(n5558), .IN2(n5559), .QN(n5525) );
  MUX21X1 U5518 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1483 ), .Q(n5559) );
  MUX21X1 U5519 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1482 ), .Q(n5558) );
  NAND2X0 U5520 ( .IN1(n5560), .IN2(n5561), .QN(n5524) );
  MUX21X1 U5521 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1480 ), .Q(n5561) );
  MUX21X1 U5522 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1481 ), .Q(n5560) );
  XOR2X1 U5523 ( .IN1(n5449), .IN2(n5450), .Q(n5488) );
  NAND2X0 U5524 ( .IN1(n5562), .IN2(n5563), .QN(n5450) );
  MUX21X1 U5525 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1475 ), .Q(n5563) );
  MUX21X1 U5526 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1474 ), .Q(n5562) );
  NAND2X0 U5527 ( .IN1(n5564), .IN2(n5565), .QN(n5449) );
  MUX21X1 U5528 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1477 ), .Q(n5565) );
  MUX21X1 U5529 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1476 ), .Q(n5564) );
  XOR2X1 U5530 ( .IN1(n5489), .IN2(n5566), .Q(n5545) );
  NAND2X0 U5531 ( .IN1(n5492), .IN2(n5493), .QN(n5566) );
  AO22X1 U5532 ( .IN1(n5567), .IN2(n5568), .IN3(n5569), .IN4(n5570), .Q(n5489)
         );
  OR2X1 U5533 ( .IN1(n5568), .IN2(n5567), .Q(n5569) );
  AO22X1 U5534 ( .IN1(n5571), .IN2(n5572), .IN3(n5573), .IN4(n3497), .Q(
        \i_m4stg_frac/a1cout[21] ) );
  AO22X1 U5535 ( .IN1(n5574), .IN2(n5575), .IN3(n5576), .IN4(n5577), .Q(n3497)
         );
  OR2X1 U5536 ( .IN1(n5574), .IN2(n5575), .Q(n5577) );
  AND2X1 U5537 ( .IN1(n5578), .IN2(n5579), .Q(n5576) );
  NAND2X0 U5538 ( .IN1(n3498), .IN2(n3496), .QN(n5573) );
  INVX0 U5539 ( .INP(n5571), .ZN(n3496) );
  INVX0 U5540 ( .INP(n3498), .ZN(n5572) );
  MUX21X1 U5541 ( .IN1(n5580), .IN2(n5581), .S(n5582), .Q(n3498) );
  INVX0 U5542 ( .INP(n5583), .ZN(n5582) );
  XOR2X1 U5543 ( .IN1(n5540), .IN2(n5538), .Q(n5571) );
  OA22X1 U5544 ( .IN1(n5584), .IN2(n5585), .IN3(n5586), .IN4(n5587), .Q(n5538)
         );
  AND2X1 U5545 ( .IN1(n5585), .IN2(n5584), .Q(n5587) );
  XNOR3X1 U5546 ( .IN1(n5588), .IN2(n5531), .IN3(n5537), .Q(n5540) );
  XOR3X1 U5547 ( .IN1(n5543), .IN2(n5542), .IN3(n5541), .Q(n5537) );
  XNOR3X1 U5548 ( .IN1(n5555), .IN2(n5553), .IN3(n5552), .Q(n5541) );
  NAND2X0 U5549 ( .IN1(n5589), .IN2(n5590), .QN(n5552) );
  MUX21X1 U5550 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1485 ), .Q(n5590) );
  MUX21X1 U5551 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1486 ), .Q(n5589) );
  NAND2X0 U5552 ( .IN1(n5591), .IN2(n5592), .QN(n5553) );
  MUX21X1 U5553 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1488 ), .Q(n5592) );
  MUX21X1 U5554 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1487 ), .Q(n5591) );
  NAND2X0 U5555 ( .IN1(n5593), .IN2(n5594), .QN(n5555) );
  MUX21X1 U5556 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1483 ), .Q(n5594) );
  MUX21X1 U5557 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1484 ), .Q(n5593) );
  AOI22X1 U5558 ( .IN1(n5595), .IN2(n5596), .IN3(n5597), .IN4(n5598), .QN(
        n5542) );
  OR2X1 U5559 ( .IN1(n5596), .IN2(n5595), .Q(n5597) );
  XNOR3X1 U5560 ( .IN1(n5567), .IN2(n5568), .IN3(n5570), .Q(n5543) );
  NAND2X0 U5561 ( .IN1(n5599), .IN2(n5600), .QN(n5570) );
  MUX21X1 U5562 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1477 ), .Q(n5600) );
  MUX21X1 U5563 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1478 ), .Q(n5599) );
  NAND2X0 U5564 ( .IN1(n5601), .IN2(n5602), .QN(n5568) );
  MUX21X1 U5565 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1482 ), .Q(n5602) );
  MUX21X1 U5566 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1481 ), .Q(n5601) );
  NAND2X0 U5567 ( .IN1(n5603), .IN2(n5604), .QN(n5567) );
  MUX21X1 U5568 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1479 ), .Q(n5604) );
  MUX21X1 U5569 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1480 ), .Q(n5603) );
  XOR2X1 U5570 ( .IN1(n5492), .IN2(n5493), .Q(n5531) );
  NAND2X0 U5571 ( .IN1(n5605), .IN2(n5606), .QN(n5493) );
  MUX21X1 U5572 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1473 ), .Q(n5606) );
  MUX21X1 U5573 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1474 ), .Q(n5605) );
  NAND2X0 U5574 ( .IN1(n5607), .IN2(n5608), .QN(n5492) );
  MUX21X1 U5575 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1476 ), .Q(n5608) );
  MUX21X1 U5576 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1475 ), .Q(n5607) );
  XOR2X1 U5577 ( .IN1(n5532), .IN2(n5609), .Q(n5588) );
  NAND2X0 U5578 ( .IN1(n5535), .IN2(n5536), .QN(n5609) );
  AO22X1 U5579 ( .IN1(n5610), .IN2(n5611), .IN3(n5612), .IN4(n5613), .Q(n5532)
         );
  OR2X1 U5580 ( .IN1(n5611), .IN2(n5610), .Q(n5612) );
  AO22X1 U5581 ( .IN1(n5614), .IN2(n5615), .IN3(n5616), .IN4(n3500), .Q(
        \i_m4stg_frac/a1cout[20] ) );
  AO22X1 U5582 ( .IN1(n5617), .IN2(n5618), .IN3(n5619), .IN4(n5620), .Q(n3500)
         );
  OR2X1 U5583 ( .IN1(n5617), .IN2(n5618), .Q(n5620) );
  AND2X1 U5584 ( .IN1(n5621), .IN2(n5622), .Q(n5619) );
  NAND2X0 U5585 ( .IN1(n3501), .IN2(n3499), .QN(n5616) );
  INVX0 U5586 ( .INP(n5614), .ZN(n3499) );
  INVX0 U5587 ( .INP(n3501), .ZN(n5615) );
  MUX21X1 U5588 ( .IN1(n5623), .IN2(n5624), .S(n5625), .Q(n3501) );
  INVX0 U5589 ( .INP(n5626), .ZN(n5625) );
  XOR2X1 U5590 ( .IN1(n5583), .IN2(n5581), .Q(n5614) );
  OA22X1 U5591 ( .IN1(n5627), .IN2(n5628), .IN3(n5629), .IN4(n5630), .Q(n5581)
         );
  AND2X1 U5592 ( .IN1(n5628), .IN2(n5627), .Q(n5630) );
  XNOR3X1 U5593 ( .IN1(n5631), .IN2(n5574), .IN3(n5580), .Q(n5583) );
  XOR3X1 U5594 ( .IN1(n5586), .IN2(n5585), .IN3(n5584), .Q(n5580) );
  XNOR3X1 U5595 ( .IN1(n5598), .IN2(n5596), .IN3(n5595), .Q(n5584) );
  NAND2X0 U5596 ( .IN1(n5632), .IN2(n5633), .QN(n5595) );
  MUX21X1 U5597 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1484 ), .Q(n5633) );
  MUX21X1 U5598 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1485 ), .Q(n5632) );
  NAND2X0 U5599 ( .IN1(n5634), .IN2(n5635), .QN(n5596) );
  MUX21X1 U5600 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1487 ), .Q(n5635) );
  MUX21X1 U5601 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1486 ), .Q(n5634) );
  NAND2X0 U5602 ( .IN1(n5636), .IN2(n5637), .QN(n5598) );
  MUX21X1 U5603 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1482 ), .Q(n5637) );
  MUX21X1 U5604 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1483 ), .Q(n5636) );
  AOI22X1 U5605 ( .IN1(n5638), .IN2(n5639), .IN3(n5640), .IN4(n5641), .QN(
        n5585) );
  OR2X1 U5606 ( .IN1(n5639), .IN2(n5638), .Q(n5640) );
  XNOR3X1 U5607 ( .IN1(n5610), .IN2(n5611), .IN3(n5613), .Q(n5586) );
  NAND2X0 U5608 ( .IN1(n5642), .IN2(n5643), .QN(n5613) );
  MUX21X1 U5609 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1476 ), .Q(n5643) );
  MUX21X1 U5610 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1477 ), .Q(n5642) );
  NAND2X0 U5611 ( .IN1(n5644), .IN2(n5645), .QN(n5611) );
  MUX21X1 U5612 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1481 ), .Q(n5645) );
  MUX21X1 U5613 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1480 ), .Q(n5644) );
  NAND2X0 U5614 ( .IN1(n5646), .IN2(n5647), .QN(n5610) );
  MUX21X1 U5615 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1478 ), .Q(n5647) );
  MUX21X1 U5616 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1479 ), .Q(n5646) );
  XOR2X1 U5617 ( .IN1(n5535), .IN2(n5536), .Q(n5574) );
  NAND2X0 U5618 ( .IN1(n5648), .IN2(n5649), .QN(n5536) );
  MUX21X1 U5619 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1473 ), .Q(n5649) );
  MUX21X1 U5620 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1472 ), .Q(n5648) );
  NAND2X0 U5621 ( .IN1(n5650), .IN2(n5651), .QN(n5535) );
  MUX21X1 U5622 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1474 ), .Q(n5651) );
  MUX21X1 U5623 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1475 ), .Q(n5650) );
  XOR2X1 U5624 ( .IN1(n5575), .IN2(n5652), .Q(n5631) );
  NAND2X0 U5625 ( .IN1(n5578), .IN2(n5579), .QN(n5652) );
  AO22X1 U5626 ( .IN1(n5653), .IN2(n5654), .IN3(n5655), .IN4(n5656), .Q(n5575)
         );
  OR2X1 U5627 ( .IN1(n5654), .IN2(n5653), .Q(n5655) );
  AO22X1 U5628 ( .IN1(n5657), .IN2(n5658), .IN3(n5659), .IN4(n3508), .Q(
        \i_m4stg_frac/a1cout[19] ) );
  AO22X1 U5629 ( .IN1(n5660), .IN2(n5661), .IN3(n5662), .IN4(n5663), .Q(n3508)
         );
  OR2X1 U5630 ( .IN1(n5660), .IN2(n5661), .Q(n5663) );
  AND2X1 U5631 ( .IN1(n5664), .IN2(n5665), .Q(n5662) );
  NAND2X0 U5632 ( .IN1(n3509), .IN2(n3507), .QN(n5659) );
  INVX0 U5633 ( .INP(n5657), .ZN(n3507) );
  INVX0 U5634 ( .INP(n3509), .ZN(n5658) );
  MUX21X1 U5635 ( .IN1(n5666), .IN2(n5667), .S(n5668), .Q(n3509) );
  INVX0 U5636 ( .INP(n5669), .ZN(n5668) );
  XOR2X1 U5637 ( .IN1(n5626), .IN2(n5624), .Q(n5657) );
  OA22X1 U5638 ( .IN1(n5670), .IN2(n5671), .IN3(n5672), .IN4(n5673), .Q(n5624)
         );
  AND2X1 U5639 ( .IN1(n5671), .IN2(n5670), .Q(n5673) );
  XNOR3X1 U5640 ( .IN1(n5674), .IN2(n5617), .IN3(n5623), .Q(n5626) );
  XOR3X1 U5641 ( .IN1(n5629), .IN2(n5628), .IN3(n5627), .Q(n5623) );
  XNOR3X1 U5642 ( .IN1(n5641), .IN2(n5639), .IN3(n5638), .Q(n5627) );
  NAND2X0 U5643 ( .IN1(n5675), .IN2(n5676), .QN(n5638) );
  MUX21X1 U5644 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1483 ), .Q(n5676) );
  MUX21X1 U5645 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1484 ), .Q(n5675) );
  NAND2X0 U5646 ( .IN1(n5677), .IN2(n5678), .QN(n5639) );
  MUX21X1 U5647 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1486 ), .Q(n5678) );
  MUX21X1 U5648 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1485 ), .Q(n5677) );
  NAND2X0 U5649 ( .IN1(n5679), .IN2(n5680), .QN(n5641) );
  MUX21X1 U5650 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1481 ), .Q(n5680) );
  MUX21X1 U5651 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1482 ), .Q(n5679) );
  AOI22X1 U5652 ( .IN1(n5681), .IN2(n5682), .IN3(n5683), .IN4(n5684), .QN(
        n5628) );
  OR2X1 U5653 ( .IN1(n5682), .IN2(n5681), .Q(n5683) );
  XNOR3X1 U5654 ( .IN1(n5653), .IN2(n5654), .IN3(n5656), .Q(n5629) );
  NAND2X0 U5655 ( .IN1(n5685), .IN2(n5686), .QN(n5656) );
  MUX21X1 U5656 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1475 ), .Q(n5686) );
  MUX21X1 U5657 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1476 ), .Q(n5685) );
  NAND2X0 U5658 ( .IN1(n5687), .IN2(n5688), .QN(n5654) );
  MUX21X1 U5659 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1480 ), .Q(n5688) );
  MUX21X1 U5660 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1479 ), .Q(n5687) );
  NAND2X0 U5661 ( .IN1(n5689), .IN2(n5690), .QN(n5653) );
  MUX21X1 U5662 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1477 ), .Q(n5690) );
  MUX21X1 U5663 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1478 ), .Q(n5689) );
  XOR2X1 U5664 ( .IN1(n5578), .IN2(n5579), .Q(n5617) );
  NAND2X0 U5665 ( .IN1(n5691), .IN2(n5692), .QN(n5579) );
  MUX21X1 U5666 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1471 ), .Q(n5692) );
  MUX21X1 U5667 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1472 ), .Q(n5691) );
  NAND2X0 U5668 ( .IN1(n5693), .IN2(n5694), .QN(n5578) );
  MUX21X1 U5669 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1474 ), .Q(n5694) );
  MUX21X1 U5670 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1473 ), .Q(n5693) );
  XOR2X1 U5671 ( .IN1(n5618), .IN2(n5695), .Q(n5674) );
  NAND2X0 U5672 ( .IN1(n5621), .IN2(n5622), .QN(n5695) );
  AO22X1 U5673 ( .IN1(n5696), .IN2(n5697), .IN3(n5698), .IN4(n5699), .Q(n5618)
         );
  OR2X1 U5674 ( .IN1(n5697), .IN2(n5696), .Q(n5698) );
  AO22X1 U5675 ( .IN1(n5700), .IN2(n5701), .IN3(n5702), .IN4(n3511), .Q(
        \i_m4stg_frac/a1cout[18] ) );
  AO22X1 U5676 ( .IN1(n5703), .IN2(n5704), .IN3(n5705), .IN4(n5706), .Q(n3511)
         );
  OR2X1 U5677 ( .IN1(n5703), .IN2(n5704), .Q(n5706) );
  AND2X1 U5678 ( .IN1(n5707), .IN2(n5708), .Q(n5705) );
  NAND2X0 U5679 ( .IN1(n3512), .IN2(n3510), .QN(n5702) );
  INVX0 U5680 ( .INP(n5700), .ZN(n3510) );
  INVX0 U5681 ( .INP(n3512), .ZN(n5701) );
  MUX21X1 U5682 ( .IN1(n5709), .IN2(n5710), .S(n5711), .Q(n3512) );
  INVX0 U5683 ( .INP(n5712), .ZN(n5711) );
  XOR2X1 U5684 ( .IN1(n5669), .IN2(n5667), .Q(n5700) );
  OA22X1 U5685 ( .IN1(n5713), .IN2(n5714), .IN3(n5715), .IN4(n5716), .Q(n5667)
         );
  AND2X1 U5686 ( .IN1(n5714), .IN2(n5713), .Q(n5716) );
  XNOR3X1 U5687 ( .IN1(n5717), .IN2(n5660), .IN3(n5666), .Q(n5669) );
  XOR3X1 U5688 ( .IN1(n5672), .IN2(n5671), .IN3(n5670), .Q(n5666) );
  XNOR3X1 U5689 ( .IN1(n5684), .IN2(n5682), .IN3(n5681), .Q(n5670) );
  NAND2X0 U5690 ( .IN1(n5718), .IN2(n5719), .QN(n5681) );
  MUX21X1 U5691 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1482 ), .Q(n5719) );
  MUX21X1 U5692 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1483 ), .Q(n5718) );
  NAND2X0 U5693 ( .IN1(n5720), .IN2(n5721), .QN(n5682) );
  MUX21X1 U5694 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1485 ), .Q(n5721) );
  MUX21X1 U5695 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1484 ), .Q(n5720) );
  NAND2X0 U5696 ( .IN1(n5722), .IN2(n5723), .QN(n5684) );
  MUX21X1 U5697 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1480 ), .Q(n5723) );
  MUX21X1 U5698 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1481 ), .Q(n5722) );
  AOI22X1 U5699 ( .IN1(n5724), .IN2(n5725), .IN3(n5726), .IN4(n5727), .QN(
        n5671) );
  OR2X1 U5700 ( .IN1(n5725), .IN2(n5724), .Q(n5726) );
  XNOR3X1 U5701 ( .IN1(n5696), .IN2(n5697), .IN3(n5699), .Q(n5672) );
  NAND2X0 U5702 ( .IN1(n5728), .IN2(n5729), .QN(n5699) );
  MUX21X1 U5703 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1474 ), .Q(n5729) );
  MUX21X1 U5704 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1475 ), .Q(n5728) );
  NAND2X0 U5705 ( .IN1(n5730), .IN2(n5731), .QN(n5697) );
  MUX21X1 U5706 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1479 ), .Q(n5731) );
  MUX21X1 U5707 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1478 ), .Q(n5730) );
  NAND2X0 U5708 ( .IN1(n5732), .IN2(n5733), .QN(n5696) );
  MUX21X1 U5709 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1476 ), .Q(n5733) );
  MUX21X1 U5710 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1477 ), .Q(n5732) );
  XOR2X1 U5711 ( .IN1(n5621), .IN2(n5622), .Q(n5660) );
  NAND2X0 U5712 ( .IN1(n5734), .IN2(n5735), .QN(n5622) );
  MUX21X1 U5713 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1470 ), .Q(n5735) );
  MUX21X1 U5714 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1471 ), .Q(n5734) );
  NAND2X0 U5715 ( .IN1(n5736), .IN2(n5737), .QN(n5621) );
  MUX21X1 U5716 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1473 ), .Q(n5737) );
  MUX21X1 U5717 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1472 ), .Q(n5736) );
  XOR2X1 U5718 ( .IN1(n5661), .IN2(n5738), .Q(n5717) );
  NAND2X0 U5719 ( .IN1(n5664), .IN2(n5665), .QN(n5738) );
  AO22X1 U5720 ( .IN1(n5739), .IN2(n5740), .IN3(n5741), .IN4(n5742), .Q(n5661)
         );
  OR2X1 U5721 ( .IN1(n5740), .IN2(n5739), .Q(n5741) );
  AO22X1 U5722 ( .IN1(n5743), .IN2(n5744), .IN3(n5745), .IN4(n3514), .Q(
        \i_m4stg_frac/a1cout[17] ) );
  AO22X1 U5723 ( .IN1(n5746), .IN2(n5747), .IN3(n5748), .IN4(n5749), .Q(n3514)
         );
  OR2X1 U5724 ( .IN1(n5746), .IN2(n5747), .Q(n5749) );
  NAND2X0 U5725 ( .IN1(n3515), .IN2(n3513), .QN(n5745) );
  INVX0 U5726 ( .INP(n5743), .ZN(n3513) );
  INVX0 U5727 ( .INP(n3515), .ZN(n5744) );
  MUX21X1 U5728 ( .IN1(n5750), .IN2(n5751), .S(n5752), .Q(n3515) );
  INVX0 U5729 ( .INP(n5753), .ZN(n5752) );
  XOR2X1 U5730 ( .IN1(n5712), .IN2(n5710), .Q(n5743) );
  OA22X1 U5731 ( .IN1(n5754), .IN2(n5755), .IN3(n5756), .IN4(n5757), .Q(n5710)
         );
  AND2X1 U5732 ( .IN1(n5755), .IN2(n5754), .Q(n5757) );
  XNOR3X1 U5733 ( .IN1(n5758), .IN2(n5703), .IN3(n5709), .Q(n5712) );
  XOR3X1 U5734 ( .IN1(n5715), .IN2(n5714), .IN3(n5713), .Q(n5709) );
  XNOR3X1 U5735 ( .IN1(n5727), .IN2(n5725), .IN3(n5724), .Q(n5713) );
  NAND2X0 U5736 ( .IN1(n5759), .IN2(n5760), .QN(n5724) );
  MUX21X1 U5737 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1481 ), .Q(n5760) );
  MUX21X1 U5738 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1482 ), .Q(n5759) );
  NAND2X0 U5739 ( .IN1(n5761), .IN2(n5762), .QN(n5725) );
  MUX21X1 U5740 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1484 ), .Q(n5762) );
  MUX21X1 U5741 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1483 ), .Q(n5761) );
  NAND2X0 U5742 ( .IN1(n5763), .IN2(n5764), .QN(n5727) );
  MUX21X1 U5743 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1479 ), .Q(n5764) );
  MUX21X1 U5744 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1480 ), .Q(n5763) );
  AOI22X1 U5745 ( .IN1(n5765), .IN2(n5766), .IN3(n5767), .IN4(n5768), .QN(
        n5714) );
  OR2X1 U5746 ( .IN1(n5766), .IN2(n5765), .Q(n5767) );
  XNOR3X1 U5747 ( .IN1(n5739), .IN2(n5740), .IN3(n5742), .Q(n5715) );
  NAND2X0 U5748 ( .IN1(n5769), .IN2(n5770), .QN(n5742) );
  MUX21X1 U5749 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1474 ), .Q(n5770) );
  MUX21X1 U5750 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1473 ), .Q(n5769) );
  NAND2X0 U5751 ( .IN1(n5771), .IN2(n5772), .QN(n5740) );
  MUX21X1 U5752 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1478 ), .Q(n5772) );
  MUX21X1 U5753 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1477 ), .Q(n5771) );
  NAND2X0 U5754 ( .IN1(n5773), .IN2(n5774), .QN(n5739) );
  MUX21X1 U5755 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1475 ), .Q(n5774) );
  MUX21X1 U5756 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1476 ), .Q(n5773) );
  XOR2X1 U5757 ( .IN1(n5664), .IN2(n5665), .Q(n5703) );
  NAND2X0 U5758 ( .IN1(n5775), .IN2(n5776), .QN(n5665) );
  MUX21X1 U5759 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1469 ), .Q(n5776) );
  MUX21X1 U5760 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1470 ), .Q(n5775) );
  NAND2X0 U5761 ( .IN1(n5777), .IN2(n5778), .QN(n5664) );
  MUX21X1 U5762 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1472 ), .Q(n5778) );
  MUX21X1 U5763 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1471 ), .Q(n5777) );
  XOR2X1 U5764 ( .IN1(n5704), .IN2(n5779), .Q(n5758) );
  NAND2X0 U5765 ( .IN1(n5707), .IN2(n5708), .QN(n5779) );
  AO22X1 U5766 ( .IN1(n5780), .IN2(n5781), .IN3(n5782), .IN4(n5783), .Q(n5704)
         );
  OR2X1 U5767 ( .IN1(n5781), .IN2(n5780), .Q(n5782) );
  AO22X1 U5768 ( .IN1(n3517), .IN2(n3518), .IN3(n5784), .IN4(n3516), .Q(
        \i_m4stg_frac/a1cout[16] ) );
  AO22X1 U5769 ( .IN1(n5785), .IN2(n5786), .IN3(n5787), .IN4(n5788), .Q(n3516)
         );
  OR2X1 U5770 ( .IN1(n5785), .IN2(n5786), .Q(n5788) );
  OR2X1 U5771 ( .IN1(n3518), .IN2(n3517), .Q(n5784) );
  INVX0 U5772 ( .INP(n5789), .ZN(n3518) );
  MUX21X1 U5773 ( .IN1(n5790), .IN2(n5791), .S(n5792), .Q(n5789) );
  INVX0 U5774 ( .INP(n5793), .ZN(n5792) );
  XNOR2X1 U5775 ( .IN1(n5753), .IN2(n5750), .Q(n3517) );
  OA22X1 U5776 ( .IN1(n5794), .IN2(n5795), .IN3(n5796), .IN4(n5797), .Q(n5750)
         );
  AND2X1 U5777 ( .IN1(n5795), .IN2(n5794), .Q(n5797) );
  XNOR3X1 U5778 ( .IN1(n5798), .IN2(n5748), .IN3(n5751), .Q(n5753) );
  XOR3X1 U5779 ( .IN1(n5756), .IN2(n5755), .IN3(n5754), .Q(n5751) );
  XNOR3X1 U5780 ( .IN1(n5768), .IN2(n5766), .IN3(n5765), .Q(n5754) );
  NAND2X0 U5781 ( .IN1(n5799), .IN2(n5800), .QN(n5765) );
  MUX21X1 U5782 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1480 ), .Q(n5800) );
  MUX21X1 U5783 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1481 ), .Q(n5799) );
  NAND2X0 U5784 ( .IN1(n5801), .IN2(n5802), .QN(n5766) );
  MUX21X1 U5785 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1483 ), .Q(n5802) );
  MUX21X1 U5786 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1482 ), .Q(n5801) );
  NAND2X0 U5787 ( .IN1(n5803), .IN2(n5804), .QN(n5768) );
  MUX21X1 U5788 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1478 ), .Q(n5804) );
  MUX21X1 U5789 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1479 ), .Q(n5803) );
  AOI22X1 U5790 ( .IN1(n5805), .IN2(n5806), .IN3(n5807), .IN4(n5808), .QN(
        n5755) );
  OR2X1 U5791 ( .IN1(n5806), .IN2(n5805), .Q(n5807) );
  XNOR3X1 U5792 ( .IN1(n5780), .IN2(n5781), .IN3(n5783), .Q(n5756) );
  NAND2X0 U5793 ( .IN1(n5809), .IN2(n5810), .QN(n5783) );
  MUX21X1 U5794 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1472 ), .Q(n5810) );
  MUX21X1 U5795 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1473 ), .Q(n5809) );
  NAND2X0 U5796 ( .IN1(n5811), .IN2(n5812), .QN(n5781) );
  MUX21X1 U5797 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1477 ), .Q(n5812) );
  MUX21X1 U5798 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1476 ), .Q(n5811) );
  NAND2X0 U5799 ( .IN1(n5813), .IN2(n5814), .QN(n5780) );
  MUX21X1 U5800 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1474 ), .Q(n5814) );
  MUX21X1 U5801 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1475 ), .Q(n5813) );
  XOR2X1 U5802 ( .IN1(n5708), .IN2(n5707), .Q(n5748) );
  NAND2X0 U5803 ( .IN1(n5815), .IN2(n5816), .QN(n5707) );
  MUX21X1 U5804 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1468 ), .Q(n5816) );
  MUX21X1 U5805 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1469 ), .Q(n5815) );
  NAND2X0 U5806 ( .IN1(n5817), .IN2(n5818), .QN(n5708) );
  MUX21X1 U5807 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1471 ), .Q(n5818) );
  MUX21X1 U5808 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1470 ), .Q(n5817) );
  XOR2X1 U5809 ( .IN1(n5747), .IN2(n5746), .Q(n5798) );
  AO22X1 U5810 ( .IN1(n5819), .IN2(n5820), .IN3(n5821), .IN4(n5822), .Q(n5746)
         );
  OR2X1 U5811 ( .IN1(n5819), .IN2(n5820), .Q(n5821) );
  AO22X1 U5812 ( .IN1(n5823), .IN2(n5824), .IN3(n5825), .IN4(n5826), .Q(n5747)
         );
  OR2X1 U5813 ( .IN1(n5824), .IN2(n5823), .Q(n5826) );
  AO22X1 U5814 ( .IN1(n3520), .IN2(n3521), .IN3(n5827), .IN4(n3519), .Q(
        \i_m4stg_frac/a1cout[15] ) );
  AO22X1 U5815 ( .IN1(n5828), .IN2(n5829), .IN3(n5830), .IN4(n5831), .Q(n3519)
         );
  OR2X1 U5816 ( .IN1(n5829), .IN2(n5828), .Q(n5831) );
  INVX0 U5817 ( .INP(n5832), .ZN(n5830) );
  OR2X1 U5818 ( .IN1(n3521), .IN2(n3520), .Q(n5827) );
  MUX21X1 U5819 ( .IN1(n5833), .IN2(n5834), .S(n5835), .Q(n3521) );
  XNOR2X1 U5820 ( .IN1(n5793), .IN2(n5790), .Q(n3520) );
  AOI22X1 U5821 ( .IN1(n5836), .IN2(n5837), .IN3(n5838), .IN4(n5839), .QN(
        n5790) );
  OR2X1 U5822 ( .IN1(n5837), .IN2(n5836), .Q(n5839) );
  XNOR3X1 U5823 ( .IN1(n5840), .IN2(n5787), .IN3(n5791), .Q(n5793) );
  XOR3X1 U5824 ( .IN1(n5796), .IN2(n5795), .IN3(n5794), .Q(n5791) );
  XNOR3X1 U5825 ( .IN1(n5808), .IN2(n5806), .IN3(n5805), .Q(n5794) );
  NAND2X0 U5826 ( .IN1(n5841), .IN2(n5842), .QN(n5805) );
  MUX21X1 U5827 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1479 ), .Q(n5842) );
  MUX21X1 U5828 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1480 ), .Q(n5841) );
  NAND2X0 U5829 ( .IN1(n5843), .IN2(n5844), .QN(n5806) );
  MUX21X1 U5830 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1482 ), .Q(n5844) );
  MUX21X1 U5831 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1481 ), .Q(n5843) );
  NAND2X0 U5832 ( .IN1(n5845), .IN2(n5846), .QN(n5808) );
  MUX21X1 U5833 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1477 ), .Q(n5846) );
  MUX21X1 U5834 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1478 ), .Q(n5845) );
  AOI22X1 U5835 ( .IN1(n5847), .IN2(n5848), .IN3(n5849), .IN4(n5850), .QN(
        n5795) );
  OR2X1 U5836 ( .IN1(n5848), .IN2(n5847), .Q(n5849) );
  XNOR3X1 U5837 ( .IN1(n5819), .IN2(n5820), .IN3(n5822), .Q(n5796) );
  NAND2X0 U5838 ( .IN1(n5851), .IN2(n5852), .QN(n5822) );
  MUX21X1 U5839 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1472 ), .Q(n5852) );
  MUX21X1 U5840 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1471 ), .Q(n5851) );
  NAND2X0 U5841 ( .IN1(n5853), .IN2(n5854), .QN(n5820) );
  MUX21X1 U5842 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1476 ), .Q(n5854) );
  MUX21X1 U5843 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1475 ), .Q(n5853) );
  NAND2X0 U5844 ( .IN1(n5855), .IN2(n5856), .QN(n5819) );
  MUX21X1 U5845 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1474 ), .Q(n5856) );
  MUX21X1 U5846 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1473 ), .Q(n5855) );
  XOR3X1 U5847 ( .IN1(n5825), .IN2(n5824), .IN3(n5823), .Q(n5787) );
  NAND2X0 U5848 ( .IN1(n5857), .IN2(n5858), .QN(n5823) );
  MUX21X1 U5849 ( .IN1(n3817), .IN2(n3818), .S(\i_m4stg_frac/n1470 ), .Q(n5858) );
  MUX21X1 U5850 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1469 ), .Q(n5857) );
  NAND2X0 U5851 ( .IN1(n5859), .IN2(n5860), .QN(n5824) );
  MUX21X1 U5852 ( .IN1(n3609), .IN2(n3759), .S(\i_m4stg_frac/n1468 ), .Q(n5860) );
  MUX21X1 U5853 ( .IN1(n3741), .IN2(n3742), .S(\i_m4stg_frac/n1467 ), .Q(n5859) );
  INVX0 U5854 ( .INP(n3741), .ZN(n5825) );
  XOR2X1 U5855 ( .IN1(n5786), .IN2(n5785), .Q(n5840) );
  AO22X1 U5856 ( .IN1(n5861), .IN2(n5862), .IN3(n5863), .IN4(n5864), .Q(n5785)
         );
  OR2X1 U5857 ( .IN1(n5861), .IN2(n5862), .Q(n5863) );
  OAI22X1 U5858 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(n3609), .IN3(n5865), .IN4(
        n5866), .QN(n5786) );
  OA21X1 U5859 ( .IN1(n1034), .IN2(n3759), .IN3(n3609), .Q(n5866) );
  AO22X1 U5860 ( .IN1(n5867), .IN2(n5868), .IN3(n5869), .IN4(n3523), .Q(
        \i_m4stg_frac/a1cout[14] ) );
  AO22X1 U5861 ( .IN1(n5870), .IN2(n5871), .IN3(n5872), .IN4(n5873), .Q(n3523)
         );
  OR2X1 U5862 ( .IN1(n5871), .IN2(n5870), .Q(n5873) );
  NAND2X0 U5863 ( .IN1(n3524), .IN2(n3522), .QN(n5869) );
  INVX0 U5864 ( .INP(n5867), .ZN(n3522) );
  INVX0 U5865 ( .INP(n3524), .ZN(n5868) );
  MUX21X1 U5866 ( .IN1(n5874), .IN2(n5875), .S(n5876), .Q(n3524) );
  INVX0 U5867 ( .INP(n5877), .ZN(n5876) );
  XNOR2X1 U5868 ( .IN1(n5835), .IN2(n5833), .Q(n5867) );
  XOR3X1 U5869 ( .IN1(n5878), .IN2(n5828), .IN3(n5834), .Q(n5835) );
  XOR3X1 U5870 ( .IN1(n5837), .IN2(n5836), .IN3(n5838), .Q(n5834) );
  XOR3X1 U5871 ( .IN1(n5861), .IN2(n5862), .IN3(n5864), .Q(n5838) );
  NAND2X0 U5872 ( .IN1(n5879), .IN2(n5880), .QN(n5864) );
  MUX21X1 U5873 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1470 ), .Q(n5880) );
  MUX21X1 U5874 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1471 ), .Q(n5879) );
  NAND2X0 U5875 ( .IN1(n5881), .IN2(n5882), .QN(n5862) );
  MUX21X1 U5876 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1474 ), .Q(n5882) );
  MUX21X1 U5877 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1475 ), .Q(n5881) );
  NAND2X0 U5878 ( .IN1(n5883), .IN2(n5884), .QN(n5861) );
  MUX21X1 U5879 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1472 ), .Q(n5884) );
  MUX21X1 U5880 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1473 ), .Q(n5883) );
  XOR3X1 U5881 ( .IN1(n5850), .IN2(n5848), .IN3(n5847), .Q(n5836) );
  NAND2X0 U5882 ( .IN1(n5885), .IN2(n5886), .QN(n5847) );
  MUX21X1 U5883 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1478 ), .Q(n5886) );
  MUX21X1 U5884 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1479 ), .Q(n5885) );
  NAND2X0 U5885 ( .IN1(n5887), .IN2(n5888), .QN(n5848) );
  MUX21X1 U5886 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1481 ), .Q(n5888) );
  MUX21X1 U5887 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1480 ), .Q(n5887) );
  NAND2X0 U5888 ( .IN1(n5889), .IN2(n5890), .QN(n5850) );
  MUX21X1 U5889 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1476 ), .Q(n5890) );
  MUX21X1 U5890 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1477 ), .Q(n5889) );
  AO22X1 U5891 ( .IN1(n5891), .IN2(n5892), .IN3(n5893), .IN4(n5894), .Q(n5837)
         );
  OR2X1 U5892 ( .IN1(n5892), .IN2(n5891), .Q(n5893) );
  XOR2X1 U5893 ( .IN1(n5895), .IN2(n5865), .Q(n5828) );
  AOI21X1 U5894 ( .IN1(n5896), .IN2(n3614), .IN3(n5897), .QN(n5865) );
  MUX21X1 U5895 ( .IN1(n3616), .IN2(n5898), .S(\i_m4stg_frac/n1469 ), .Q(n5897) );
  INVX0 U5896 ( .INP(n3818), .ZN(n5898) );
  INVX0 U5897 ( .INP(n3817), .ZN(n3616) );
  NAND3X0 U5898 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(n938), .IN3(
        \i_m4stg_frac/n656 ), .QN(n5895) );
  XOR2X1 U5899 ( .IN1(n5832), .IN2(n5829), .Q(n5878) );
  AO22X1 U5900 ( .IN1(n5899), .IN2(n5900), .IN3(n5901), .IN4(n5902), .Q(n5829)
         );
  OR2X1 U5901 ( .IN1(n5900), .IN2(n5899), .Q(n5901) );
  AO22X1 U5902 ( .IN1(n3526), .IN2(n3527), .IN3(n5903), .IN4(n3525), .Q(
        \i_m4stg_frac/a1cout[13] ) );
  AO22X1 U5903 ( .IN1(n5904), .IN2(n5905), .IN3(n5906), .IN4(n5907), .Q(n3525)
         );
  OR2X1 U5904 ( .IN1(n5905), .IN2(n5904), .Q(n5907) );
  OR2X1 U5905 ( .IN1(n3527), .IN2(n3526), .Q(n5903) );
  INVX0 U5906 ( .INP(n5908), .ZN(n3527) );
  MUX21X1 U5907 ( .IN1(n5909), .IN2(n5910), .S(n5911), .Q(n5908) );
  INVX0 U5908 ( .INP(n5912), .ZN(n5911) );
  XOR2X1 U5909 ( .IN1(n5877), .IN2(n5875), .Q(n3526) );
  INVX0 U5910 ( .INP(n5913), .ZN(n5875) );
  XNOR3X1 U5911 ( .IN1(n5914), .IN2(n5870), .IN3(n5874), .Q(n5877) );
  AO21X1 U5912 ( .IN1(n5915), .IN2(n5916), .IN3(n5833), .Q(n5874) );
  NOR2X0 U5913 ( .IN1(n5916), .IN2(n5915), .QN(n5833) );
  XNOR3X1 U5914 ( .IN1(n5894), .IN2(n5892), .IN3(n5891), .Q(n5916) );
  NAND2X0 U5915 ( .IN1(n5917), .IN2(n5918), .QN(n5891) );
  MUX21X1 U5916 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1477 ), .Q(n5918) );
  MUX21X1 U5917 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1478 ), .Q(n5917) );
  NAND2X0 U5918 ( .IN1(n5919), .IN2(n5920), .QN(n5892) );
  MUX21X1 U5919 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1480 ), .Q(n5920) );
  MUX21X1 U5920 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1479 ), .Q(n5919) );
  NAND2X0 U5921 ( .IN1(n5921), .IN2(n5922), .QN(n5894) );
  MUX21X1 U5922 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1475 ), .Q(n5922) );
  MUX21X1 U5923 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1476 ), .Q(n5921) );
  AOI22X1 U5924 ( .IN1(n5923), .IN2(n5924), .IN3(n5925), .IN4(n5926), .QN(
        n5915) );
  OR2X1 U5925 ( .IN1(n5924), .IN2(n5923), .Q(n5925) );
  XOR3X1 U5926 ( .IN1(n5899), .IN2(n5900), .IN3(n5902), .Q(n5870) );
  NAND2X0 U5927 ( .IN1(n5927), .IN2(n5928), .QN(n5902) );
  MUX21X1 U5928 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1469 ), .Q(n5928) );
  MUX21X1 U5929 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1470 ), .Q(n5927) );
  NAND2X0 U5930 ( .IN1(n5929), .IN2(n5930), .QN(n5900) );
  MUX21X1 U5931 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1474 ), .Q(n5930) );
  MUX21X1 U5932 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1473 ), .Q(n5929) );
  NAND2X0 U5933 ( .IN1(n5931), .IN2(n5932), .QN(n5899) );
  MUX21X1 U5934 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1472 ), .Q(n5932) );
  MUX21X1 U5935 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1471 ), .Q(n5931) );
  XNOR2X1 U5936 ( .IN1(n5872), .IN2(n5871), .Q(n5914) );
  AO22X1 U5937 ( .IN1(n5933), .IN2(n5934), .IN3(n5935), .IN4(n5936), .Q(n5871)
         );
  OR2X1 U5938 ( .IN1(n5934), .IN2(n5933), .Q(n5935) );
  AND2X1 U5939 ( .IN1(n5937), .IN2(n5832), .Q(n5872) );
  NAND3X0 U5940 ( .IN1(n5938), .IN2(n5939), .IN3(n3312), .QN(n5832) );
  AO21X1 U5941 ( .IN1(n3312), .IN2(n5938), .IN3(n5939), .Q(n5937) );
  NAND2X0 U5942 ( .IN1(n5940), .IN2(n5941), .QN(n5939) );
  NAND3X0 U5943 ( .IN1(\i_m4stg_frac/n659 ), .IN2(n1133), .IN3(n5896), .QN(
        n5941) );
  XOR2X1 U5944 ( .IN1(n1039), .IN2(\i_m4stg_frac/n1468 ), .Q(n5896) );
  MUX21X1 U5945 ( .IN1(n3781), .IN2(n3782), .S(\i_m4stg_frac/n1467 ), .Q(n5940) );
  NOR2X0 U5946 ( .IN1(\i_m4stg_frac/n659 ), .IN2(\i_m4stg_frac/n658 ), .QN(
        n3614) );
  NOR2X0 U5947 ( .IN1(\i_m4stg_frac/n658 ), .IN2(\i_m4stg_frac/n657 ), .QN(
        n3312) );
  AO22X1 U5948 ( .IN1(n3529), .IN2(n3530), .IN3(n5942), .IN4(n3528), .Q(
        \i_m4stg_frac/a1cout[12] ) );
  AO22X1 U5949 ( .IN1(n5943), .IN2(n5944), .IN3(n5945), .IN4(n5946), .Q(n3528)
         );
  NAND2X0 U5950 ( .IN1(n5947), .IN2(n3844), .QN(n5946) );
  OR2X1 U5951 ( .IN1(n3530), .IN2(n3529), .Q(n5942) );
  INVX0 U5952 ( .INP(n5948), .ZN(n3530) );
  MUX21X1 U5953 ( .IN1(n5949), .IN2(n5950), .S(n5951), .Q(n5948) );
  INVX0 U5954 ( .INP(n5952), .ZN(n5951) );
  XOR2X1 U5955 ( .IN1(n5912), .IN2(n5910), .Q(n3529) );
  INVX0 U5956 ( .INP(n5953), .ZN(n5910) );
  XNOR3X1 U5957 ( .IN1(n5954), .IN2(n5904), .IN3(n5909), .Q(n5912) );
  AO21X1 U5958 ( .IN1(n5955), .IN2(n5956), .IN3(n5913), .Q(n5909) );
  NOR2X0 U5959 ( .IN1(n5956), .IN2(n5955), .QN(n5913) );
  XNOR3X1 U5960 ( .IN1(n5926), .IN2(n5924), .IN3(n5923), .Q(n5956) );
  NAND2X0 U5961 ( .IN1(n5957), .IN2(n5958), .QN(n5923) );
  MUX21X1 U5962 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1476 ), .Q(n5958) );
  MUX21X1 U5963 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1477 ), .Q(n5957) );
  NAND2X0 U5964 ( .IN1(n5959), .IN2(n5960), .QN(n5924) );
  MUX21X1 U5965 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1479 ), .Q(n5960) );
  MUX21X1 U5966 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1478 ), .Q(n5959) );
  NAND2X0 U5967 ( .IN1(n5961), .IN2(n5962), .QN(n5926) );
  MUX21X1 U5968 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1474 ), .Q(n5962) );
  MUX21X1 U5969 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1475 ), .Q(n5961) );
  AOI22X1 U5970 ( .IN1(n5963), .IN2(n5964), .IN3(n5965), .IN4(n5966), .QN(
        n5955) );
  OR2X1 U5971 ( .IN1(n5964), .IN2(n5963), .Q(n5965) );
  XOR3X1 U5972 ( .IN1(n5933), .IN2(n5934), .IN3(n5936), .Q(n5904) );
  NAND2X0 U5973 ( .IN1(n5967), .IN2(n5968), .QN(n5936) );
  MUX21X1 U5974 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1468 ), .Q(n5968) );
  MUX21X1 U5975 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1469 ), .Q(n5967) );
  NAND2X0 U5976 ( .IN1(n5969), .IN2(n5970), .QN(n5934) );
  MUX21X1 U5977 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1472 ), .Q(n5970) );
  MUX21X1 U5978 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1473 ), .Q(n5969) );
  NAND2X0 U5979 ( .IN1(n5971), .IN2(n5972), .QN(n5933) );
  MUX21X1 U5980 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1470 ), .Q(n5972) );
  MUX21X1 U5981 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1471 ), .Q(n5971) );
  XNOR2X1 U5982 ( .IN1(n5906), .IN2(n5905), .Q(n5954) );
  AO22X1 U5983 ( .IN1(n5973), .IN2(n5974), .IN3(n5975), .IN4(n5976), .Q(n5905)
         );
  OR2X1 U5984 ( .IN1(n5974), .IN2(n5973), .Q(n5975) );
  NOR2X0 U5985 ( .IN1(n5938), .IN2(\i_m4stg_frac/n658 ), .QN(n5906) );
  NAND2X0 U5986 ( .IN1(\i_m4stg_frac/n659 ), .IN2(\i_m4stg_frac/n1467 ), .QN(
        n5938) );
  NOR2X0 U5987 ( .IN1(n3531), .IN2(n3532), .QN(\i_m4stg_frac/a1cout[11] ) );
  OAI22X1 U5988 ( .IN1(n5977), .IN2(n5978), .IN3(n5979), .IN4(n5980), .QN(
        n3532) );
  AND2X1 U5989 ( .IN1(n5978), .IN2(n5977), .Q(n5980) );
  XOR2X1 U5990 ( .IN1(n5952), .IN2(n5949), .Q(n3531) );
  INVX0 U5991 ( .INP(n5981), .ZN(n5949) );
  XNOR3X1 U5992 ( .IN1(n5982), .IN2(n5945), .IN3(n5950), .Q(n5952) );
  AO21X1 U5993 ( .IN1(n5983), .IN2(n5984), .IN3(n5953), .Q(n5950) );
  NOR2X0 U5994 ( .IN1(n5984), .IN2(n5983), .QN(n5953) );
  XNOR3X1 U5995 ( .IN1(n5966), .IN2(n5964), .IN3(n5963), .Q(n5984) );
  NAND2X0 U5996 ( .IN1(n5985), .IN2(n5986), .QN(n5963) );
  MUX21X1 U5997 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1475 ), .Q(n5986) );
  MUX21X1 U5998 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1476 ), .Q(n5985) );
  NAND2X0 U5999 ( .IN1(n5987), .IN2(n5988), .QN(n5964) );
  MUX21X1 U6000 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1478 ), .Q(n5988) );
  MUX21X1 U6001 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1477 ), .Q(n5987) );
  NAND2X0 U6002 ( .IN1(n5989), .IN2(n5990), .QN(n5966) );
  MUX21X1 U6003 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1474 ), .Q(n5990) );
  MUX21X1 U6004 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1473 ), .Q(n5989) );
  AOI22X1 U6005 ( .IN1(n5991), .IN2(n5992), .IN3(n5993), .IN4(n5994), .QN(
        n5983) );
  OR2X1 U6006 ( .IN1(n5992), .IN2(n5991), .Q(n5993) );
  XOR3X1 U6007 ( .IN1(n5973), .IN2(n5974), .IN3(n5976), .Q(n5945) );
  NAND2X0 U6008 ( .IN1(n5995), .IN2(n5996), .QN(n5976) );
  MUX21X1 U6009 ( .IN1(n3844), .IN2(n3845), .S(\i_m4stg_frac/n1467 ), .Q(n5996) );
  MUX21X1 U6010 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1468 ), .Q(n5995) );
  NAND2X0 U6011 ( .IN1(n5997), .IN2(n5998), .QN(n5974) );
  MUX21X1 U6012 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1472 ), .Q(n5998) );
  MUX21X1 U6013 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1471 ), .Q(n5997) );
  NAND2X0 U6014 ( .IN1(n5999), .IN2(n6000), .QN(n5973) );
  MUX21X1 U6015 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1469 ), .Q(n6000) );
  MUX21X1 U6016 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1470 ), .Q(n5999) );
  XOR2X1 U6017 ( .IN1(n5944), .IN2(n5943), .Q(n5982) );
  INVX0 U6018 ( .INP(n5947), .ZN(n5943) );
  AO22X1 U6019 ( .IN1(n6001), .IN2(n6002), .IN3(n6003), .IN4(n6004), .Q(n5947)
         );
  OR2X1 U6020 ( .IN1(n6002), .IN2(n6001), .Q(n6004) );
  NOR2X0 U6021 ( .IN1(n3610), .IN2(\i_m4stg_frac/n662 ), .QN(n5944) );
  AO22X1 U6022 ( .IN1(n3535), .IN2(n3534), .IN3(n3533), .IN4(n6005), .Q(
        \i_m4stg_frac/a1cout[10] ) );
  OR2X1 U6023 ( .IN1(n3535), .IN2(n3534), .Q(n6005) );
  AOI21X1 U6024 ( .IN1(n6006), .IN2(n6007), .IN3(n5981), .QN(n3533) );
  NOR2X0 U6025 ( .IN1(n6007), .IN2(n6006), .QN(n5981) );
  XNOR3X1 U6026 ( .IN1(n5994), .IN2(n5992), .IN3(n5991), .Q(n6007) );
  NAND2X0 U6027 ( .IN1(n6008), .IN2(n6009), .QN(n5991) );
  MUX21X1 U6028 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1474 ), .Q(n6009) );
  MUX21X1 U6029 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1475 ), .Q(n6008) );
  NAND2X0 U6030 ( .IN1(n6010), .IN2(n6011), .QN(n5992) );
  MUX21X1 U6031 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1477 ), .Q(n6011) );
  MUX21X1 U6032 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1476 ), .Q(n6010) );
  NAND2X0 U6033 ( .IN1(n6012), .IN2(n6013), .QN(n5994) );
  MUX21X1 U6034 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1472 ), .Q(n6013) );
  MUX21X1 U6035 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1473 ), .Q(n6012) );
  AOI22X1 U6036 ( .IN1(n6014), .IN2(n6015), .IN3(n6016), .IN4(n6017), .QN(
        n6006) );
  OR2X1 U6037 ( .IN1(n6014), .IN2(n6015), .Q(n6016) );
  AO22X1 U6038 ( .IN1(n3541), .IN2(n3540), .IN3(n6018), .IN4(n3539), .Q(n3534)
         );
  AO22X1 U6039 ( .IN1(n3559), .IN2(n3558), .IN3(n6019), .IN4(n3557), .Q(n3539)
         );
  NAND2X0 U6040 ( .IN1(n6020), .IN2(n6021), .QN(n3557) );
  MUX21X1 U6041 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1472 ), .Q(n6021) );
  MUX21X1 U6042 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1473 ), .Q(n6020) );
  OR2X1 U6043 ( .IN1(n3558), .IN2(n3559), .Q(n6019) );
  NAND2X0 U6044 ( .IN1(n6022), .IN2(n6023), .QN(n3558) );
  MUX21X1 U6045 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1474 ), .Q(n6023) );
  MUX21X1 U6046 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1475 ), .Q(n6022) );
  NAND2X0 U6047 ( .IN1(n6024), .IN2(n6025), .QN(n3559) );
  MUX21X1 U6048 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1470 ), .Q(n6025) );
  MUX21X1 U6049 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1471 ), .Q(n6024) );
  OR2X1 U6050 ( .IN1(n3540), .IN2(n3541), .Q(n6018) );
  XNOR3X1 U6051 ( .IN1(n3890), .IN2(n6026), .IN3(n6027), .Q(n3540) );
  XOR3X1 U6052 ( .IN1(n6017), .IN2(n6015), .IN3(n6014), .Q(n3541) );
  NAND2X0 U6053 ( .IN1(n6028), .IN2(n6029), .QN(n6014) );
  MUX21X1 U6054 ( .IN1(n3593), .IN2(n3594), .S(\i_m4stg_frac/n1472 ), .Q(n6029) );
  NOR2X0 U6055 ( .IN1(n948), .IN2(n3665), .QN(n3942) );
  MUX21X1 U6056 ( .IN1(n3591), .IN2(n3592), .S(\i_m4stg_frac/n1471 ), .Q(n6028) );
  NOR2X0 U6057 ( .IN1(n3665), .IN2(\i_m4stg_frac/n671 ), .QN(n3687) );
  NAND2X0 U6058 ( .IN1(n1142), .IN2(n937), .QN(n3665) );
  NAND2X0 U6059 ( .IN1(n6030), .IN2(n6031), .QN(n6015) );
  MUX21X1 U6060 ( .IN1(n3585), .IN2(n3586), .S(\i_m4stg_frac/n1476 ), .Q(n6031) );
  NOR2X0 U6061 ( .IN1(\i_m4stg_frac/n676 ), .IN2(\i_m4stg_frac/n675 ), .QN(
        n3506) );
  MUX21X1 U6062 ( .IN1(n3587), .IN2(n3588), .S(\i_m4stg_frac/n1475 ), .Q(n6030) );
  NOR2X0 U6063 ( .IN1(\i_m4stg_frac/n677 ), .IN2(\i_m4stg_frac/n676 ), .QN(
        n3820) );
  NAND2X0 U6064 ( .IN1(n6032), .IN2(n6033), .QN(n6017) );
  MUX21X1 U6065 ( .IN1(n3579), .IN2(n3580), .S(\i_m4stg_frac/n1474 ), .Q(n6033) );
  MUX21X1 U6066 ( .IN1(n3581), .IN2(n3582), .S(\i_m4stg_frac/n1473 ), .Q(n6032) );
  NOR2X0 U6067 ( .IN1(\i_m4stg_frac/n672 ), .IN2(\i_m4stg_frac/n673 ), .QN(
        n3721) );
  XNOR3X1 U6068 ( .IN1(n3868), .IN2(n5977), .IN3(n5979), .Q(n3535) );
  XNOR3X1 U6069 ( .IN1(n6002), .IN2(n6001), .IN3(n6003), .Q(n5979) );
  AND2X1 U6070 ( .IN1(n6034), .IN2(n6035), .Q(n6003) );
  MUX21X1 U6071 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1468 ), .Q(n6035) );
  MUX21X1 U6072 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1469 ), .Q(n6034) );
  AND2X1 U6073 ( .IN1(n6036), .IN2(n6037), .Q(n6001) );
  MUX21X1 U6074 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1471 ), .Q(n6037) );
  MUX21X1 U6075 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1470 ), .Q(n6036) );
  MUX21X1 U6076 ( .IN1(n3868), .IN2(n3869), .S(\i_m4stg_frac/n1467 ), .Q(n6002) );
  AO22X1 U6077 ( .IN1(n6038), .IN2(n6039), .IN3(n6040), .IN4(n6041), .Q(n5977)
         );
  NAND2X0 U6078 ( .IN1(n6027), .IN2(n6026), .QN(n6041) );
  INVX0 U6079 ( .INP(n6039), .ZN(n6026) );
  INVX0 U6080 ( .INP(n6038), .ZN(n6027) );
  INVX0 U6081 ( .INP(n3890), .ZN(n6040) );
  NAND2X0 U6082 ( .IN1(n6042), .IN2(n6043), .QN(n6039) );
  MUX21X1 U6083 ( .IN1(n3890), .IN2(n3891), .S(\i_m4stg_frac/n1467 ), .Q(n6043) );
  MUX21X1 U6084 ( .IN1(n3647), .IN2(n3550), .S(\i_m4stg_frac/n1468 ), .Q(n6042) );
  NOR2X0 U6085 ( .IN1(\i_m4stg_frac/n663 ), .IN2(\i_m4stg_frac/n664 ), .QN(
        n3630) );
  NAND2X0 U6086 ( .IN1(n6044), .IN2(n6045), .QN(n6038) );
  MUX21X1 U6087 ( .IN1(n3569), .IN2(n3570), .S(\i_m4stg_frac/n1470 ), .Q(n6045) );
  AND2X1 U6088 ( .IN1(\i_m4stg_frac/n668 ), .IN2(n1168), .Q(n3606) );
  INVX0 U6089 ( .INP(n3651), .ZN(n3602) );
  NAND2X0 U6090 ( .IN1(n1168), .IN2(n912), .QN(n3651) );
  MUX21X1 U6091 ( .IN1(n3567), .IN2(n3568), .S(\i_m4stg_frac/n1469 ), .Q(n6044) );
  NOR2X0 U6092 ( .IN1(\i_m4stg_frac/n667 ), .IN2(\i_m4stg_frac/n668 ), .QN(
        n3670) );
  NOR2X0 U6093 ( .IN1(n949), .IN2(n3610), .QN(n5978) );
  NAND2X0 U6094 ( .IN1(n1143), .IN2(n934), .QN(n3610) );
  XOR3X1 U6095 ( .IN1(n6046), .IN2(n6047), .IN3(n6048), .Q(
        \i_m4stg_frac/a0sum[9] ) );
  XOR3X1 U6096 ( .IN1(n6049), .IN2(n6050), .IN3(n6051), .Q(
        \i_m4stg_frac/a0sum[8] ) );
  XOR2X1 U6097 ( .IN1(n6052), .IN2(n6053), .Q(\i_m4stg_frac/a0sum[7] ) );
  XOR2X1 U6098 ( .IN1(n6054), .IN2(n6055), .Q(\i_m4stg_frac/a0sum[79] ) );
  XNOR2X1 U6099 ( .IN1(n6055), .IN2(n6056), .Q(\i_m4stg_frac/a0sum[78] ) );
  NAND2X0 U6100 ( .IN1(n6057), .IN2(n6058), .QN(n6056) );
  XOR3X1 U6101 ( .IN1(n6059), .IN2(n6060), .IN3(n6061), .Q(
        \i_m4stg_frac/a0sum[77] ) );
  XNOR2X1 U6102 ( .IN1(n6062), .IN2(n6063), .Q(\i_m4stg_frac/a0sum[76] ) );
  NAND2X0 U6103 ( .IN1(n6064), .IN2(n6065), .QN(n6063) );
  XOR2X1 U6104 ( .IN1(n6066), .IN2(n6067), .Q(\i_m4stg_frac/a0sum[75] ) );
  AND2X1 U6105 ( .IN1(n6068), .IN2(n6069), .Q(n6066) );
  XOR3X1 U6106 ( .IN1(n6070), .IN2(n6071), .IN3(n6072), .Q(
        \i_m4stg_frac/a0sum[74] ) );
  XNOR2X1 U6107 ( .IN1(n6073), .IN2(n6074), .Q(\i_m4stg_frac/a0sum[73] ) );
  NOR2X0 U6108 ( .IN1(n6075), .IN2(n6076), .QN(n6074) );
  XNOR3X1 U6109 ( .IN1(n6077), .IN2(n6078), .IN3(n6079), .Q(
        \i_m4stg_frac/a0sum[72] ) );
  XOR3X1 U6110 ( .IN1(n6080), .IN2(n6081), .IN3(n6082), .Q(
        \i_m4stg_frac/a0sum[71] ) );
  XOR3X1 U6111 ( .IN1(n6083), .IN2(n6084), .IN3(n6085), .Q(
        \i_m4stg_frac/a0sum[70] ) );
  XOR2X1 U6112 ( .IN1(n6086), .IN2(n6087), .Q(\i_m4stg_frac/a0sum[6] ) );
  XOR3X1 U6113 ( .IN1(n6088), .IN2(n6089), .IN3(n6090), .Q(
        \i_m4stg_frac/a0sum[69] ) );
  XOR3X1 U6114 ( .IN1(n6091), .IN2(n6092), .IN3(n6093), .Q(
        \i_m4stg_frac/a0sum[68] ) );
  XOR3X1 U6115 ( .IN1(n6094), .IN2(n6095), .IN3(n6096), .Q(
        \i_m4stg_frac/a0sum[67] ) );
  XOR3X1 U6116 ( .IN1(n6097), .IN2(n6098), .IN3(n6099), .Q(
        \i_m4stg_frac/a0sum[66] ) );
  XOR3X1 U6117 ( .IN1(n6100), .IN2(n6101), .IN3(n6102), .Q(
        \i_m4stg_frac/a0sum[65] ) );
  XOR3X1 U6118 ( .IN1(n6103), .IN2(n6104), .IN3(n6105), .Q(
        \i_m4stg_frac/a0sum[64] ) );
  XOR3X1 U6119 ( .IN1(n6106), .IN2(n6107), .IN3(n6108), .Q(
        \i_m4stg_frac/a0sum[63] ) );
  XOR3X1 U6120 ( .IN1(n6109), .IN2(n6110), .IN3(n6111), .Q(
        \i_m4stg_frac/a0sum[62] ) );
  XOR3X1 U6121 ( .IN1(n6112), .IN2(n6113), .IN3(n6114), .Q(
        \i_m4stg_frac/a0sum[61] ) );
  XOR3X1 U6122 ( .IN1(n6115), .IN2(n6116), .IN3(n6117), .Q(
        \i_m4stg_frac/a0sum[60] ) );
  XOR2X1 U6123 ( .IN1(n6118), .IN2(n6119), .Q(\i_m4stg_frac/a0sum[5] ) );
  XOR3X1 U6124 ( .IN1(n6120), .IN2(n6121), .IN3(n6122), .Q(
        \i_m4stg_frac/a0sum[59] ) );
  XOR3X1 U6125 ( .IN1(n6123), .IN2(n6124), .IN3(n6125), .Q(
        \i_m4stg_frac/a0sum[58] ) );
  XOR3X1 U6126 ( .IN1(n6126), .IN2(n6127), .IN3(n6128), .Q(
        \i_m4stg_frac/a0sum[57] ) );
  XOR3X1 U6127 ( .IN1(n6129), .IN2(n6130), .IN3(n6131), .Q(
        \i_m4stg_frac/a0sum[56] ) );
  XOR3X1 U6128 ( .IN1(n6132), .IN2(n6133), .IN3(n6134), .Q(
        \i_m4stg_frac/a0sum[55] ) );
  XOR3X1 U6129 ( .IN1(n6135), .IN2(n6136), .IN3(n6137), .Q(
        \i_m4stg_frac/a0sum[54] ) );
  XOR3X1 U6130 ( .IN1(n6138), .IN2(n6139), .IN3(n6140), .Q(
        \i_m4stg_frac/a0sum[53] ) );
  XOR3X1 U6131 ( .IN1(n6141), .IN2(n6142), .IN3(n6143), .Q(
        \i_m4stg_frac/a0sum[52] ) );
  XOR3X1 U6132 ( .IN1(n6144), .IN2(n6145), .IN3(n6146), .Q(
        \i_m4stg_frac/a0sum[51] ) );
  XOR3X1 U6133 ( .IN1(n6147), .IN2(n6148), .IN3(n6149), .Q(
        \i_m4stg_frac/a0sum[50] ) );
  XOR2X1 U6134 ( .IN1(n6150), .IN2(n6151), .Q(\i_m4stg_frac/a0sum[4] ) );
  XOR3X1 U6135 ( .IN1(n6152), .IN2(n6153), .IN3(n6154), .Q(
        \i_m4stg_frac/a0sum[49] ) );
  XOR3X1 U6136 ( .IN1(n6155), .IN2(n6156), .IN3(n6157), .Q(
        \i_m4stg_frac/a0sum[48] ) );
  XOR3X1 U6137 ( .IN1(n6158), .IN2(n6159), .IN3(n6160), .Q(
        \i_m4stg_frac/a0sum[47] ) );
  XOR3X1 U6138 ( .IN1(n6161), .IN2(n6162), .IN3(n6163), .Q(
        \i_m4stg_frac/a0sum[46] ) );
  XOR3X1 U6139 ( .IN1(n6164), .IN2(n6165), .IN3(n6166), .Q(
        \i_m4stg_frac/a0sum[45] ) );
  XOR3X1 U6140 ( .IN1(n6167), .IN2(n6168), .IN3(n6169), .Q(
        \i_m4stg_frac/a0sum[44] ) );
  XOR3X1 U6141 ( .IN1(n6170), .IN2(n6171), .IN3(n6172), .Q(
        \i_m4stg_frac/a0sum[43] ) );
  XOR3X1 U6142 ( .IN1(n6173), .IN2(n6174), .IN3(n6175), .Q(
        \i_m4stg_frac/a0sum[42] ) );
  XOR3X1 U6143 ( .IN1(n6176), .IN2(n6177), .IN3(n6178), .Q(
        \i_m4stg_frac/a0sum[41] ) );
  XOR3X1 U6144 ( .IN1(n6179), .IN2(n6180), .IN3(n6181), .Q(
        \i_m4stg_frac/a0sum[40] ) );
  XOR3X1 U6145 ( .IN1(n6182), .IN2(n6183), .IN3(n6184), .Q(
        \i_m4stg_frac/a0sum[3] ) );
  XOR3X1 U6146 ( .IN1(n6185), .IN2(n6186), .IN3(n6187), .Q(
        \i_m4stg_frac/a0sum[39] ) );
  XOR3X1 U6147 ( .IN1(n6188), .IN2(n6189), .IN3(n6190), .Q(
        \i_m4stg_frac/a0sum[38] ) );
  XOR3X1 U6148 ( .IN1(n6191), .IN2(n6192), .IN3(n6193), .Q(
        \i_m4stg_frac/a0sum[37] ) );
  XOR3X1 U6149 ( .IN1(n6194), .IN2(n6195), .IN3(n6196), .Q(
        \i_m4stg_frac/a0sum[36] ) );
  XOR3X1 U6150 ( .IN1(n6197), .IN2(n6198), .IN3(n6199), .Q(
        \i_m4stg_frac/a0sum[35] ) );
  XOR3X1 U6151 ( .IN1(n6200), .IN2(n6201), .IN3(n6202), .Q(
        \i_m4stg_frac/a0sum[34] ) );
  XOR3X1 U6152 ( .IN1(n6203), .IN2(n6204), .IN3(n6205), .Q(
        \i_m4stg_frac/a0sum[33] ) );
  XOR3X1 U6153 ( .IN1(n6206), .IN2(n6207), .IN3(n6208), .Q(
        \i_m4stg_frac/a0sum[32] ) );
  XOR3X1 U6154 ( .IN1(n6209), .IN2(n6210), .IN3(n6211), .Q(
        \i_m4stg_frac/a0sum[31] ) );
  XOR3X1 U6155 ( .IN1(n6212), .IN2(n6213), .IN3(n6214), .Q(
        \i_m4stg_frac/a0sum[30] ) );
  OA21X1 U6156 ( .IN1(n6215), .IN2(n6216), .IN3(n6183), .Q(
        \i_m4stg_frac/a0sum[2] ) );
  XOR3X1 U6157 ( .IN1(n6217), .IN2(n6218), .IN3(n6219), .Q(
        \i_m4stg_frac/a0sum[29] ) );
  XOR3X1 U6158 ( .IN1(n6220), .IN2(n6221), .IN3(n6222), .Q(
        \i_m4stg_frac/a0sum[28] ) );
  XOR3X1 U6159 ( .IN1(n6223), .IN2(n6224), .IN3(n6225), .Q(
        \i_m4stg_frac/a0sum[27] ) );
  XOR3X1 U6160 ( .IN1(n6226), .IN2(n6227), .IN3(n6228), .Q(
        \i_m4stg_frac/a0sum[26] ) );
  XOR3X1 U6161 ( .IN1(n6229), .IN2(n6230), .IN3(n6231), .Q(
        \i_m4stg_frac/a0sum[25] ) );
  XOR3X1 U6162 ( .IN1(n6232), .IN2(n6233), .IN3(n6234), .Q(
        \i_m4stg_frac/a0sum[24] ) );
  XOR3X1 U6163 ( .IN1(n6235), .IN2(n6236), .IN3(n6237), .Q(
        \i_m4stg_frac/a0sum[23] ) );
  XOR3X1 U6164 ( .IN1(n6238), .IN2(n6239), .IN3(n6240), .Q(
        \i_m4stg_frac/a0sum[22] ) );
  XOR3X1 U6165 ( .IN1(n6241), .IN2(n6242), .IN3(n6243), .Q(
        \i_m4stg_frac/a0sum[21] ) );
  XOR3X1 U6166 ( .IN1(n6244), .IN2(n6245), .IN3(n6246), .Q(
        \i_m4stg_frac/a0sum[20] ) );
  NOR2X0 U6167 ( .IN1(n6215), .IN2(n6247), .QN(\i_m4stg_frac/a0sum[1] ) );
  AOI21X1 U6168 ( .IN1(n1034), .IN2(n6248), .IN3(n6249), .QN(n6247) );
  XOR3X1 U6169 ( .IN1(n6250), .IN2(n6251), .IN3(n6252), .Q(
        \i_m4stg_frac/a0sum[19] ) );
  XOR3X1 U6170 ( .IN1(n6253), .IN2(n6254), .IN3(n6255), .Q(
        \i_m4stg_frac/a0sum[18] ) );
  XOR3X1 U6171 ( .IN1(n6256), .IN2(n6257), .IN3(n6258), .Q(
        \i_m4stg_frac/a0sum[17] ) );
  XOR3X1 U6172 ( .IN1(n6259), .IN2(n6260), .IN3(n6261), .Q(
        \i_m4stg_frac/a0sum[16] ) );
  XOR3X1 U6173 ( .IN1(n6262), .IN2(n6263), .IN3(n6264), .Q(
        \i_m4stg_frac/a0sum[15] ) );
  XOR3X1 U6174 ( .IN1(n6265), .IN2(n6266), .IN3(n6267), .Q(
        \i_m4stg_frac/a0sum[14] ) );
  XOR3X1 U6175 ( .IN1(n6268), .IN2(n6269), .IN3(n6270), .Q(
        \i_m4stg_frac/a0sum[13] ) );
  XOR3X1 U6176 ( .IN1(n6271), .IN2(n6272), .IN3(n6273), .Q(
        \i_m4stg_frac/a0sum[12] ) );
  XOR2X1 U6177 ( .IN1(n6274), .IN2(n6275), .Q(\i_m4stg_frac/a0sum[11] ) );
  XOR3X1 U6178 ( .IN1(n6276), .IN2(n6277), .IN3(n6278), .Q(
        \i_m4stg_frac/a0sum[10] ) );
  NOR2X0 U6179 ( .IN1(n1034), .IN2(n6279), .QN(\i_m4stg_frac/a0sum[0] ) );
  AO22X1 U6180 ( .IN1(n6280), .IN2(n6281), .IN3(n6048), .IN4(n6282), .Q(
        \i_m4stg_frac/a0cout[9] ) );
  NAND2X0 U6181 ( .IN1(n6047), .IN2(n6046), .QN(n6282) );
  INVX0 U6182 ( .INP(n6280), .ZN(n6047) );
  XNOR3X1 U6183 ( .IN1(n6283), .IN2(n6284), .IN3(n6285), .Q(n6048) );
  INVX0 U6184 ( .INP(n6046), .ZN(n6281) );
  OA22X1 U6185 ( .IN1(n6286), .IN2(n6287), .IN3(n6288), .IN4(n6289), .Q(n6046)
         );
  AND2X1 U6186 ( .IN1(n6287), .IN2(n6286), .Q(n6289) );
  NAND2X0 U6187 ( .IN1(n6290), .IN2(n6291), .QN(n6280) );
  NAND3X0 U6188 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(n6292), .IN3(n6293), .QN(
        n6291) );
  INVX0 U6189 ( .INP(n6294), .ZN(n6293) );
  OAI21X1 U6190 ( .IN1(n6292), .IN2(n1034), .IN3(n6295), .QN(n6290) );
  AO22X1 U6191 ( .IN1(n6051), .IN2(n6049), .IN3(n6050), .IN4(n6296), .Q(
        \i_m4stg_frac/a0cout[8] ) );
  OR2X1 U6192 ( .IN1(n6049), .IN2(n6051), .Q(n6296) );
  INVX0 U6193 ( .INP(n6297), .ZN(n6050) );
  AO22X1 U6194 ( .IN1(n6298), .IN2(n6299), .IN3(n6300), .IN4(n6301), .Q(n6049)
         );
  OR2X1 U6195 ( .IN1(n6299), .IN2(n6298), .Q(n6301) );
  XNOR3X1 U6196 ( .IN1(n6288), .IN2(n6287), .IN3(n6286), .Q(n6051) );
  XNOR3X1 U6197 ( .IN1(n6302), .IN2(n6303), .IN3(n6304), .Q(n6286) );
  AOI22X1 U6198 ( .IN1(n6305), .IN2(n6306), .IN3(n6307), .IN4(n6308), .QN(
        n6287) );
  OR2X1 U6199 ( .IN1(n6306), .IN2(n6305), .Q(n6307) );
  XOR2X1 U6200 ( .IN1(n6309), .IN2(n6292), .Q(n6288) );
  NAND2X0 U6201 ( .IN1(n6310), .IN2(n6311), .QN(n6292) );
  MUX21X1 U6202 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1468 ), .Q(n6311) );
  MUX21X1 U6203 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1469 ), .Q(n6310) );
  NAND3X0 U6204 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(n1118), .IN3(
        \i_m4stg_frac/n1009 ), .QN(n6309) );
  NOR2X0 U6205 ( .IN1(n6053), .IN2(n6052), .QN(\i_m4stg_frac/a0cout[7] ) );
  AO22X1 U6206 ( .IN1(n6316), .IN2(n6317), .IN3(n6318), .IN4(n6319), .Q(n6052)
         );
  NAND2X0 U6207 ( .IN1(n6320), .IN2(n6321), .QN(n6318) );
  INVX0 U6208 ( .INP(n6320), .ZN(n6317) );
  INVX0 U6209 ( .INP(n6321), .ZN(n6316) );
  XNOR3X1 U6210 ( .IN1(n6300), .IN2(n6299), .IN3(n6298), .Q(n6053) );
  XOR3X1 U6211 ( .IN1(n6305), .IN2(n6306), .IN3(n6308), .Q(n6298) );
  NAND2X0 U6212 ( .IN1(n6322), .IN2(n6323), .QN(n6308) );
  MUX21X1 U6213 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1469 ), .Q(n6323) );
  MUX21X1 U6214 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1470 ), .Q(n6322) );
  NAND2X0 U6215 ( .IN1(n6328), .IN2(n6329), .QN(n6306) );
  MUX21X1 U6216 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1474 ), .Q(n6329) );
  MUX21X1 U6217 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1473 ), .Q(n6328) );
  NAND2X0 U6218 ( .IN1(n6334), .IN2(n6335), .QN(n6305) );
  MUX21X1 U6219 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1472 ), .Q(n6335) );
  MUX21X1 U6220 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1471 ), .Q(n6334) );
  AO22X1 U6221 ( .IN1(n6340), .IN2(n6341), .IN3(n6342), .IN4(n6343), .Q(n6299)
         );
  OR2X1 U6222 ( .IN1(n6341), .IN2(n6340), .Q(n6342) );
  AND2X1 U6223 ( .IN1(n6344), .IN2(n6297), .Q(n6300) );
  NAND3X0 U6224 ( .IN1(n6345), .IN2(n6346), .IN3(n6347), .QN(n6297) );
  AO21X1 U6225 ( .IN1(n6347), .IN2(n6345), .IN3(n6346), .Q(n6344) );
  NAND2X0 U6226 ( .IN1(n6348), .IN2(n6349), .QN(n6346) );
  MUX21X1 U6227 ( .IN1(n6350), .IN2(n6315), .S(\i_m4stg_frac/n1468 ), .Q(n6349) );
  NAND2X0 U6228 ( .IN1(n6351), .IN2(n913), .QN(n6350) );
  MUX21X1 U6229 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1467 ), .Q(n6348) );
  NAND2X0 U6230 ( .IN1(\i_m4stg_frac/n1012 ), .IN2(\i_m4stg_frac/n1467 ), .QN(
        n6345) );
  NOR2X0 U6231 ( .IN1(n6054), .IN2(n6055), .QN(\i_m4stg_frac/a0cout[79] ) );
  AND3X1 U6232 ( .IN1(n6055), .IN2(n6058), .IN3(n6057), .Q(
        \i_m4stg_frac/a0cout[78] ) );
  OA21X1 U6233 ( .IN1(n6352), .IN2(\i_m4stg_frac/n1000 ), .IN3(n6353), .Q(
        n6055) );
  OAI21X1 U6234 ( .IN1(n6061), .IN2(n6354), .IN3(n6060), .QN(
        \i_m4stg_frac/a0cout[77] ) );
  INVX0 U6235 ( .INP(n6059), .ZN(n6354) );
  XOR2X1 U6236 ( .IN1(n6058), .IN2(n6352), .Q(n6061) );
  INVX0 U6237 ( .INP(n6355), .ZN(n6058) );
  OAI22X1 U6238 ( .IN1(n6064), .IN2(n6062), .IN3(n6062), .IN4(n6065), .QN(
        \i_m4stg_frac/a0cout[76] ) );
  NAND2X0 U6239 ( .IN1(n6067), .IN2(n6356), .QN(n6065) );
  OA21X1 U6240 ( .IN1(n6357), .IN2(n6358), .IN3(n6059), .Q(n6062) );
  NAND2X0 U6241 ( .IN1(n6358), .IN2(n6357), .QN(n6059) );
  NAND2X0 U6242 ( .IN1(n6359), .IN2(n6060), .QN(n6358) );
  AO21X1 U6243 ( .IN1(n6360), .IN2(n6361), .IN3(n6352), .Q(n6060) );
  NAND3X0 U6244 ( .IN1(n6352), .IN2(n6361), .IN3(n6360), .QN(n6359) );
  NAND2X0 U6245 ( .IN1(n6362), .IN2(n6363), .QN(n6360) );
  NAND2X0 U6246 ( .IN1(n6364), .IN2(n6365), .QN(n6064) );
  OAI22X1 U6247 ( .IN1(n6067), .IN2(n6069), .IN3(n6067), .IN4(n6068), .QN(
        \i_m4stg_frac/a0cout[75] ) );
  INVX0 U6248 ( .INP(n6366), .ZN(n6068) );
  NAND2X0 U6249 ( .IN1(n6365), .IN2(n6367), .QN(n6069) );
  XOR3X1 U6250 ( .IN1(n6368), .IN2(n6356), .IN3(n6369), .Q(n6067) );
  XOR2X1 U6251 ( .IN1(n6364), .IN2(n6370), .Q(n6369) );
  OA21X1 U6252 ( .IN1(n6072), .IN2(n6071), .IN3(n6070), .Q(
        \i_m4stg_frac/a0cout[74] ) );
  AOI21X1 U6253 ( .IN1(n6371), .IN2(n6364), .IN3(n6366), .QN(n6070) );
  NOR2X0 U6254 ( .IN1(n6371), .IN2(n6364), .QN(n6366) );
  AND2X1 U6255 ( .IN1(n6372), .IN2(n6373), .Q(n6364) );
  MUX21X1 U6256 ( .IN1(n6374), .IN2(n936), .S(\i_m4stg_frac/n1006 ), .Q(n6372)
         );
  NAND2X0 U6257 ( .IN1(\i_m4stg_frac/n1530 ), .IN2(n936), .QN(n6374) );
  MUX21X1 U6258 ( .IN1(n6375), .IN2(n6365), .S(n6367), .Q(n6371) );
  NOR2X0 U6259 ( .IN1(n6376), .IN2(n6377), .QN(n6367) );
  NOR2X0 U6260 ( .IN1(n6368), .IN2(n6378), .QN(n6375) );
  AND2X1 U6261 ( .IN1(n6379), .IN2(n6365), .Q(n6071) );
  NOR2X0 U6262 ( .IN1(n6073), .IN2(n6380), .QN(n6072) );
  AO22X1 U6263 ( .IN1(n6073), .IN2(n6076), .IN3(n6075), .IN4(n6381), .Q(
        \i_m4stg_frac/a0cout[73] ) );
  OR2X1 U6264 ( .IN1(n6073), .IN2(n6076), .Q(n6381) );
  AND2X1 U6265 ( .IN1(n6077), .IN2(n6382), .Q(n6075) );
  AND2X1 U6266 ( .IN1(n6383), .IN2(n6365), .Q(n6076) );
  XOR3X1 U6267 ( .IN1(n6384), .IN2(n6368), .IN3(n6385), .Q(n6073) );
  XOR2X1 U6268 ( .IN1(n6378), .IN2(n6380), .Q(n6384) );
  XOR2X1 U6269 ( .IN1(n6377), .IN2(n6386), .Q(n6380) );
  OAI22X1 U6270 ( .IN1(n6077), .IN2(n6078), .IN3(n6079), .IN4(n6387), .QN(
        \i_m4stg_frac/a0cout[72] ) );
  AND2X1 U6271 ( .IN1(n6077), .IN2(n6078), .Q(n6387) );
  MUX21X1 U6272 ( .IN1(n6388), .IN2(n6389), .S(n6390), .Q(n6079) );
  INVX0 U6273 ( .INP(n6391), .ZN(n6390) );
  NAND2X0 U6274 ( .IN1(n6392), .IN2(n6365), .QN(n6078) );
  XOR3X1 U6275 ( .IN1(n6393), .IN2(n6368), .IN3(n6382), .Q(n6077) );
  AO221X1 U6276 ( .IN1(n6394), .IN2(n915), .IN3(n6386), .IN4(n6295), .IN5(
        n6385), .Q(n6382) );
  INVX0 U6277 ( .INP(n6379), .ZN(n6385) );
  NAND3X0 U6278 ( .IN1(n6376), .IN2(n6395), .IN3(n6396), .QN(n6379) );
  NAND2X0 U6279 ( .IN1(n6397), .IN2(n915), .QN(n6396) );
  INVX0 U6280 ( .INP(n6395), .ZN(n6295) );
  XOR2X1 U6281 ( .IN1(n6383), .IN2(n6370), .Q(n6393) );
  AO21X1 U6282 ( .IN1(n6398), .IN2(n6399), .IN3(n6394), .Q(n6383) );
  AO22X1 U6283 ( .IN1(n6080), .IN2(n6081), .IN3(n6082), .IN4(n6400), .Q(
        \i_m4stg_frac/a0cout[71] ) );
  NAND2X0 U6284 ( .IN1(n6401), .IN2(n6084), .QN(n6400) );
  XOR2X1 U6285 ( .IN1(n6391), .IN2(n6389), .Q(n6082) );
  INVX0 U6286 ( .INP(n6402), .ZN(n6389) );
  XOR3X1 U6287 ( .IN1(n6403), .IN2(n6368), .IN3(n6392), .Q(n6391) );
  AO21X1 U6288 ( .IN1(n6404), .IN2(n6398), .IN3(n6394), .Q(n6392) );
  XOR2X1 U6289 ( .IN1(n6378), .IN2(n6388), .Q(n6403) );
  XOR2X1 U6290 ( .IN1(n6347), .IN2(n6405), .Q(n6388) );
  INVX0 U6291 ( .INP(n6401), .ZN(n6080) );
  MUX21X1 U6292 ( .IN1(n6406), .IN2(n6402), .S(n6407), .Q(n6401) );
  AO22X1 U6293 ( .IN1(n6408), .IN2(n6081), .IN3(n6083), .IN4(n6409), .Q(
        \i_m4stg_frac/a0cout[70] ) );
  NAND2X0 U6294 ( .IN1(n6085), .IN2(n6084), .QN(n6409) );
  XOR2X1 U6295 ( .IN1(n6407), .IN2(n6406), .Q(n6083) );
  AOI22X1 U6296 ( .IN1(n6410), .IN2(n6411), .IN3(n6412), .IN4(n6413), .QN(
        n6406) );
  NAND2X0 U6297 ( .IN1(n6414), .IN2(n6415), .QN(n6412) );
  XNOR3X1 U6298 ( .IN1(n6416), .IN2(n6378), .IN3(n6402), .Q(n6407) );
  XOR2X1 U6299 ( .IN1(n6405), .IN2(n6404), .Q(n6402) );
  AO21X1 U6300 ( .IN1(n6417), .IN2(n6418), .IN3(n6419), .Q(n6404) );
  INVX0 U6301 ( .INP(n6314), .ZN(n6419) );
  INVX0 U6302 ( .INP(n6084), .ZN(n6081) );
  NAND2X0 U6303 ( .IN1(n6420), .IN2(n6365), .QN(n6084) );
  NAND2X0 U6304 ( .IN1(n6370), .IN2(n6357), .QN(n6365) );
  INVX0 U6305 ( .INP(n6378), .ZN(n6370) );
  INVX0 U6306 ( .INP(n6085), .ZN(n6408) );
  MUX21X1 U6307 ( .IN1(n6421), .IN2(n6422), .S(n6423), .Q(n6085) );
  NOR2X0 U6308 ( .IN1(n6087), .IN2(n6086), .QN(\i_m4stg_frac/a0cout[6] ) );
  XOR3X1 U6309 ( .IN1(n6319), .IN2(n6321), .IN3(n6320), .Q(n6086) );
  XOR3X1 U6310 ( .IN1(n6343), .IN2(n6341), .IN3(n6340), .Q(n6320) );
  NAND2X0 U6311 ( .IN1(n6424), .IN2(n6425), .QN(n6340) );
  MUX21X1 U6312 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1472 ), .Q(n6425) );
  MUX21X1 U6313 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1473 ), .Q(n6424) );
  NAND2X0 U6314 ( .IN1(n6426), .IN2(n6427), .QN(n6341) );
  MUX21X1 U6315 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1468 ), .Q(n6427) );
  MUX21X1 U6316 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1469 ), .Q(n6426) );
  NAND2X0 U6317 ( .IN1(n6428), .IN2(n6429), .QN(n6343) );
  MUX21X1 U6318 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1471 ), .Q(n6429) );
  MUX21X1 U6319 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1470 ), .Q(n6428) );
  AO22X1 U6320 ( .IN1(n6430), .IN2(n6431), .IN3(n6432), .IN4(n6433), .Q(n6321)
         );
  OR2X1 U6321 ( .IN1(n6431), .IN2(n6430), .Q(n6432) );
  NAND2X0 U6322 ( .IN1(n6351), .IN2(\i_m4stg_frac/n1467 ), .QN(n6319) );
  AOI22X1 U6323 ( .IN1(n6434), .IN2(n6435), .IN3(n6436), .IN4(n6437), .QN(
        n6087) );
  OR2X1 U6324 ( .IN1(n6435), .IN2(n6434), .Q(n6437) );
  AO22X1 U6325 ( .IN1(n6089), .IN2(n6090), .IN3(n6438), .IN4(n6088), .Q(
        \i_m4stg_frac/a0cout[69] ) );
  AO22X1 U6326 ( .IN1(n6439), .IN2(n6378), .IN3(n6440), .IN4(n6420), .Q(n6088)
         );
  OR2X1 U6327 ( .IN1(n6378), .IN2(n6439), .Q(n6440) );
  OR2X1 U6328 ( .IN1(n6090), .IN2(n6089), .Q(n6438) );
  INVX0 U6329 ( .INP(n6441), .ZN(n6090) );
  MUX21X1 U6330 ( .IN1(n6442), .IN2(n6443), .S(n6444), .Q(n6441) );
  XNOR2X1 U6331 ( .IN1(n6423), .IN2(n6422), .Q(n6089) );
  AOI22X1 U6332 ( .IN1(n6445), .IN2(n6415), .IN3(n6411), .IN4(n6446), .QN(
        n6422) );
  OR2X1 U6333 ( .IN1(n6445), .IN2(n6415), .Q(n6446) );
  XOR3X1 U6334 ( .IN1(n6416), .IN2(n6378), .IN3(n6421), .Q(n6423) );
  XOR2X1 U6335 ( .IN1(n6447), .IN2(n6413), .Q(n6421) );
  XOR2X1 U6336 ( .IN1(n6368), .IN2(n6448), .Q(n6416) );
  INVX0 U6337 ( .INP(n6357), .ZN(n6368) );
  NAND2X0 U6338 ( .IN1(n6449), .IN2(n6057), .QN(n6357) );
  INVX0 U6339 ( .INP(n6352), .ZN(n6057) );
  AO22X1 U6340 ( .IN1(n6092), .IN2(n6093), .IN3(n6450), .IN4(n6091), .Q(
        \i_m4stg_frac/a0cout[68] ) );
  AO22X1 U6341 ( .IN1(n6451), .IN2(n6420), .IN3(n6452), .IN4(n6449), .Q(n6091)
         );
  OA21X1 U6342 ( .IN1(n6451), .IN2(n6420), .IN3(n6453), .Q(n6452) );
  OR2X1 U6343 ( .IN1(n6093), .IN2(n6092), .Q(n6450) );
  INVX0 U6344 ( .INP(n6454), .ZN(n6093) );
  MUX21X1 U6345 ( .IN1(n6455), .IN2(n6456), .S(n6457), .Q(n6454) );
  INVX0 U6346 ( .INP(n6458), .ZN(n6457) );
  XOR2X1 U6347 ( .IN1(n6444), .IN2(n6442), .Q(n6092) );
  OA22X1 U6348 ( .IN1(n6459), .IN2(n6460), .IN3(n6414), .IN4(n6461), .Q(n6442)
         );
  AND2X1 U6349 ( .IN1(n6460), .IN2(n6459), .Q(n6461) );
  XOR3X1 U6350 ( .IN1(n6378), .IN2(n6443), .IN3(n6462), .Q(n6444) );
  XOR2X1 U6351 ( .IN1(n6420), .IN2(n6439), .Q(n6462) );
  XNOR2X1 U6352 ( .IN1(n6447), .IN2(n6445), .Q(n6443) );
  AO22X1 U6353 ( .IN1(n6463), .IN2(n6464), .IN3(n6465), .IN4(n6466), .Q(n6445)
         );
  OR2X1 U6354 ( .IN1(n6463), .IN2(n6464), .Q(n6465) );
  XOR2X1 U6355 ( .IN1(n6414), .IN2(n6410), .Q(n6447) );
  INVX0 U6356 ( .INP(n6415), .ZN(n6410) );
  NAND2X0 U6357 ( .IN1(n6467), .IN2(n6468), .QN(n6415) );
  MUX21X1 U6358 ( .IN1(n6469), .IN2(n935), .S(\i_m4stg_frac/n1015 ), .Q(n6467)
         );
  NAND2X0 U6359 ( .IN1(\i_m4stg_frac/n1530 ), .IN2(n935), .QN(n6469) );
  XNOR2X1 U6360 ( .IN1(n6352), .IN2(n6449), .Q(n6378) );
  NAND2X0 U6361 ( .IN1(n6470), .IN2(n976), .QN(n6352) );
  XOR2X1 U6362 ( .IN1(\i_m4stg_frac/n998 ), .IN2(n907), .Q(n6470) );
  AO22X1 U6363 ( .IN1(n6471), .IN2(n6472), .IN3(n6473), .IN4(n6095), .Q(
        \i_m4stg_frac/a0cout[67] ) );
  AO22X1 U6364 ( .IN1(n6474), .IN2(n6420), .IN3(n6475), .IN4(n6476), .Q(n6095)
         );
  NAND2X0 U6365 ( .IN1(n6448), .IN2(n6477), .QN(n6476) );
  NAND2X0 U6366 ( .IN1(n6094), .IN2(n6096), .QN(n6473) );
  INVX0 U6367 ( .INP(n6094), .ZN(n6472) );
  MUX21X1 U6368 ( .IN1(n6478), .IN2(n6479), .S(n6480), .Q(n6094) );
  INVX0 U6369 ( .INP(n6481), .ZN(n6480) );
  INVX0 U6370 ( .INP(n6096), .ZN(n6471) );
  XOR2X1 U6371 ( .IN1(n6458), .IN2(n6455), .Q(n6096) );
  OA22X1 U6372 ( .IN1(n6482), .IN2(n6483), .IN3(n6414), .IN4(n6484), .Q(n6455)
         );
  AND2X1 U6373 ( .IN1(n6483), .IN2(n6482), .Q(n6484) );
  XOR3X1 U6374 ( .IN1(n6485), .IN2(n6456), .IN3(n6486), .Q(n6458) );
  XOR2X1 U6375 ( .IN1(n6451), .IN2(n6420), .Q(n6486) );
  AOI21X1 U6376 ( .IN1(n6487), .IN2(n6488), .IN3(n6439), .QN(n6451) );
  NOR2X0 U6377 ( .IN1(n6488), .IN2(n6487), .QN(n6439) );
  AND2X1 U6378 ( .IN1(n6489), .IN2(n6490), .Q(n6487) );
  MUX21X1 U6379 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1519 ), .Q(n6490) );
  MUX21X1 U6380 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1530 ), .Q(n6489) );
  XOR3X1 U6381 ( .IN1(n6459), .IN2(n6414), .IN3(n6460), .Q(n6456) );
  OA22X1 U6382 ( .IN1(n6464), .IN2(n6494), .IN3(n6495), .IN4(n6496), .Q(n6460)
         );
  AND2X1 U6383 ( .IN1(n6494), .IN2(n6464), .Q(n6496) );
  XOR2X1 U6384 ( .IN1(n6497), .IN2(n6466), .Q(n6459) );
  NAND2X0 U6385 ( .IN1(n6449), .IN2(n6453), .QN(n6485) );
  INVX0 U6386 ( .INP(n6488), .ZN(n6449) );
  AO22X1 U6387 ( .IN1(n6098), .IN2(n6099), .IN3(n6498), .IN4(n6097), .Q(
        \i_m4stg_frac/a0cout[66] ) );
  AO22X1 U6388 ( .IN1(n6499), .IN2(n6420), .IN3(n6500), .IN4(n6501), .Q(n6097)
         );
  NAND2X0 U6389 ( .IN1(n6448), .IN2(n6502), .QN(n6501) );
  AND2X1 U6390 ( .IN1(n6503), .IN2(n6504), .Q(n6500) );
  INVX0 U6391 ( .INP(n6502), .ZN(n6499) );
  OR2X1 U6392 ( .IN1(n6099), .IN2(n6098), .Q(n6498) );
  INVX0 U6393 ( .INP(n6505), .ZN(n6099) );
  MUX21X1 U6394 ( .IN1(n6506), .IN2(n6507), .S(n6508), .Q(n6505) );
  INVX0 U6395 ( .INP(n6509), .ZN(n6508) );
  XNOR2X1 U6396 ( .IN1(n6481), .IN2(n6478), .Q(n6098) );
  AOI22X1 U6397 ( .IN1(n6510), .IN2(n6511), .IN3(n6411), .IN4(n6512), .QN(
        n6478) );
  OR2X1 U6398 ( .IN1(n6511), .IN2(n6510), .Q(n6512) );
  XOR3X1 U6399 ( .IN1(n6448), .IN2(n6475), .IN3(n6513), .Q(n6481) );
  XOR2X1 U6400 ( .IN1(n6474), .IN2(n6479), .Q(n6513) );
  XOR3X1 U6401 ( .IN1(n6483), .IN2(n6414), .IN3(n6482), .Q(n6479) );
  XOR2X1 U6402 ( .IN1(n6497), .IN2(n6494), .Q(n6482) );
  OA21X1 U6403 ( .IN1(n6514), .IN2(\i_m4stg_frac/n1018 ), .IN3(n6336), .Q(
        n6494) );
  XOR2X1 U6404 ( .IN1(n6464), .IN2(n6495), .Q(n6497) );
  AOI21X1 U6405 ( .IN1(n6515), .IN2(n6516), .IN3(n6517), .QN(n6483) );
  INVX0 U6406 ( .INP(n6477), .ZN(n6474) );
  XOR2X1 U6407 ( .IN1(n6488), .IN2(n6453), .Q(n6477) );
  NAND2X0 U6408 ( .IN1(n6518), .IN2(n6519), .QN(n6453) );
  MUX21X1 U6409 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1519 ), .Q(n6519) );
  MUX21X1 U6410 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1518 ), .Q(n6518) );
  NAND2X0 U6411 ( .IN1(n6363), .IN2(n1229), .QN(n6488) );
  AO22X1 U6412 ( .IN1(n6102), .IN2(n6101), .IN3(n6520), .IN4(n6100), .Q(
        \i_m4stg_frac/a0cout[65] ) );
  AO22X1 U6413 ( .IN1(n6521), .IN2(n6522), .IN3(n6523), .IN4(n6524), .Q(n6100)
         );
  OR2X1 U6414 ( .IN1(n6521), .IN2(n6522), .Q(n6524) );
  OR2X1 U6415 ( .IN1(n6101), .IN2(n6102), .Q(n6520) );
  INVX0 U6416 ( .INP(n6525), .ZN(n6101) );
  MUX21X1 U6417 ( .IN1(n6526), .IN2(n6527), .S(n6528), .Q(n6525) );
  INVX0 U6418 ( .INP(n6529), .ZN(n6528) );
  XOR2X1 U6419 ( .IN1(n6509), .IN2(n6507), .Q(n6102) );
  AOI22X1 U6420 ( .IN1(n6530), .IN2(n6411), .IN3(n6531), .IN4(n6532), .QN(
        n6507) );
  OR2X1 U6421 ( .IN1(n6411), .IN2(n6530), .Q(n6531) );
  XNOR3X1 U6422 ( .IN1(n6533), .IN2(n6506), .IN3(n6534), .Q(n6509) );
  XOR2X1 U6423 ( .IN1(n6502), .IN2(n6448), .Q(n6534) );
  INVX0 U6424 ( .INP(n6420), .ZN(n6448) );
  AO21X1 U6425 ( .IN1(n6535), .IN2(n6398), .IN3(n6394), .Q(n6420) );
  INVX0 U6426 ( .INP(n6536), .ZN(n6398) );
  AO21X1 U6427 ( .IN1(n6537), .IN2(n6538), .IN3(n6475), .Q(n6502) );
  NOR2X0 U6428 ( .IN1(n6537), .IN2(n6538), .QN(n6475) );
  AND2X1 U6429 ( .IN1(n6539), .IN2(n6540), .Q(n6538) );
  MUX21X1 U6430 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1517 ), .Q(n6540) );
  MUX21X1 U6431 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1518 ), .Q(n6539) );
  AOI21X1 U6432 ( .IN1(n6541), .IN2(n6363), .IN3(n6542), .QN(n6537) );
  MUX21X1 U6433 ( .IN1(n6543), .IN2(n6544), .S(\i_m4stg_frac/n1519 ), .Q(n6542) );
  XNOR2X1 U6434 ( .IN1(n1038), .IN2(n907), .Q(n6363) );
  XNOR3X1 U6435 ( .IN1(n6510), .IN2(n6411), .IN3(n6511), .Q(n6506) );
  AO21X1 U6436 ( .IN1(n6545), .IN2(n6516), .IN3(n6517), .Q(n6511) );
  INVX0 U6437 ( .INP(n6414), .ZN(n6411) );
  XOR2X1 U6438 ( .IN1(n6515), .IN2(n6546), .Q(n6510) );
  AOI21X1 U6439 ( .IN1(\i_m4stg_frac/n1464 ), .IN2(n6248), .IN3(n6464), .QN(
        n6515) );
  NOR2X0 U6440 ( .IN1(\i_m4stg_frac/n1464 ), .IN2(n6248), .QN(n6464) );
  NAND2X0 U6441 ( .IN1(n6503), .IN2(n6504), .QN(n6533) );
  AO22X1 U6442 ( .IN1(n6104), .IN2(n6105), .IN3(n6547), .IN4(n6103), .Q(
        \i_m4stg_frac/a0cout[64] ) );
  AO22X1 U6443 ( .IN1(n6548), .IN2(n6549), .IN3(n6550), .IN4(n6551), .Q(n6103)
         );
  OR2X1 U6444 ( .IN1(n6548), .IN2(n6549), .Q(n6551) );
  OR2X1 U6445 ( .IN1(n6105), .IN2(n6104), .Q(n6547) );
  INVX0 U6446 ( .INP(n6552), .ZN(n6105) );
  MUX21X1 U6447 ( .IN1(n6553), .IN2(n6554), .S(n6555), .Q(n6552) );
  INVX0 U6448 ( .INP(n6556), .ZN(n6555) );
  XNOR2X1 U6449 ( .IN1(n6529), .IN2(n6526), .Q(n6104) );
  AOI21X1 U6450 ( .IN1(n6557), .IN2(n6558), .IN3(n6559), .QN(n6526) );
  XNOR3X1 U6451 ( .IN1(n6522), .IN2(n6523), .IN3(n6560), .Q(n6529) );
  XOR2X1 U6452 ( .IN1(n6527), .IN2(n6521), .Q(n6560) );
  XOR2X1 U6453 ( .IN1(n6504), .IN2(n6503), .Q(n6521) );
  NAND2X0 U6454 ( .IN1(n6561), .IN2(n6562), .QN(n6503) );
  MUX21X1 U6455 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1517 ), .Q(n6562) );
  MUX21X1 U6456 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1516 ), .Q(n6561) );
  NAND2X0 U6457 ( .IN1(n6563), .IN2(n6564), .QN(n6504) );
  MUX21X1 U6458 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1519 ), .Q(n6564) );
  MUX21X1 U6459 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1518 ), .Q(n6563) );
  XOR3X1 U6460 ( .IN1(n6532), .IN2(n6414), .IN3(n6530), .Q(n6527) );
  XOR2X1 U6461 ( .IN1(n6545), .IN2(n6546), .Q(n6530) );
  AO21X1 U6462 ( .IN1(n6568), .IN2(n6569), .IN3(n6570), .Q(n6545) );
  XOR2X1 U6463 ( .IN1(n6571), .IN2(n6405), .Q(n6414) );
  NOR2X0 U6464 ( .IN1(n6536), .IN2(n6394), .QN(n6405) );
  NOR2X0 U6465 ( .IN1(n6572), .IN2(n6376), .QN(n6394) );
  NOR2X0 U6466 ( .IN1(n6397), .IN2(n6386), .QN(n6536) );
  NOR2X0 U6467 ( .IN1(n6573), .IN2(n6574), .QN(n6523) );
  AO22X1 U6468 ( .IN1(n6535), .IN2(n6397), .IN3(n6575), .IN4(n6576), .Q(n6522)
         );
  AO22X1 U6469 ( .IN1(n6577), .IN2(n6578), .IN3(n6579), .IN4(n6107), .Q(
        \i_m4stg_frac/a0cout[63] ) );
  AO22X1 U6470 ( .IN1(n6580), .IN2(n6581), .IN3(n6582), .IN4(n6583), .Q(n6107)
         );
  OR2X1 U6471 ( .IN1(n6580), .IN2(n6581), .Q(n6583) );
  NAND2X0 U6472 ( .IN1(n6108), .IN2(n6106), .QN(n6579) );
  INVX0 U6473 ( .INP(n6577), .ZN(n6106) );
  INVX0 U6474 ( .INP(n6108), .ZN(n6578) );
  MUX21X1 U6475 ( .IN1(n6584), .IN2(n6585), .S(n6586), .Q(n6108) );
  INVX0 U6476 ( .INP(n6587), .ZN(n6586) );
  XOR2X1 U6477 ( .IN1(n6556), .IN2(n6554), .Q(n6577) );
  AOI21X1 U6478 ( .IN1(n6588), .IN2(n6558), .IN3(n6559), .QN(n6554) );
  XNOR3X1 U6479 ( .IN1(n6549), .IN2(n6550), .IN3(n6589), .Q(n6556) );
  XNOR2X1 U6480 ( .IN1(n6553), .IN2(n6548), .Q(n6589) );
  XOR2X1 U6481 ( .IN1(n6573), .IN2(n6574), .Q(n6548) );
  AND2X1 U6482 ( .IN1(n6590), .IN2(n6591), .Q(n6574) );
  MUX21X1 U6483 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1516 ), .Q(n6591) );
  MUX21X1 U6484 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1515 ), .Q(n6590) );
  AND2X1 U6485 ( .IN1(n6592), .IN2(n6593), .Q(n6573) );
  MUX21X1 U6486 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1518 ), .Q(n6593) );
  MUX21X1 U6487 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1517 ), .Q(n6592) );
  XNOR2X1 U6488 ( .IN1(n6557), .IN2(n6594), .Q(n6553) );
  XOR2X1 U6489 ( .IN1(n6595), .IN2(n6575), .Q(n6557) );
  OAI21X1 U6490 ( .IN1(n6376), .IN2(n951), .IN3(n6596), .QN(n6575) );
  MUX21X1 U6491 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1519 ), .Q(n6596) );
  INVX0 U6492 ( .INP(n6386), .ZN(n6376) );
  OA21X1 U6493 ( .IN1(n907), .IN2(\i_m4stg_frac/n1004 ), .IN3(n6373), .Q(n6386) );
  OA21X1 U6494 ( .IN1(n936), .IN2(\i_m4stg_frac/n1530 ), .IN3(n1145), .Q(n6373) );
  NOR2X0 U6495 ( .IN1(n6599), .IN2(n6600), .QN(n6550) );
  AO22X1 U6496 ( .IN1(n6535), .IN2(n6397), .IN3(n6601), .IN4(n6576), .Q(n6549)
         );
  INVX0 U6497 ( .INP(n6572), .ZN(n6397) );
  AO22X1 U6498 ( .IN1(n6602), .IN2(n6603), .IN3(n6604), .IN4(n6110), .Q(
        \i_m4stg_frac/a0cout[62] ) );
  AO22X1 U6499 ( .IN1(n6605), .IN2(n6606), .IN3(n6607), .IN4(n6608), .Q(n6110)
         );
  OR2X1 U6500 ( .IN1(n6605), .IN2(n6606), .Q(n6608) );
  NAND2X0 U6501 ( .IN1(n6111), .IN2(n6109), .QN(n6604) );
  INVX0 U6502 ( .INP(n6602), .ZN(n6109) );
  INVX0 U6503 ( .INP(n6111), .ZN(n6603) );
  MUX21X1 U6504 ( .IN1(n6609), .IN2(n6610), .S(n6611), .Q(n6111) );
  INVX0 U6505 ( .INP(n6612), .ZN(n6611) );
  XOR2X1 U6506 ( .IN1(n6587), .IN2(n6585), .Q(n6602) );
  AOI21X1 U6507 ( .IN1(n6613), .IN2(n6558), .IN3(n6559), .QN(n6585) );
  XNOR3X1 U6508 ( .IN1(n6581), .IN2(n6582), .IN3(n6614), .Q(n6587) );
  XNOR2X1 U6509 ( .IN1(n6584), .IN2(n6580), .Q(n6614) );
  XOR2X1 U6510 ( .IN1(n6599), .IN2(n6600), .Q(n6580) );
  AND2X1 U6511 ( .IN1(n6615), .IN2(n6616), .Q(n6600) );
  MUX21X1 U6512 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1515 ), .Q(n6616) );
  MUX21X1 U6513 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1514 ), .Q(n6615) );
  AND2X1 U6514 ( .IN1(n6617), .IN2(n6618), .Q(n6599) );
  MUX21X1 U6515 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1517 ), .Q(n6618) );
  MUX21X1 U6516 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1516 ), .Q(n6617) );
  XNOR2X1 U6517 ( .IN1(n6588), .IN2(n6594), .Q(n6584) );
  XOR2X1 U6518 ( .IN1(n6601), .IN2(n6595), .Q(n6588) );
  OA21X1 U6519 ( .IN1(n6571), .IN2(n6572), .IN3(n6576), .Q(n6595) );
  NAND2X0 U6520 ( .IN1(n6571), .IN2(n6572), .QN(n6576) );
  NAND2X0 U6521 ( .IN1(n6619), .IN2(n6620), .QN(n6601) );
  MUX21X1 U6522 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1518 ), .Q(n6620) );
  MUX21X1 U6523 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1519 ), .Q(n6619) );
  NOR2X0 U6524 ( .IN1(n6623), .IN2(n6624), .QN(n6582) );
  AO22X1 U6525 ( .IN1(n6625), .IN2(n6626), .IN3(n6535), .IN4(n6627), .Q(n6581)
         );
  OR2X1 U6526 ( .IN1(n6626), .IN2(n6625), .Q(n6627) );
  AO22X1 U6527 ( .IN1(n6113), .IN2(n6114), .IN3(n6628), .IN4(n6112), .Q(
        \i_m4stg_frac/a0cout[61] ) );
  AO22X1 U6528 ( .IN1(n6629), .IN2(n6630), .IN3(n6631), .IN4(n6632), .Q(n6112)
         );
  OR2X1 U6529 ( .IN1(n6629), .IN2(n6630), .Q(n6632) );
  OR2X1 U6530 ( .IN1(n6114), .IN2(n6113), .Q(n6628) );
  INVX0 U6531 ( .INP(n6633), .ZN(n6114) );
  MUX21X1 U6532 ( .IN1(n6634), .IN2(n6635), .S(n6636), .Q(n6633) );
  INVX0 U6533 ( .INP(n6637), .ZN(n6636) );
  XNOR2X1 U6534 ( .IN1(n6612), .IN2(n6609), .Q(n6113) );
  AOI21X1 U6535 ( .IN1(n6638), .IN2(n6558), .IN3(n6559), .QN(n6609) );
  XOR3X1 U6536 ( .IN1(n6639), .IN2(n6605), .IN3(n6610), .Q(n6612) );
  XNOR2X1 U6537 ( .IN1(n6613), .IN2(n6594), .Q(n6610) );
  XOR3X1 U6538 ( .IN1(n6625), .IN2(n6535), .IN3(n6626), .Q(n6613) );
  NAND2X0 U6539 ( .IN1(n6640), .IN2(n6641), .QN(n6626) );
  MUX21X1 U6540 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1517 ), .Q(n6641) );
  MUX21X1 U6541 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1518 ), .Q(n6640) );
  OAI21X1 U6542 ( .IN1(n6572), .IN2(n915), .IN3(n6642), .QN(n6625) );
  MUX21X1 U6543 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1519 ), .Q(n6642) );
  NAND2X0 U6544 ( .IN1(n6645), .IN2(n1118), .QN(n6572) );
  XOR2X1 U6545 ( .IN1(\i_m4stg_frac/n1007 ), .IN2(n907), .Q(n6645) );
  XOR2X1 U6546 ( .IN1(n6623), .IN2(n6624), .Q(n6605) );
  AND2X1 U6547 ( .IN1(n6646), .IN2(n6647), .Q(n6624) );
  MUX21X1 U6548 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1514 ), .Q(n6647) );
  MUX21X1 U6549 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1513 ), .Q(n6646) );
  AND2X1 U6550 ( .IN1(n6648), .IN2(n6649), .Q(n6623) );
  MUX21X1 U6551 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1516 ), .Q(n6649) );
  MUX21X1 U6552 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1515 ), .Q(n6648) );
  XNOR2X1 U6553 ( .IN1(n6606), .IN2(n6607), .Q(n6639) );
  NOR2X0 U6554 ( .IN1(n6650), .IN2(n6651), .QN(n6607) );
  AO22X1 U6555 ( .IN1(n6535), .IN2(n6652), .IN3(n6653), .IN4(n6654), .Q(n6606)
         );
  OR2X1 U6556 ( .IN1(n6652), .IN2(n6535), .Q(n6653) );
  INVX0 U6557 ( .INP(n6571), .ZN(n6535) );
  AO22X1 U6558 ( .IN1(n6116), .IN2(n6117), .IN3(n6655), .IN4(n6115), .Q(
        \i_m4stg_frac/a0cout[60] ) );
  AO22X1 U6559 ( .IN1(n6656), .IN2(n6657), .IN3(n6658), .IN4(n6659), .Q(n6115)
         );
  OR2X1 U6560 ( .IN1(n6656), .IN2(n6657), .Q(n6659) );
  AND2X1 U6561 ( .IN1(n6660), .IN2(n6661), .Q(n6658) );
  OR2X1 U6562 ( .IN1(n6117), .IN2(n6116), .Q(n6655) );
  INVX0 U6563 ( .INP(n6662), .ZN(n6117) );
  MUX21X1 U6564 ( .IN1(n6663), .IN2(n6664), .S(n6665), .Q(n6662) );
  INVX0 U6565 ( .INP(n6666), .ZN(n6665) );
  XNOR2X1 U6566 ( .IN1(n6637), .IN2(n6634), .Q(n6116) );
  AOI21X1 U6567 ( .IN1(n6667), .IN2(n6558), .IN3(n6559), .QN(n6634) );
  INVX0 U6568 ( .INP(n6668), .ZN(n6558) );
  XOR3X1 U6569 ( .IN1(n6669), .IN2(n6629), .IN3(n6635), .Q(n6637) );
  XNOR2X1 U6570 ( .IN1(n6638), .IN2(n6594), .Q(n6635) );
  XNOR3X1 U6571 ( .IN1(n6654), .IN2(n6652), .IN3(n6571), .Q(n6638) );
  NAND2X0 U6572 ( .IN1(n6417), .IN2(n1169), .QN(n6571) );
  NAND2X0 U6573 ( .IN1(n6670), .IN2(n6671), .QN(n6652) );
  MUX21X1 U6574 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1518 ), .Q(n6671) );
  MUX21X1 U6575 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1519 ), .Q(n6670) );
  NAND2X0 U6576 ( .IN1(n6672), .IN2(n6673), .QN(n6654) );
  MUX21X1 U6577 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1516 ), .Q(n6673) );
  MUX21X1 U6578 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1517 ), .Q(n6672) );
  XOR2X1 U6579 ( .IN1(n6650), .IN2(n6651), .Q(n6629) );
  AND2X1 U6580 ( .IN1(n6674), .IN2(n6675), .Q(n6651) );
  MUX21X1 U6581 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1513 ), .Q(n6675) );
  MUX21X1 U6582 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1512 ), .Q(n6674) );
  AND2X1 U6583 ( .IN1(n6676), .IN2(n6677), .Q(n6650) );
  MUX21X1 U6584 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1515 ), .Q(n6677) );
  MUX21X1 U6585 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1514 ), .Q(n6676) );
  XNOR2X1 U6586 ( .IN1(n6630), .IN2(n6631), .Q(n6669) );
  NOR2X0 U6587 ( .IN1(n6678), .IN2(n6679), .QN(n6631) );
  AO22X1 U6588 ( .IN1(n6680), .IN2(n6681), .IN3(n6682), .IN4(n6683), .Q(n6630)
         );
  OR2X1 U6589 ( .IN1(n6680), .IN2(n6681), .Q(n6682) );
  NOR2X0 U6590 ( .IN1(n6119), .IN2(n6118), .QN(\i_m4stg_frac/a0cout[5] ) );
  XOR3X1 U6591 ( .IN1(n6324), .IN2(n6435), .IN3(n6436), .Q(n6118) );
  XOR3X1 U6592 ( .IN1(n6430), .IN2(n6431), .IN3(n6433), .Q(n6436) );
  NAND2X0 U6593 ( .IN1(n6684), .IN2(n6685), .QN(n6433) );
  MUX21X1 U6594 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1468 ), .Q(n6685) );
  MUX21X1 U6595 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1467 ), .Q(n6684) );
  NAND2X0 U6596 ( .IN1(n6686), .IN2(n6687), .QN(n6431) );
  MUX21X1 U6597 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1472 ), .Q(n6687) );
  MUX21X1 U6598 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1471 ), .Q(n6686) );
  NAND2X0 U6599 ( .IN1(n6688), .IN2(n6689), .QN(n6430) );
  MUX21X1 U6600 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1470 ), .Q(n6689) );
  MUX21X1 U6601 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1469 ), .Q(n6688) );
  AO22X1 U6602 ( .IN1(n6690), .IN2(n6691), .IN3(n6692), .IN4(n6693), .Q(n6435)
         );
  OR2X1 U6603 ( .IN1(n6691), .IN2(n6690), .Q(n6692) );
  AOI22X1 U6604 ( .IN1(n6694), .IN2(n6695), .IN3(n6696), .IN4(n6697), .QN(
        n6119) );
  OR2X1 U6605 ( .IN1(n6695), .IN2(n6694), .Q(n6697) );
  AO22X1 U6606 ( .IN1(n6698), .IN2(n6699), .IN3(n6700), .IN4(n6121), .Q(
        \i_m4stg_frac/a0cout[59] ) );
  AO22X1 U6607 ( .IN1(n6701), .IN2(n6702), .IN3(n6703), .IN4(n6704), .Q(n6121)
         );
  OR2X1 U6608 ( .IN1(n6701), .IN2(n6702), .Q(n6704) );
  AND2X1 U6609 ( .IN1(n6705), .IN2(n6706), .Q(n6703) );
  NAND2X0 U6610 ( .IN1(n6122), .IN2(n6120), .QN(n6700) );
  INVX0 U6611 ( .INP(n6698), .ZN(n6120) );
  INVX0 U6612 ( .INP(n6122), .ZN(n6699) );
  MUX21X1 U6613 ( .IN1(n6707), .IN2(n6708), .S(n6709), .Q(n6122) );
  INVX0 U6614 ( .INP(n6710), .ZN(n6709) );
  XOR2X1 U6615 ( .IN1(n6666), .IN2(n6664), .Q(n6698) );
  AOI22X1 U6616 ( .IN1(n6711), .IN2(n6712), .IN3(n6713), .IN4(n6714), .QN(
        n6664) );
  OR2X1 U6617 ( .IN1(n6712), .IN2(n6711), .Q(n6714) );
  XNOR3X1 U6618 ( .IN1(n6715), .IN2(n6656), .IN3(n6663), .Q(n6666) );
  XNOR2X1 U6619 ( .IN1(n6667), .IN2(n6594), .Q(n6663) );
  NOR2X0 U6620 ( .IN1(n6668), .IN2(n6559), .QN(n6594) );
  AND2X1 U6621 ( .IN1(n6711), .IN2(n6532), .Q(n6559) );
  NOR2X0 U6622 ( .IN1(n6532), .IN2(n6711), .QN(n6668) );
  AO21X1 U6623 ( .IN1(n6716), .IN2(n6516), .IN3(n6517), .Q(n6532) );
  INVX0 U6624 ( .INP(n6717), .ZN(n6516) );
  XOR3X1 U6625 ( .IN1(n6683), .IN2(n6681), .IN3(n6680), .Q(n6667) );
  NAND2X0 U6626 ( .IN1(n6718), .IN2(n6719), .QN(n6680) );
  MUX21X1 U6627 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1518 ), .Q(n6719) );
  MUX21X1 U6628 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1517 ), .Q(n6718) );
  AO21X1 U6629 ( .IN1(n6417), .IN2(n6351), .IN3(n6720), .Q(n6681) );
  INVX0 U6630 ( .INP(n6721), .ZN(n6720) );
  MUX21X1 U6631 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1519 ), .Q(n6721) );
  XOR2X1 U6632 ( .IN1(n913), .IN2(\i_m4stg_frac/n1530 ), .Q(n6417) );
  NAND2X0 U6633 ( .IN1(n6722), .IN2(n6723), .QN(n6683) );
  MUX21X1 U6634 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1515 ), .Q(n6723) );
  MUX21X1 U6635 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1516 ), .Q(n6722) );
  XOR2X1 U6636 ( .IN1(n6678), .IN2(n6679), .Q(n6656) );
  AND2X1 U6637 ( .IN1(n6724), .IN2(n6725), .Q(n6679) );
  MUX21X1 U6638 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1512 ), .Q(n6725) );
  MUX21X1 U6639 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1511 ), .Q(n6724) );
  AND2X1 U6640 ( .IN1(n6726), .IN2(n6727), .Q(n6678) );
  MUX21X1 U6641 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1514 ), .Q(n6727) );
  MUX21X1 U6642 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1513 ), .Q(n6726) );
  XOR2X1 U6643 ( .IN1(n6657), .IN2(n6728), .Q(n6715) );
  NAND2X0 U6644 ( .IN1(n6660), .IN2(n6661), .QN(n6728) );
  AO22X1 U6645 ( .IN1(n6729), .IN2(n6730), .IN3(n6731), .IN4(n6732), .Q(n6657)
         );
  OR2X1 U6646 ( .IN1(n6730), .IN2(n6729), .Q(n6731) );
  AO22X1 U6647 ( .IN1(n6124), .IN2(n6125), .IN3(n6733), .IN4(n6123), .Q(
        \i_m4stg_frac/a0cout[58] ) );
  AO22X1 U6648 ( .IN1(n6734), .IN2(n6735), .IN3(n6736), .IN4(n6737), .Q(n6123)
         );
  OR2X1 U6649 ( .IN1(n6734), .IN2(n6735), .Q(n6737) );
  AND2X1 U6650 ( .IN1(n6738), .IN2(n6739), .Q(n6736) );
  OR2X1 U6651 ( .IN1(n6125), .IN2(n6124), .Q(n6733) );
  INVX0 U6652 ( .INP(n6740), .ZN(n6125) );
  MUX21X1 U6653 ( .IN1(n6741), .IN2(n6742), .S(n6743), .Q(n6740) );
  INVX0 U6654 ( .INP(n6744), .ZN(n6743) );
  XNOR2X1 U6655 ( .IN1(n6710), .IN2(n6707), .Q(n6124) );
  AOI22X1 U6656 ( .IN1(n6745), .IN2(n6746), .IN3(n6747), .IN4(n6748), .QN(
        n6707) );
  OR2X1 U6657 ( .IN1(n6746), .IN2(n6745), .Q(n6748) );
  XOR3X1 U6658 ( .IN1(n6749), .IN2(n6701), .IN3(n6708), .Q(n6710) );
  XNOR3X1 U6659 ( .IN1(n6712), .IN2(n6711), .IN3(n6713), .Q(n6708) );
  XOR3X1 U6660 ( .IN1(n6729), .IN2(n6730), .IN3(n6732), .Q(n6713) );
  NAND2X0 U6661 ( .IN1(n6750), .IN2(n6751), .QN(n6732) );
  MUX21X1 U6662 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1514 ), .Q(n6751) );
  MUX21X1 U6663 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1515 ), .Q(n6750) );
  NAND2X0 U6664 ( .IN1(n6752), .IN2(n6753), .QN(n6730) );
  MUX21X1 U6665 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1518 ), .Q(n6753) );
  MUX21X1 U6666 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1519 ), .Q(n6752) );
  NAND2X0 U6667 ( .IN1(n6754), .IN2(n6755), .QN(n6729) );
  MUX21X1 U6668 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1516 ), .Q(n6755) );
  MUX21X1 U6669 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1517 ), .Q(n6754) );
  XNOR2X1 U6670 ( .IN1(n6756), .IN2(n6546), .Q(n6711) );
  NOR2X0 U6671 ( .IN1(n6717), .IN2(n6517), .QN(n6546) );
  NOR2X0 U6672 ( .IN1(n6514), .IN2(n6495), .QN(n6517) );
  NOR2X0 U6673 ( .IN1(n6757), .IN2(n6463), .QN(n6717) );
  AO22X1 U6674 ( .IN1(n6716), .IN2(n6757), .IN3(n6758), .IN4(n6759), .Q(n6712)
         );
  XOR2X1 U6675 ( .IN1(n6661), .IN2(n6660), .Q(n6701) );
  NAND2X0 U6676 ( .IN1(n6760), .IN2(n6761), .QN(n6660) );
  MUX21X1 U6677 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1511 ), .Q(n6761) );
  MUX21X1 U6678 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1510 ), .Q(n6760) );
  NAND2X0 U6679 ( .IN1(n6762), .IN2(n6763), .QN(n6661) );
  MUX21X1 U6680 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1513 ), .Q(n6763) );
  MUX21X1 U6681 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1512 ), .Q(n6762) );
  XOR2X1 U6682 ( .IN1(n6702), .IN2(n6764), .Q(n6749) );
  NAND2X0 U6683 ( .IN1(n6705), .IN2(n6706), .QN(n6764) );
  AO22X1 U6684 ( .IN1(n6765), .IN2(n6766), .IN3(n6767), .IN4(n6768), .Q(n6702)
         );
  OR2X1 U6685 ( .IN1(n6765), .IN2(n6766), .Q(n6767) );
  AO22X1 U6686 ( .IN1(n6769), .IN2(n6770), .IN3(n6771), .IN4(n6127), .Q(
        \i_m4stg_frac/a0cout[57] ) );
  AO22X1 U6687 ( .IN1(n6772), .IN2(n6773), .IN3(n6774), .IN4(n6775), .Q(n6127)
         );
  OR2X1 U6688 ( .IN1(n6772), .IN2(n6773), .Q(n6775) );
  AND2X1 U6689 ( .IN1(n6776), .IN2(n6777), .Q(n6774) );
  NAND2X0 U6690 ( .IN1(n6128), .IN2(n6126), .QN(n6771) );
  INVX0 U6691 ( .INP(n6769), .ZN(n6126) );
  INVX0 U6692 ( .INP(n6128), .ZN(n6770) );
  MUX21X1 U6693 ( .IN1(n6778), .IN2(n6779), .S(n6780), .Q(n6128) );
  INVX0 U6694 ( .INP(n6781), .ZN(n6780) );
  XOR2X1 U6695 ( .IN1(n6744), .IN2(n6742), .Q(n6769) );
  AOI22X1 U6696 ( .IN1(n6782), .IN2(n6783), .IN3(n6784), .IN4(n6785), .QN(
        n6742) );
  OR2X1 U6697 ( .IN1(n6783), .IN2(n6782), .Q(n6785) );
  XNOR3X1 U6698 ( .IN1(n6786), .IN2(n6734), .IN3(n6741), .Q(n6744) );
  XNOR3X1 U6699 ( .IN1(n6746), .IN2(n6745), .IN3(n6747), .Q(n6741) );
  XOR3X1 U6700 ( .IN1(n6765), .IN2(n6766), .IN3(n6768), .Q(n6747) );
  NAND2X0 U6701 ( .IN1(n6787), .IN2(n6788), .QN(n6768) );
  MUX21X1 U6702 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1513 ), .Q(n6788) );
  MUX21X1 U6703 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1514 ), .Q(n6787) );
  NAND2X0 U6704 ( .IN1(n6789), .IN2(n6790), .QN(n6766) );
  MUX21X1 U6705 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1518 ), .Q(n6790) );
  MUX21X1 U6706 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1517 ), .Q(n6789) );
  NAND2X0 U6707 ( .IN1(n6791), .IN2(n6792), .QN(n6765) );
  MUX21X1 U6708 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1515 ), .Q(n6792) );
  MUX21X1 U6709 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1516 ), .Q(n6791) );
  XOR2X1 U6710 ( .IN1(n6793), .IN2(n6758), .Q(n6745) );
  OAI21X1 U6711 ( .IN1(n6495), .IN2(n950), .IN3(n6794), .QN(n6758) );
  MUX21X1 U6712 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1519 ), .Q(n6794) );
  INVX0 U6713 ( .INP(n6463), .ZN(n6495) );
  OA21X1 U6714 ( .IN1(n907), .IN2(\i_m4stg_frac/n1013 ), .IN3(n6468), .Q(n6463) );
  OA21X1 U6715 ( .IN1(n935), .IN2(\i_m4stg_frac/n1530 ), .IN3(n1144), .Q(n6468) );
  AO22X1 U6716 ( .IN1(n6716), .IN2(n6757), .IN3(n6795), .IN4(n6759), .Q(n6746)
         );
  INVX0 U6717 ( .INP(n6514), .ZN(n6757) );
  XOR2X1 U6718 ( .IN1(n6706), .IN2(n6705), .Q(n6734) );
  NAND2X0 U6719 ( .IN1(n6796), .IN2(n6797), .QN(n6705) );
  MUX21X1 U6720 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1510 ), .Q(n6797) );
  MUX21X1 U6721 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1509 ), .Q(n6796) );
  NAND2X0 U6722 ( .IN1(n6798), .IN2(n6799), .QN(n6706) );
  MUX21X1 U6723 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1512 ), .Q(n6799) );
  MUX21X1 U6724 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1511 ), .Q(n6798) );
  XOR2X1 U6725 ( .IN1(n6735), .IN2(n6800), .Q(n6786) );
  NAND2X0 U6726 ( .IN1(n6738), .IN2(n6739), .QN(n6800) );
  AO22X1 U6727 ( .IN1(n6801), .IN2(n6802), .IN3(n6803), .IN4(n6804), .Q(n6735)
         );
  OR2X1 U6728 ( .IN1(n6802), .IN2(n6801), .Q(n6803) );
  AO22X1 U6729 ( .IN1(n6130), .IN2(n6131), .IN3(n6805), .IN4(n6129), .Q(
        \i_m4stg_frac/a0cout[56] ) );
  AO22X1 U6730 ( .IN1(n6806), .IN2(n6807), .IN3(n6808), .IN4(n6809), .Q(n6129)
         );
  OR2X1 U6731 ( .IN1(n6806), .IN2(n6807), .Q(n6809) );
  AND2X1 U6732 ( .IN1(n6810), .IN2(n6811), .Q(n6808) );
  OR2X1 U6733 ( .IN1(n6131), .IN2(n6130), .Q(n6805) );
  INVX0 U6734 ( .INP(n6812), .ZN(n6131) );
  MUX21X1 U6735 ( .IN1(n6813), .IN2(n6814), .S(n6815), .Q(n6812) );
  INVX0 U6736 ( .INP(n6816), .ZN(n6815) );
  XOR2X1 U6737 ( .IN1(n6781), .IN2(n6779), .Q(n6130) );
  AOI22X1 U6738 ( .IN1(n6817), .IN2(n6818), .IN3(n6819), .IN4(n6820), .QN(
        n6779) );
  OR2X1 U6739 ( .IN1(n6818), .IN2(n6817), .Q(n6820) );
  XNOR3X1 U6740 ( .IN1(n6821), .IN2(n6772), .IN3(n6778), .Q(n6781) );
  XNOR3X1 U6741 ( .IN1(n6783), .IN2(n6782), .IN3(n6784), .Q(n6778) );
  XOR3X1 U6742 ( .IN1(n6801), .IN2(n6802), .IN3(n6804), .Q(n6784) );
  NAND2X0 U6743 ( .IN1(n6822), .IN2(n6823), .QN(n6804) );
  MUX21X1 U6744 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1512 ), .Q(n6823) );
  MUX21X1 U6745 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1513 ), .Q(n6822) );
  NAND2X0 U6746 ( .IN1(n6824), .IN2(n6825), .QN(n6802) );
  MUX21X1 U6747 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1517 ), .Q(n6825) );
  MUX21X1 U6748 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1516 ), .Q(n6824) );
  NAND2X0 U6749 ( .IN1(n6826), .IN2(n6827), .QN(n6801) );
  MUX21X1 U6750 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1514 ), .Q(n6827) );
  MUX21X1 U6751 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1515 ), .Q(n6826) );
  XOR2X1 U6752 ( .IN1(n6795), .IN2(n6793), .Q(n6782) );
  OA21X1 U6753 ( .IN1(n6756), .IN2(n6514), .IN3(n6759), .Q(n6793) );
  NAND2X0 U6754 ( .IN1(n6756), .IN2(n6514), .QN(n6759) );
  INVX0 U6755 ( .INP(n6716), .ZN(n6756) );
  NAND2X0 U6756 ( .IN1(n6828), .IN2(n6829), .QN(n6795) );
  MUX21X1 U6757 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1518 ), .Q(n6829) );
  MUX21X1 U6758 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1519 ), .Q(n6828) );
  AO22X1 U6759 ( .IN1(n6830), .IN2(n6831), .IN3(n6716), .IN4(n6832), .Q(n6783)
         );
  OR2X1 U6760 ( .IN1(n6831), .IN2(n6830), .Q(n6832) );
  XOR2X1 U6761 ( .IN1(n6739), .IN2(n6738), .Q(n6772) );
  NAND2X0 U6762 ( .IN1(n6833), .IN2(n6834), .QN(n6738) );
  MUX21X1 U6763 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1509 ), .Q(n6834) );
  MUX21X1 U6764 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1508 ), .Q(n6833) );
  NAND2X0 U6765 ( .IN1(n6835), .IN2(n6836), .QN(n6739) );
  MUX21X1 U6766 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1511 ), .Q(n6836) );
  MUX21X1 U6767 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1510 ), .Q(n6835) );
  XOR2X1 U6768 ( .IN1(n6773), .IN2(n6837), .Q(n6821) );
  NAND2X0 U6769 ( .IN1(n6776), .IN2(n6777), .QN(n6837) );
  AO22X1 U6770 ( .IN1(n6838), .IN2(n6839), .IN3(n6840), .IN4(n6841), .Q(n6773)
         );
  OR2X1 U6771 ( .IN1(n6839), .IN2(n6838), .Q(n6840) );
  AO22X1 U6772 ( .IN1(n6133), .IN2(n6134), .IN3(n6842), .IN4(n6132), .Q(
        \i_m4stg_frac/a0cout[55] ) );
  AO22X1 U6773 ( .IN1(n6843), .IN2(n6844), .IN3(n6845), .IN4(n6846), .Q(n6132)
         );
  OR2X1 U6774 ( .IN1(n6843), .IN2(n6844), .Q(n6846) );
  AND2X1 U6775 ( .IN1(n6847), .IN2(n6848), .Q(n6845) );
  OR2X1 U6776 ( .IN1(n6134), .IN2(n6133), .Q(n6842) );
  INVX0 U6777 ( .INP(n6849), .ZN(n6134) );
  MUX21X1 U6778 ( .IN1(n6850), .IN2(n6851), .S(n6852), .Q(n6849) );
  INVX0 U6779 ( .INP(n6853), .ZN(n6852) );
  XNOR2X1 U6780 ( .IN1(n6816), .IN2(n6813), .Q(n6133) );
  OA22X1 U6781 ( .IN1(n6854), .IN2(n6855), .IN3(n6856), .IN4(n6857), .Q(n6813)
         );
  AND2X1 U6782 ( .IN1(n6855), .IN2(n6854), .Q(n6857) );
  XOR3X1 U6783 ( .IN1(n6858), .IN2(n6806), .IN3(n6814), .Q(n6816) );
  XNOR3X1 U6784 ( .IN1(n6818), .IN2(n6817), .IN3(n6819), .Q(n6814) );
  XOR3X1 U6785 ( .IN1(n6838), .IN2(n6839), .IN3(n6841), .Q(n6819) );
  NAND2X0 U6786 ( .IN1(n6859), .IN2(n6860), .QN(n6841) );
  MUX21X1 U6787 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1511 ), .Q(n6860) );
  MUX21X1 U6788 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1512 ), .Q(n6859) );
  NAND2X0 U6789 ( .IN1(n6861), .IN2(n6862), .QN(n6839) );
  MUX21X1 U6790 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1516 ), .Q(n6862) );
  MUX21X1 U6791 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1515 ), .Q(n6861) );
  NAND2X0 U6792 ( .IN1(n6863), .IN2(n6864), .QN(n6838) );
  MUX21X1 U6793 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1513 ), .Q(n6864) );
  MUX21X1 U6794 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1514 ), .Q(n6863) );
  XOR3X1 U6795 ( .IN1(n6830), .IN2(n6716), .IN3(n6831), .Q(n6817) );
  NAND2X0 U6796 ( .IN1(n6865), .IN2(n6866), .QN(n6831) );
  MUX21X1 U6797 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1517 ), .Q(n6866) );
  MUX21X1 U6798 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1518 ), .Q(n6865) );
  OAI21X1 U6799 ( .IN1(n6514), .IN2(n1135), .IN3(n6867), .QN(n6830) );
  MUX21X1 U6800 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1519 ), .Q(n6867) );
  NAND2X0 U6801 ( .IN1(n6868), .IN2(n933), .QN(n6514) );
  XOR2X1 U6802 ( .IN1(\i_m4stg_frac/n1016 ), .IN2(n907), .Q(n6868) );
  AO22X1 U6803 ( .IN1(n6716), .IN2(n6869), .IN3(n6870), .IN4(n6871), .Q(n6818)
         );
  OR2X1 U6804 ( .IN1(n6869), .IN2(n6716), .Q(n6870) );
  XOR2X1 U6805 ( .IN1(n6777), .IN2(n6776), .Q(n6806) );
  NAND2X0 U6806 ( .IN1(n6872), .IN2(n6873), .QN(n6776) );
  MUX21X1 U6807 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1508 ), .Q(n6873) );
  MUX21X1 U6808 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1507 ), .Q(n6872) );
  NAND2X0 U6809 ( .IN1(n6874), .IN2(n6875), .QN(n6777) );
  MUX21X1 U6810 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1510 ), .Q(n6875) );
  MUX21X1 U6811 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1509 ), .Q(n6874) );
  XOR2X1 U6812 ( .IN1(n6807), .IN2(n6876), .Q(n6858) );
  NAND2X0 U6813 ( .IN1(n6810), .IN2(n6811), .QN(n6876) );
  AO22X1 U6814 ( .IN1(n6877), .IN2(n6878), .IN3(n6879), .IN4(n6880), .Q(n6807)
         );
  OR2X1 U6815 ( .IN1(n6877), .IN2(n6878), .Q(n6879) );
  AO22X1 U6816 ( .IN1(n6136), .IN2(n6137), .IN3(n6881), .IN4(n6135), .Q(
        \i_m4stg_frac/a0cout[54] ) );
  AO22X1 U6817 ( .IN1(n6882), .IN2(n6883), .IN3(n6884), .IN4(n6885), .Q(n6135)
         );
  OR2X1 U6818 ( .IN1(n6882), .IN2(n6883), .Q(n6885) );
  AND2X1 U6819 ( .IN1(n6886), .IN2(n6887), .Q(n6884) );
  OR2X1 U6820 ( .IN1(n6137), .IN2(n6136), .Q(n6881) );
  INVX0 U6821 ( .INP(n6888), .ZN(n6137) );
  MUX21X1 U6822 ( .IN1(n6889), .IN2(n6890), .S(n6891), .Q(n6888) );
  INVX0 U6823 ( .INP(n6892), .ZN(n6891) );
  XNOR2X1 U6824 ( .IN1(n6853), .IN2(n6850), .Q(n6136) );
  OA22X1 U6825 ( .IN1(n6893), .IN2(n6894), .IN3(n6895), .IN4(n6896), .Q(n6850)
         );
  AND2X1 U6826 ( .IN1(n6894), .IN2(n6893), .Q(n6896) );
  XOR3X1 U6827 ( .IN1(n6897), .IN2(n6843), .IN3(n6851), .Q(n6853) );
  XOR3X1 U6828 ( .IN1(n6856), .IN2(n6855), .IN3(n6854), .Q(n6851) );
  XNOR3X1 U6829 ( .IN1(n6871), .IN2(n6869), .IN3(n6716), .Q(n6854) );
  NOR2X0 U6830 ( .IN1(n6898), .IN2(\i_m4stg_frac/n1020 ), .QN(n6716) );
  NAND2X0 U6831 ( .IN1(n6899), .IN2(n6900), .QN(n6869) );
  MUX21X1 U6832 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1518 ), .Q(n6900) );
  MUX21X1 U6833 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1519 ), .Q(n6899) );
  NAND2X0 U6834 ( .IN1(n6901), .IN2(n6902), .QN(n6871) );
  MUX21X1 U6835 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1516 ), .Q(n6902) );
  MUX21X1 U6836 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1517 ), .Q(n6901) );
  AOI22X1 U6837 ( .IN1(n6903), .IN2(n6904), .IN3(n6905), .IN4(n6906), .QN(
        n6855) );
  OR2X1 U6838 ( .IN1(n6904), .IN2(n6903), .Q(n6905) );
  XNOR3X1 U6839 ( .IN1(n6877), .IN2(n6878), .IN3(n6880), .Q(n6856) );
  NAND2X0 U6840 ( .IN1(n6907), .IN2(n6908), .QN(n6880) );
  MUX21X1 U6841 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1510 ), .Q(n6908) );
  MUX21X1 U6842 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1511 ), .Q(n6907) );
  NAND2X0 U6843 ( .IN1(n6909), .IN2(n6910), .QN(n6878) );
  MUX21X1 U6844 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1515 ), .Q(n6910) );
  MUX21X1 U6845 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1514 ), .Q(n6909) );
  NAND2X0 U6846 ( .IN1(n6911), .IN2(n6912), .QN(n6877) );
  MUX21X1 U6847 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1512 ), .Q(n6912) );
  MUX21X1 U6848 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1513 ), .Q(n6911) );
  XOR2X1 U6849 ( .IN1(n6811), .IN2(n6810), .Q(n6843) );
  NAND2X0 U6850 ( .IN1(n6913), .IN2(n6914), .QN(n6810) );
  MUX21X1 U6851 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1507 ), .Q(n6914) );
  MUX21X1 U6852 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1506 ), .Q(n6913) );
  NAND2X0 U6853 ( .IN1(n6915), .IN2(n6916), .QN(n6811) );
  MUX21X1 U6854 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1509 ), .Q(n6916) );
  MUX21X1 U6855 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1508 ), .Q(n6915) );
  XOR2X1 U6856 ( .IN1(n6844), .IN2(n6917), .Q(n6897) );
  NAND2X0 U6857 ( .IN1(n6847), .IN2(n6848), .QN(n6917) );
  AO22X1 U6858 ( .IN1(n6918), .IN2(n6919), .IN3(n6920), .IN4(n6921), .Q(n6844)
         );
  OR2X1 U6859 ( .IN1(n6918), .IN2(n6919), .Q(n6920) );
  AO22X1 U6860 ( .IN1(n6922), .IN2(n6923), .IN3(n6924), .IN4(n6139), .Q(
        \i_m4stg_frac/a0cout[53] ) );
  AO22X1 U6861 ( .IN1(n6925), .IN2(n6926), .IN3(n6927), .IN4(n6928), .Q(n6139)
         );
  OR2X1 U6862 ( .IN1(n6925), .IN2(n6926), .Q(n6928) );
  AND2X1 U6863 ( .IN1(n6929), .IN2(n6930), .Q(n6927) );
  NAND2X0 U6864 ( .IN1(n6140), .IN2(n6138), .QN(n6924) );
  INVX0 U6865 ( .INP(n6922), .ZN(n6138) );
  INVX0 U6866 ( .INP(n6140), .ZN(n6923) );
  MUX21X1 U6867 ( .IN1(n6931), .IN2(n6932), .S(n6933), .Q(n6140) );
  INVX0 U6868 ( .INP(n6934), .ZN(n6933) );
  XOR2X1 U6869 ( .IN1(n6892), .IN2(n6890), .Q(n6922) );
  OA22X1 U6870 ( .IN1(n6935), .IN2(n6936), .IN3(n6937), .IN4(n6938), .Q(n6890)
         );
  AND2X1 U6871 ( .IN1(n6936), .IN2(n6935), .Q(n6938) );
  XNOR3X1 U6872 ( .IN1(n6939), .IN2(n6882), .IN3(n6889), .Q(n6892) );
  XOR3X1 U6873 ( .IN1(n6895), .IN2(n6894), .IN3(n6893), .Q(n6889) );
  XNOR3X1 U6874 ( .IN1(n6906), .IN2(n6904), .IN3(n6903), .Q(n6893) );
  NAND2X0 U6875 ( .IN1(n6940), .IN2(n6941), .QN(n6903) );
  MUX21X1 U6876 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1517 ), .Q(n6941) );
  MUX21X1 U6877 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1518 ), .Q(n6940) );
  OAI21X1 U6878 ( .IN1(n6898), .IN2(n6279), .IN3(n6942), .QN(n6904) );
  MUX21X1 U6879 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1519 ), .Q(n6942) );
  INVX0 U6880 ( .INP(n6568), .ZN(n6898) );
  XNOR2X1 U6881 ( .IN1(n1053), .IN2(n907), .Q(n6568) );
  NAND2X0 U6882 ( .IN1(n6943), .IN2(n6944), .QN(n6906) );
  MUX21X1 U6883 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1515 ), .Q(n6944) );
  MUX21X1 U6884 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1516 ), .Q(n6943) );
  AOI22X1 U6885 ( .IN1(n6945), .IN2(n6946), .IN3(n6947), .IN4(n6948), .QN(
        n6894) );
  OR2X1 U6886 ( .IN1(n6946), .IN2(n6945), .Q(n6947) );
  XNOR3X1 U6887 ( .IN1(n6918), .IN2(n6919), .IN3(n6921), .Q(n6895) );
  NAND2X0 U6888 ( .IN1(n6949), .IN2(n6950), .QN(n6921) );
  MUX21X1 U6889 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1509 ), .Q(n6950) );
  MUX21X1 U6890 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1510 ), .Q(n6949) );
  NAND2X0 U6891 ( .IN1(n6951), .IN2(n6952), .QN(n6919) );
  MUX21X1 U6892 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1514 ), .Q(n6952) );
  MUX21X1 U6893 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1513 ), .Q(n6951) );
  NAND2X0 U6894 ( .IN1(n6953), .IN2(n6954), .QN(n6918) );
  MUX21X1 U6895 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1511 ), .Q(n6954) );
  MUX21X1 U6896 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1512 ), .Q(n6953) );
  XOR2X1 U6897 ( .IN1(n6848), .IN2(n6847), .Q(n6882) );
  NAND2X0 U6898 ( .IN1(n6955), .IN2(n6956), .QN(n6847) );
  MUX21X1 U6899 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1506 ), .Q(n6956) );
  MUX21X1 U6900 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1505 ), .Q(n6955) );
  NAND2X0 U6901 ( .IN1(n6957), .IN2(n6958), .QN(n6848) );
  MUX21X1 U6902 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1508 ), .Q(n6958) );
  MUX21X1 U6903 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1507 ), .Q(n6957) );
  XOR2X1 U6904 ( .IN1(n6883), .IN2(n6959), .Q(n6939) );
  NAND2X0 U6905 ( .IN1(n6886), .IN2(n6887), .QN(n6959) );
  AO22X1 U6906 ( .IN1(n6960), .IN2(n6961), .IN3(n6962), .IN4(n6963), .Q(n6883)
         );
  OR2X1 U6907 ( .IN1(n6961), .IN2(n6960), .Q(n6962) );
  AO22X1 U6908 ( .IN1(n6964), .IN2(n6965), .IN3(n6966), .IN4(n6142), .Q(
        \i_m4stg_frac/a0cout[52] ) );
  AO22X1 U6909 ( .IN1(n6967), .IN2(n6968), .IN3(n6969), .IN4(n6970), .Q(n6142)
         );
  OR2X1 U6910 ( .IN1(n6967), .IN2(n6968), .Q(n6970) );
  AND2X1 U6911 ( .IN1(n6971), .IN2(n6972), .Q(n6969) );
  NAND2X0 U6912 ( .IN1(n6143), .IN2(n6141), .QN(n6966) );
  INVX0 U6913 ( .INP(n6964), .ZN(n6141) );
  INVX0 U6914 ( .INP(n6143), .ZN(n6965) );
  MUX21X1 U6915 ( .IN1(n6973), .IN2(n6974), .S(n6975), .Q(n6143) );
  INVX0 U6916 ( .INP(n6976), .ZN(n6975) );
  XOR2X1 U6917 ( .IN1(n6934), .IN2(n6932), .Q(n6964) );
  OA22X1 U6918 ( .IN1(n6977), .IN2(n6978), .IN3(n6979), .IN4(n6980), .Q(n6932)
         );
  AND2X1 U6919 ( .IN1(n6978), .IN2(n6977), .Q(n6980) );
  XNOR3X1 U6920 ( .IN1(n6981), .IN2(n6925), .IN3(n6931), .Q(n6934) );
  XOR3X1 U6921 ( .IN1(n6937), .IN2(n6936), .IN3(n6935), .Q(n6931) );
  XNOR3X1 U6922 ( .IN1(n6948), .IN2(n6946), .IN3(n6945), .Q(n6935) );
  NAND2X0 U6923 ( .IN1(n6982), .IN2(n6983), .QN(n6945) );
  MUX21X1 U6924 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1518 ), .Q(n6983) );
  MUX21X1 U6925 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1519 ), .Q(n6982) );
  NAND2X0 U6926 ( .IN1(n6984), .IN2(n6985), .QN(n6946) );
  MUX21X1 U6927 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1514 ), .Q(n6985) );
  MUX21X1 U6928 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1515 ), .Q(n6984) );
  NAND2X0 U6929 ( .IN1(n6986), .IN2(n6987), .QN(n6948) );
  MUX21X1 U6930 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1517 ), .Q(n6987) );
  MUX21X1 U6931 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1516 ), .Q(n6986) );
  AOI22X1 U6932 ( .IN1(n6988), .IN2(n6989), .IN3(n6990), .IN4(n6991), .QN(
        n6936) );
  OR2X1 U6933 ( .IN1(n6989), .IN2(n6988), .Q(n6990) );
  XNOR3X1 U6934 ( .IN1(n6960), .IN2(n6961), .IN3(n6963), .Q(n6937) );
  NAND2X0 U6935 ( .IN1(n6992), .IN2(n6993), .QN(n6963) );
  MUX21X1 U6936 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1508 ), .Q(n6993) );
  MUX21X1 U6937 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1509 ), .Q(n6992) );
  NAND2X0 U6938 ( .IN1(n6994), .IN2(n6995), .QN(n6961) );
  MUX21X1 U6939 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1513 ), .Q(n6995) );
  MUX21X1 U6940 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1512 ), .Q(n6994) );
  NAND2X0 U6941 ( .IN1(n6996), .IN2(n6997), .QN(n6960) );
  MUX21X1 U6942 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1510 ), .Q(n6997) );
  MUX21X1 U6943 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1511 ), .Q(n6996) );
  XOR2X1 U6944 ( .IN1(n6887), .IN2(n6886), .Q(n6925) );
  NAND2X0 U6945 ( .IN1(n6998), .IN2(n6999), .QN(n6886) );
  MUX21X1 U6946 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1505 ), .Q(n6999) );
  MUX21X1 U6947 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1504 ), .Q(n6998) );
  NAND2X0 U6948 ( .IN1(n7000), .IN2(n7001), .QN(n6887) );
  MUX21X1 U6949 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1507 ), .Q(n7001) );
  MUX21X1 U6950 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1506 ), .Q(n7000) );
  XOR2X1 U6951 ( .IN1(n6926), .IN2(n7002), .Q(n6981) );
  NAND2X0 U6952 ( .IN1(n6929), .IN2(n6930), .QN(n7002) );
  AO22X1 U6953 ( .IN1(n7003), .IN2(n7004), .IN3(n7005), .IN4(n7006), .Q(n6926)
         );
  OR2X1 U6954 ( .IN1(n7004), .IN2(n7003), .Q(n7005) );
  AO22X1 U6955 ( .IN1(n7007), .IN2(n7008), .IN3(n7009), .IN4(n6145), .Q(
        \i_m4stg_frac/a0cout[51] ) );
  AO22X1 U6956 ( .IN1(n7010), .IN2(n7011), .IN3(n7012), .IN4(n7013), .Q(n6145)
         );
  OR2X1 U6957 ( .IN1(n7010), .IN2(n7011), .Q(n7013) );
  AND2X1 U6958 ( .IN1(n7014), .IN2(n7015), .Q(n7012) );
  NAND2X0 U6959 ( .IN1(n6146), .IN2(n6144), .QN(n7009) );
  INVX0 U6960 ( .INP(n7007), .ZN(n6144) );
  INVX0 U6961 ( .INP(n6146), .ZN(n7008) );
  MUX21X1 U6962 ( .IN1(n7016), .IN2(n7017), .S(n7018), .Q(n6146) );
  INVX0 U6963 ( .INP(n7019), .ZN(n7018) );
  XOR2X1 U6964 ( .IN1(n6976), .IN2(n6974), .Q(n7007) );
  OA22X1 U6965 ( .IN1(n7020), .IN2(n7021), .IN3(n7022), .IN4(n7023), .Q(n6974)
         );
  AND2X1 U6966 ( .IN1(n7021), .IN2(n7020), .Q(n7023) );
  XNOR3X1 U6967 ( .IN1(n7024), .IN2(n6967), .IN3(n6973), .Q(n6976) );
  XOR3X1 U6968 ( .IN1(n6979), .IN2(n6978), .IN3(n6977), .Q(n6973) );
  XNOR3X1 U6969 ( .IN1(n6988), .IN2(n6989), .IN3(n6991), .Q(n6977) );
  NAND2X0 U6970 ( .IN1(n7025), .IN2(n7026), .QN(n6991) );
  MUX21X1 U6971 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1513 ), .Q(n7026) );
  MUX21X1 U6972 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1514 ), .Q(n7025) );
  NAND2X0 U6973 ( .IN1(n7027), .IN2(n7028), .QN(n6989) );
  MUX21X1 U6974 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1518 ), .Q(n7028) );
  MUX21X1 U6975 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1517 ), .Q(n7027) );
  NAND2X0 U6976 ( .IN1(n7029), .IN2(n7030), .QN(n6988) );
  MUX21X1 U6977 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1516 ), .Q(n7030) );
  MUX21X1 U6978 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1515 ), .Q(n7029) );
  AOI22X1 U6979 ( .IN1(n7031), .IN2(n7032), .IN3(n7033), .IN4(n7034), .QN(
        n6978) );
  OR2X1 U6980 ( .IN1(n7032), .IN2(n7031), .Q(n7033) );
  XNOR3X1 U6981 ( .IN1(n7003), .IN2(n7004), .IN3(n7006), .Q(n6979) );
  NAND2X0 U6982 ( .IN1(n7035), .IN2(n7036), .QN(n7006) );
  MUX21X1 U6983 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1507 ), .Q(n7036) );
  MUX21X1 U6984 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1508 ), .Q(n7035) );
  NAND2X0 U6985 ( .IN1(n7037), .IN2(n7038), .QN(n7004) );
  MUX21X1 U6986 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1512 ), .Q(n7038) );
  MUX21X1 U6987 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1511 ), .Q(n7037) );
  NAND2X0 U6988 ( .IN1(n7039), .IN2(n7040), .QN(n7003) );
  MUX21X1 U6989 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1509 ), .Q(n7040) );
  MUX21X1 U6990 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1510 ), .Q(n7039) );
  XOR2X1 U6991 ( .IN1(n6930), .IN2(n6929), .Q(n6967) );
  NAND2X0 U6992 ( .IN1(n7041), .IN2(n7042), .QN(n6929) );
  MUX21X1 U6993 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1504 ), .Q(n7042) );
  MUX21X1 U6994 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1503 ), .Q(n7041) );
  NAND2X0 U6995 ( .IN1(n7043), .IN2(n7044), .QN(n6930) );
  MUX21X1 U6996 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1506 ), .Q(n7044) );
  MUX21X1 U6997 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1505 ), .Q(n7043) );
  XOR2X1 U6998 ( .IN1(n6968), .IN2(n7045), .Q(n7024) );
  NAND2X0 U6999 ( .IN1(n6971), .IN2(n6972), .QN(n7045) );
  AO22X1 U7000 ( .IN1(n7046), .IN2(n7047), .IN3(n7048), .IN4(n7049), .Q(n6968)
         );
  OR2X1 U7001 ( .IN1(n7047), .IN2(n7046), .Q(n7048) );
  AO22X1 U7002 ( .IN1(n7050), .IN2(n7051), .IN3(n7052), .IN4(n6148), .Q(
        \i_m4stg_frac/a0cout[50] ) );
  AO22X1 U7003 ( .IN1(n7053), .IN2(n7054), .IN3(n7055), .IN4(n7056), .Q(n6148)
         );
  OR2X1 U7004 ( .IN1(n7053), .IN2(n7054), .Q(n7056) );
  AND2X1 U7005 ( .IN1(n7057), .IN2(n7058), .Q(n7055) );
  NAND2X0 U7006 ( .IN1(n6149), .IN2(n6147), .QN(n7052) );
  INVX0 U7007 ( .INP(n7050), .ZN(n6147) );
  INVX0 U7008 ( .INP(n6149), .ZN(n7051) );
  MUX21X1 U7009 ( .IN1(n7059), .IN2(n7060), .S(n7061), .Q(n6149) );
  INVX0 U7010 ( .INP(n7062), .ZN(n7061) );
  XOR2X1 U7011 ( .IN1(n7019), .IN2(n7017), .Q(n7050) );
  OA22X1 U7012 ( .IN1(n7063), .IN2(n7064), .IN3(n7065), .IN4(n7066), .Q(n7017)
         );
  AND2X1 U7013 ( .IN1(n7064), .IN2(n7063), .Q(n7066) );
  XNOR3X1 U7014 ( .IN1(n7067), .IN2(n7010), .IN3(n7016), .Q(n7019) );
  XOR3X1 U7015 ( .IN1(n7022), .IN2(n7021), .IN3(n7020), .Q(n7016) );
  XNOR3X1 U7016 ( .IN1(n7031), .IN2(n7032), .IN3(n7034), .Q(n7020) );
  NAND2X0 U7017 ( .IN1(n7068), .IN2(n7069), .QN(n7034) );
  MUX21X1 U7018 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1512 ), .Q(n7069) );
  MUX21X1 U7019 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1513 ), .Q(n7068) );
  NAND2X0 U7020 ( .IN1(n7070), .IN2(n7071), .QN(n7032) );
  MUX21X1 U7021 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1517 ), .Q(n7071) );
  MUX21X1 U7022 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1516 ), .Q(n7070) );
  NAND2X0 U7023 ( .IN1(n7072), .IN2(n7073), .QN(n7031) );
  MUX21X1 U7024 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1515 ), .Q(n7073) );
  MUX21X1 U7025 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1514 ), .Q(n7072) );
  AOI22X1 U7026 ( .IN1(n7074), .IN2(n7075), .IN3(n7076), .IN4(n7077), .QN(
        n7021) );
  OR2X1 U7027 ( .IN1(n7075), .IN2(n7074), .Q(n7076) );
  XNOR3X1 U7028 ( .IN1(n7046), .IN2(n7047), .IN3(n7049), .Q(n7022) );
  NAND2X0 U7029 ( .IN1(n7078), .IN2(n7079), .QN(n7049) );
  MUX21X1 U7030 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1506 ), .Q(n7079) );
  MUX21X1 U7031 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1507 ), .Q(n7078) );
  NAND2X0 U7032 ( .IN1(n7080), .IN2(n7081), .QN(n7047) );
  MUX21X1 U7033 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1511 ), .Q(n7081) );
  MUX21X1 U7034 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1510 ), .Q(n7080) );
  NAND2X0 U7035 ( .IN1(n7082), .IN2(n7083), .QN(n7046) );
  MUX21X1 U7036 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1508 ), .Q(n7083) );
  MUX21X1 U7037 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1509 ), .Q(n7082) );
  XOR2X1 U7038 ( .IN1(n6972), .IN2(n6971), .Q(n7010) );
  NAND2X0 U7039 ( .IN1(n7084), .IN2(n7085), .QN(n6971) );
  MUX21X1 U7040 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1503 ), .Q(n7085) );
  MUX21X1 U7041 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1502 ), .Q(n7084) );
  NAND2X0 U7042 ( .IN1(n7086), .IN2(n7087), .QN(n6972) );
  MUX21X1 U7043 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1505 ), .Q(n7087) );
  MUX21X1 U7044 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1504 ), .Q(n7086) );
  XOR2X1 U7045 ( .IN1(n7011), .IN2(n7088), .Q(n7067) );
  NAND2X0 U7046 ( .IN1(n7014), .IN2(n7015), .QN(n7088) );
  AO22X1 U7047 ( .IN1(n7089), .IN2(n7090), .IN3(n7091), .IN4(n7092), .Q(n7011)
         );
  OR2X1 U7048 ( .IN1(n7090), .IN2(n7089), .Q(n7091) );
  NOR2X0 U7049 ( .IN1(n6150), .IN2(n6151), .QN(\i_m4stg_frac/a0cout[4] ) );
  XNOR3X1 U7050 ( .IN1(n6694), .IN2(n6695), .IN3(n6696), .Q(n6151) );
  XOR3X1 U7051 ( .IN1(n6690), .IN2(n6691), .IN3(n6693), .Q(n6696) );
  NAND2X0 U7052 ( .IN1(n7093), .IN2(n7094), .QN(n6693) );
  MUX21X1 U7053 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1468 ), .Q(n7094) );
  MUX21X1 U7054 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1469 ), .Q(n7093) );
  NAND2X0 U7055 ( .IN1(n7095), .IN2(n7096), .QN(n6691) );
  MUX21X1 U7056 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1471 ), .Q(n7096) );
  MUX21X1 U7057 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1470 ), .Q(n7095) );
  INVX0 U7058 ( .INP(n7097), .ZN(n6690) );
  MUX21X1 U7059 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1467 ), .Q(n7097) );
  AO22X1 U7060 ( .IN1(n7098), .IN2(n7099), .IN3(n7100), .IN4(n7101), .Q(n6695)
         );
  OR2X1 U7061 ( .IN1(n7099), .IN2(n7098), .Q(n7101) );
  AOI22X1 U7062 ( .IN1(n7102), .IN2(n7103), .IN3(n7104), .IN4(n6182), .QN(
        n6150) );
  NAND2X0 U7063 ( .IN1(n7105), .IN2(n7106), .QN(n6182) );
  NAND3X0 U7064 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(n7107), .IN3(n7108), .QN(
        n7106) );
  INVX0 U7065 ( .INP(n6337), .ZN(n7108) );
  OAI21X1 U7066 ( .IN1(n7107), .IN2(n1034), .IN3(n7109), .QN(n7105) );
  NAND2X0 U7067 ( .IN1(n6184), .IN2(n6183), .QN(n7104) );
  INVX0 U7068 ( .INP(n6184), .ZN(n7103) );
  XOR3X1 U7069 ( .IN1(n6338), .IN2(n7099), .IN3(n7098), .Q(n6184) );
  NAND2X0 U7070 ( .IN1(n7110), .IN2(n7111), .QN(n7098) );
  MUX21X1 U7071 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1470 ), .Q(n7111) );
  MUX21X1 U7072 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1469 ), .Q(n7110) );
  NAND2X0 U7073 ( .IN1(n7112), .IN2(n7113), .QN(n7099) );
  MUX21X1 U7074 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1468 ), .Q(n7113) );
  MUX21X1 U7075 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1467 ), .Q(n7112) );
  INVX0 U7076 ( .INP(n6183), .ZN(n7102) );
  NAND2X0 U7077 ( .IN1(n6215), .IN2(n6216), .QN(n6183) );
  XNOR2X1 U7078 ( .IN1(n7114), .IN2(n7107), .Q(n6216) );
  NAND2X0 U7079 ( .IN1(n7115), .IN2(n7116), .QN(n7107) );
  MUX21X1 U7080 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1468 ), .Q(n7116) );
  MUX21X1 U7081 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1469 ), .Q(n7115) );
  NAND3X0 U7082 ( .IN1(\i_m4stg_frac/n1467 ), .IN2(n933), .IN3(
        \i_m4stg_frac/n1018 ), .QN(n7114) );
  AND3X1 U7083 ( .IN1(n6249), .IN2(n1034), .IN3(n6248), .Q(n6215) );
  NOR2X0 U7084 ( .IN1(\i_m4stg_frac/n1020 ), .IN2(\i_m4stg_frac/n1019 ), .QN(
        n6248) );
  NAND3X0 U7085 ( .IN1(n7117), .IN2(n6332), .IN3(n7118), .QN(n6249) );
  MUX21X1 U7086 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1468 ), .Q(n7118) );
  OR2X1 U7087 ( .IN1(n6333), .IN2(n1034), .Q(n7117) );
  AO22X1 U7088 ( .IN1(n7119), .IN2(n7120), .IN3(n7121), .IN4(n6153), .Q(
        \i_m4stg_frac/a0cout[49] ) );
  AO22X1 U7089 ( .IN1(n7122), .IN2(n7123), .IN3(n7124), .IN4(n7125), .Q(n6153)
         );
  OR2X1 U7090 ( .IN1(n7122), .IN2(n7123), .Q(n7125) );
  AND2X1 U7091 ( .IN1(n7126), .IN2(n7127), .Q(n7124) );
  NAND2X0 U7092 ( .IN1(n6154), .IN2(n6152), .QN(n7121) );
  INVX0 U7093 ( .INP(n7119), .ZN(n6152) );
  INVX0 U7094 ( .INP(n6154), .ZN(n7120) );
  MUX21X1 U7095 ( .IN1(n7128), .IN2(n7129), .S(n7130), .Q(n6154) );
  INVX0 U7096 ( .INP(n7131), .ZN(n7130) );
  XOR2X1 U7097 ( .IN1(n7062), .IN2(n7060), .Q(n7119) );
  OA22X1 U7098 ( .IN1(n7132), .IN2(n7133), .IN3(n7134), .IN4(n7135), .Q(n7060)
         );
  AND2X1 U7099 ( .IN1(n7133), .IN2(n7132), .Q(n7135) );
  XNOR3X1 U7100 ( .IN1(n7136), .IN2(n7053), .IN3(n7059), .Q(n7062) );
  XOR3X1 U7101 ( .IN1(n7065), .IN2(n7064), .IN3(n7063), .Q(n7059) );
  XNOR3X1 U7102 ( .IN1(n7074), .IN2(n7075), .IN3(n7077), .Q(n7063) );
  NAND2X0 U7103 ( .IN1(n7137), .IN2(n7138), .QN(n7077) );
  MUX21X1 U7104 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1511 ), .Q(n7138) );
  MUX21X1 U7105 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1512 ), .Q(n7137) );
  NAND2X0 U7106 ( .IN1(n7139), .IN2(n7140), .QN(n7075) );
  MUX21X1 U7107 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1516 ), .Q(n7140) );
  MUX21X1 U7108 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1515 ), .Q(n7139) );
  NAND2X0 U7109 ( .IN1(n7141), .IN2(n7142), .QN(n7074) );
  MUX21X1 U7110 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1514 ), .Q(n7142) );
  MUX21X1 U7111 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1513 ), .Q(n7141) );
  AOI22X1 U7112 ( .IN1(n7143), .IN2(n7144), .IN3(n7145), .IN4(n7146), .QN(
        n7064) );
  OR2X1 U7113 ( .IN1(n7144), .IN2(n7143), .Q(n7145) );
  XNOR3X1 U7114 ( .IN1(n7089), .IN2(n7090), .IN3(n7092), .Q(n7065) );
  NAND2X0 U7115 ( .IN1(n7147), .IN2(n7148), .QN(n7092) );
  MUX21X1 U7116 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1505 ), .Q(n7148) );
  MUX21X1 U7117 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1506 ), .Q(n7147) );
  NAND2X0 U7118 ( .IN1(n7149), .IN2(n7150), .QN(n7090) );
  MUX21X1 U7119 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1510 ), .Q(n7150) );
  MUX21X1 U7120 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1509 ), .Q(n7149) );
  NAND2X0 U7121 ( .IN1(n7151), .IN2(n7152), .QN(n7089) );
  MUX21X1 U7122 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1507 ), .Q(n7152) );
  MUX21X1 U7123 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1508 ), .Q(n7151) );
  XOR2X1 U7124 ( .IN1(n7015), .IN2(n7014), .Q(n7053) );
  NAND2X0 U7125 ( .IN1(n7153), .IN2(n7154), .QN(n7014) );
  MUX21X1 U7126 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1502 ), .Q(n7154) );
  MUX21X1 U7127 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1501 ), .Q(n7153) );
  NAND2X0 U7128 ( .IN1(n7155), .IN2(n7156), .QN(n7015) );
  MUX21X1 U7129 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1504 ), .Q(n7156) );
  MUX21X1 U7130 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1503 ), .Q(n7155) );
  XOR2X1 U7131 ( .IN1(n7054), .IN2(n7157), .Q(n7136) );
  NAND2X0 U7132 ( .IN1(n7057), .IN2(n7058), .QN(n7157) );
  AO22X1 U7133 ( .IN1(n7158), .IN2(n7159), .IN3(n7160), .IN4(n7161), .Q(n7054)
         );
  OR2X1 U7134 ( .IN1(n7159), .IN2(n7158), .Q(n7160) );
  AO22X1 U7135 ( .IN1(n7162), .IN2(n7163), .IN3(n7164), .IN4(n6156), .Q(
        \i_m4stg_frac/a0cout[48] ) );
  AO22X1 U7136 ( .IN1(n7165), .IN2(n7166), .IN3(n7167), .IN4(n7168), .Q(n6156)
         );
  OR2X1 U7137 ( .IN1(n7165), .IN2(n7166), .Q(n7168) );
  AND2X1 U7138 ( .IN1(n7169), .IN2(n7170), .Q(n7167) );
  NAND2X0 U7139 ( .IN1(n6157), .IN2(n6155), .QN(n7164) );
  INVX0 U7140 ( .INP(n7162), .ZN(n6155) );
  INVX0 U7141 ( .INP(n6157), .ZN(n7163) );
  MUX21X1 U7142 ( .IN1(n7171), .IN2(n7172), .S(n7173), .Q(n6157) );
  INVX0 U7143 ( .INP(n7174), .ZN(n7173) );
  XOR2X1 U7144 ( .IN1(n7131), .IN2(n7129), .Q(n7162) );
  OA22X1 U7145 ( .IN1(n7175), .IN2(n7176), .IN3(n7177), .IN4(n7178), .Q(n7129)
         );
  AND2X1 U7146 ( .IN1(n7176), .IN2(n7175), .Q(n7178) );
  XNOR3X1 U7147 ( .IN1(n7179), .IN2(n7122), .IN3(n7128), .Q(n7131) );
  XOR3X1 U7148 ( .IN1(n7134), .IN2(n7133), .IN3(n7132), .Q(n7128) );
  XNOR3X1 U7149 ( .IN1(n7143), .IN2(n7144), .IN3(n7146), .Q(n7132) );
  NAND2X0 U7150 ( .IN1(n7180), .IN2(n7181), .QN(n7146) );
  MUX21X1 U7151 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1510 ), .Q(n7181) );
  MUX21X1 U7152 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1511 ), .Q(n7180) );
  NAND2X0 U7153 ( .IN1(n7182), .IN2(n7183), .QN(n7144) );
  MUX21X1 U7154 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1515 ), .Q(n7183) );
  MUX21X1 U7155 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1514 ), .Q(n7182) );
  NAND2X0 U7156 ( .IN1(n7184), .IN2(n7185), .QN(n7143) );
  MUX21X1 U7157 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1513 ), .Q(n7185) );
  MUX21X1 U7158 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1512 ), .Q(n7184) );
  AOI22X1 U7159 ( .IN1(n7186), .IN2(n7187), .IN3(n7188), .IN4(n7189), .QN(
        n7133) );
  OR2X1 U7160 ( .IN1(n7187), .IN2(n7186), .Q(n7188) );
  XNOR3X1 U7161 ( .IN1(n7158), .IN2(n7159), .IN3(n7161), .Q(n7134) );
  NAND2X0 U7162 ( .IN1(n7190), .IN2(n7191), .QN(n7161) );
  MUX21X1 U7163 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1504 ), .Q(n7191) );
  MUX21X1 U7164 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1505 ), .Q(n7190) );
  NAND2X0 U7165 ( .IN1(n7192), .IN2(n7193), .QN(n7159) );
  MUX21X1 U7166 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1509 ), .Q(n7193) );
  MUX21X1 U7167 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1508 ), .Q(n7192) );
  NAND2X0 U7168 ( .IN1(n7194), .IN2(n7195), .QN(n7158) );
  MUX21X1 U7169 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1506 ), .Q(n7195) );
  MUX21X1 U7170 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1507 ), .Q(n7194) );
  XOR2X1 U7171 ( .IN1(n7058), .IN2(n7057), .Q(n7122) );
  NAND2X0 U7172 ( .IN1(n7196), .IN2(n7197), .QN(n7057) );
  MUX21X1 U7173 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1501 ), .Q(n7197) );
  MUX21X1 U7174 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1500 ), .Q(n7196) );
  NAND2X0 U7175 ( .IN1(n7198), .IN2(n7199), .QN(n7058) );
  MUX21X1 U7176 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1503 ), .Q(n7199) );
  MUX21X1 U7177 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1502 ), .Q(n7198) );
  XOR2X1 U7178 ( .IN1(n7123), .IN2(n7200), .Q(n7179) );
  NAND2X0 U7179 ( .IN1(n7126), .IN2(n7127), .QN(n7200) );
  AO22X1 U7180 ( .IN1(n7201), .IN2(n7202), .IN3(n7203), .IN4(n7204), .Q(n7123)
         );
  OR2X1 U7181 ( .IN1(n7202), .IN2(n7201), .Q(n7203) );
  AO22X1 U7182 ( .IN1(n7205), .IN2(n7206), .IN3(n7207), .IN4(n6159), .Q(
        \i_m4stg_frac/a0cout[47] ) );
  AO22X1 U7183 ( .IN1(n7208), .IN2(n7209), .IN3(n7210), .IN4(n7211), .Q(n6159)
         );
  OR2X1 U7184 ( .IN1(n7208), .IN2(n7209), .Q(n7211) );
  AND2X1 U7185 ( .IN1(n7212), .IN2(n7213), .Q(n7210) );
  NAND2X0 U7186 ( .IN1(n6160), .IN2(n6158), .QN(n7207) );
  INVX0 U7187 ( .INP(n7205), .ZN(n6158) );
  INVX0 U7188 ( .INP(n6160), .ZN(n7206) );
  MUX21X1 U7189 ( .IN1(n7214), .IN2(n7215), .S(n7216), .Q(n6160) );
  INVX0 U7190 ( .INP(n7217), .ZN(n7216) );
  XOR2X1 U7191 ( .IN1(n7174), .IN2(n7172), .Q(n7205) );
  OA22X1 U7192 ( .IN1(n7218), .IN2(n7219), .IN3(n7220), .IN4(n7221), .Q(n7172)
         );
  AND2X1 U7193 ( .IN1(n7219), .IN2(n7218), .Q(n7221) );
  XNOR3X1 U7194 ( .IN1(n7222), .IN2(n7165), .IN3(n7171), .Q(n7174) );
  XOR3X1 U7195 ( .IN1(n7177), .IN2(n7176), .IN3(n7175), .Q(n7171) );
  XNOR3X1 U7196 ( .IN1(n7186), .IN2(n7187), .IN3(n7189), .Q(n7175) );
  NAND2X0 U7197 ( .IN1(n7223), .IN2(n7224), .QN(n7189) );
  MUX21X1 U7198 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1509 ), .Q(n7224) );
  MUX21X1 U7199 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1510 ), .Q(n7223) );
  NAND2X0 U7200 ( .IN1(n7225), .IN2(n7226), .QN(n7187) );
  MUX21X1 U7201 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1514 ), .Q(n7226) );
  MUX21X1 U7202 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1513 ), .Q(n7225) );
  NAND2X0 U7203 ( .IN1(n7227), .IN2(n7228), .QN(n7186) );
  MUX21X1 U7204 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1512 ), .Q(n7228) );
  MUX21X1 U7205 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1511 ), .Q(n7227) );
  AOI22X1 U7206 ( .IN1(n7229), .IN2(n7230), .IN3(n7231), .IN4(n7232), .QN(
        n7176) );
  OR2X1 U7207 ( .IN1(n7230), .IN2(n7229), .Q(n7231) );
  XNOR3X1 U7208 ( .IN1(n7201), .IN2(n7202), .IN3(n7204), .Q(n7177) );
  NAND2X0 U7209 ( .IN1(n7233), .IN2(n7234), .QN(n7204) );
  MUX21X1 U7210 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1503 ), .Q(n7234) );
  MUX21X1 U7211 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1504 ), .Q(n7233) );
  NAND2X0 U7212 ( .IN1(n7235), .IN2(n7236), .QN(n7202) );
  MUX21X1 U7213 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1508 ), .Q(n7236) );
  MUX21X1 U7214 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1507 ), .Q(n7235) );
  NAND2X0 U7215 ( .IN1(n7237), .IN2(n7238), .QN(n7201) );
  MUX21X1 U7216 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1505 ), .Q(n7238) );
  MUX21X1 U7217 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1506 ), .Q(n7237) );
  XOR2X1 U7218 ( .IN1(n7127), .IN2(n7126), .Q(n7165) );
  NAND2X0 U7219 ( .IN1(n7239), .IN2(n7240), .QN(n7126) );
  MUX21X1 U7220 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1500 ), .Q(n7240) );
  MUX21X1 U7221 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1499 ), .Q(n7239) );
  NAND2X0 U7222 ( .IN1(n7241), .IN2(n7242), .QN(n7127) );
  MUX21X1 U7223 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1502 ), .Q(n7242) );
  MUX21X1 U7224 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1501 ), .Q(n7241) );
  XOR2X1 U7225 ( .IN1(n7166), .IN2(n7243), .Q(n7222) );
  NAND2X0 U7226 ( .IN1(n7169), .IN2(n7170), .QN(n7243) );
  AO22X1 U7227 ( .IN1(n7244), .IN2(n7245), .IN3(n7246), .IN4(n7247), .Q(n7166)
         );
  OR2X1 U7228 ( .IN1(n7245), .IN2(n7244), .Q(n7246) );
  AO22X1 U7229 ( .IN1(n7248), .IN2(n7249), .IN3(n7250), .IN4(n6162), .Q(
        \i_m4stg_frac/a0cout[46] ) );
  AO22X1 U7230 ( .IN1(n7251), .IN2(n7252), .IN3(n7253), .IN4(n7254), .Q(n6162)
         );
  OR2X1 U7231 ( .IN1(n7251), .IN2(n7252), .Q(n7254) );
  AND2X1 U7232 ( .IN1(n7255), .IN2(n7256), .Q(n7253) );
  NAND2X0 U7233 ( .IN1(n6163), .IN2(n6161), .QN(n7250) );
  INVX0 U7234 ( .INP(n7248), .ZN(n6161) );
  INVX0 U7235 ( .INP(n6163), .ZN(n7249) );
  MUX21X1 U7236 ( .IN1(n7257), .IN2(n7258), .S(n7259), .Q(n6163) );
  INVX0 U7237 ( .INP(n7260), .ZN(n7259) );
  XOR2X1 U7238 ( .IN1(n7217), .IN2(n7215), .Q(n7248) );
  OA22X1 U7239 ( .IN1(n7261), .IN2(n7262), .IN3(n7263), .IN4(n7264), .Q(n7215)
         );
  AND2X1 U7240 ( .IN1(n7262), .IN2(n7261), .Q(n7264) );
  XNOR3X1 U7241 ( .IN1(n7265), .IN2(n7208), .IN3(n7214), .Q(n7217) );
  XOR3X1 U7242 ( .IN1(n7220), .IN2(n7219), .IN3(n7218), .Q(n7214) );
  XNOR3X1 U7243 ( .IN1(n7229), .IN2(n7230), .IN3(n7232), .Q(n7218) );
  NAND2X0 U7244 ( .IN1(n7266), .IN2(n7267), .QN(n7232) );
  MUX21X1 U7245 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1508 ), .Q(n7267) );
  MUX21X1 U7246 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1509 ), .Q(n7266) );
  NAND2X0 U7247 ( .IN1(n7268), .IN2(n7269), .QN(n7230) );
  MUX21X1 U7248 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1513 ), .Q(n7269) );
  MUX21X1 U7249 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1512 ), .Q(n7268) );
  NAND2X0 U7250 ( .IN1(n7270), .IN2(n7271), .QN(n7229) );
  MUX21X1 U7251 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1511 ), .Q(n7271) );
  MUX21X1 U7252 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1510 ), .Q(n7270) );
  AOI22X1 U7253 ( .IN1(n7272), .IN2(n7273), .IN3(n7274), .IN4(n7275), .QN(
        n7219) );
  OR2X1 U7254 ( .IN1(n7273), .IN2(n7272), .Q(n7274) );
  XNOR3X1 U7255 ( .IN1(n7244), .IN2(n7245), .IN3(n7247), .Q(n7220) );
  NAND2X0 U7256 ( .IN1(n7276), .IN2(n7277), .QN(n7247) );
  MUX21X1 U7257 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1502 ), .Q(n7277) );
  MUX21X1 U7258 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1503 ), .Q(n7276) );
  NAND2X0 U7259 ( .IN1(n7278), .IN2(n7279), .QN(n7245) );
  MUX21X1 U7260 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1507 ), .Q(n7279) );
  MUX21X1 U7261 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1506 ), .Q(n7278) );
  NAND2X0 U7262 ( .IN1(n7280), .IN2(n7281), .QN(n7244) );
  MUX21X1 U7263 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1504 ), .Q(n7281) );
  MUX21X1 U7264 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1505 ), .Q(n7280) );
  XOR2X1 U7265 ( .IN1(n7170), .IN2(n7169), .Q(n7208) );
  NAND2X0 U7266 ( .IN1(n7282), .IN2(n7283), .QN(n7169) );
  MUX21X1 U7267 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1499 ), .Q(n7283) );
  MUX21X1 U7268 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1498 ), .Q(n7282) );
  NAND2X0 U7269 ( .IN1(n7284), .IN2(n7285), .QN(n7170) );
  MUX21X1 U7270 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1501 ), .Q(n7285) );
  MUX21X1 U7271 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1500 ), .Q(n7284) );
  XOR2X1 U7272 ( .IN1(n7209), .IN2(n7286), .Q(n7265) );
  NAND2X0 U7273 ( .IN1(n7212), .IN2(n7213), .QN(n7286) );
  AO22X1 U7274 ( .IN1(n7287), .IN2(n7288), .IN3(n7289), .IN4(n7290), .Q(n7209)
         );
  OR2X1 U7275 ( .IN1(n7288), .IN2(n7287), .Q(n7289) );
  AO22X1 U7276 ( .IN1(n7291), .IN2(n7292), .IN3(n7293), .IN4(n6165), .Q(
        \i_m4stg_frac/a0cout[45] ) );
  AO22X1 U7277 ( .IN1(n7294), .IN2(n7295), .IN3(n7296), .IN4(n7297), .Q(n6165)
         );
  OR2X1 U7278 ( .IN1(n7294), .IN2(n7295), .Q(n7297) );
  AND2X1 U7279 ( .IN1(n7298), .IN2(n7299), .Q(n7296) );
  NAND2X0 U7280 ( .IN1(n6166), .IN2(n6164), .QN(n7293) );
  INVX0 U7281 ( .INP(n7291), .ZN(n6164) );
  INVX0 U7282 ( .INP(n6166), .ZN(n7292) );
  MUX21X1 U7283 ( .IN1(n7300), .IN2(n7301), .S(n7302), .Q(n6166) );
  INVX0 U7284 ( .INP(n7303), .ZN(n7302) );
  XOR2X1 U7285 ( .IN1(n7260), .IN2(n7258), .Q(n7291) );
  OA22X1 U7286 ( .IN1(n7304), .IN2(n7305), .IN3(n7306), .IN4(n7307), .Q(n7258)
         );
  AND2X1 U7287 ( .IN1(n7305), .IN2(n7304), .Q(n7307) );
  XNOR3X1 U7288 ( .IN1(n7308), .IN2(n7251), .IN3(n7257), .Q(n7260) );
  XOR3X1 U7289 ( .IN1(n7263), .IN2(n7262), .IN3(n7261), .Q(n7257) );
  XNOR3X1 U7290 ( .IN1(n7272), .IN2(n7273), .IN3(n7275), .Q(n7261) );
  NAND2X0 U7291 ( .IN1(n7309), .IN2(n7310), .QN(n7275) );
  MUX21X1 U7292 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1507 ), .Q(n7310) );
  MUX21X1 U7293 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1508 ), .Q(n7309) );
  NAND2X0 U7294 ( .IN1(n7311), .IN2(n7312), .QN(n7273) );
  MUX21X1 U7295 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1512 ), .Q(n7312) );
  MUX21X1 U7296 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1511 ), .Q(n7311) );
  NAND2X0 U7297 ( .IN1(n7313), .IN2(n7314), .QN(n7272) );
  MUX21X1 U7298 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1510 ), .Q(n7314) );
  MUX21X1 U7299 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1509 ), .Q(n7313) );
  AOI22X1 U7300 ( .IN1(n7315), .IN2(n7316), .IN3(n7317), .IN4(n7318), .QN(
        n7262) );
  OR2X1 U7301 ( .IN1(n7316), .IN2(n7315), .Q(n7317) );
  XNOR3X1 U7302 ( .IN1(n7287), .IN2(n7288), .IN3(n7290), .Q(n7263) );
  NAND2X0 U7303 ( .IN1(n7319), .IN2(n7320), .QN(n7290) );
  MUX21X1 U7304 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1501 ), .Q(n7320) );
  MUX21X1 U7305 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1502 ), .Q(n7319) );
  NAND2X0 U7306 ( .IN1(n7321), .IN2(n7322), .QN(n7288) );
  MUX21X1 U7307 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1506 ), .Q(n7322) );
  MUX21X1 U7308 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1505 ), .Q(n7321) );
  NAND2X0 U7309 ( .IN1(n7323), .IN2(n7324), .QN(n7287) );
  MUX21X1 U7310 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1503 ), .Q(n7324) );
  MUX21X1 U7311 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1504 ), .Q(n7323) );
  XOR2X1 U7312 ( .IN1(n7213), .IN2(n7212), .Q(n7251) );
  NAND2X0 U7313 ( .IN1(n7325), .IN2(n7326), .QN(n7212) );
  MUX21X1 U7314 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1498 ), .Q(n7326) );
  MUX21X1 U7315 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1497 ), .Q(n7325) );
  NAND2X0 U7316 ( .IN1(n7327), .IN2(n7328), .QN(n7213) );
  MUX21X1 U7317 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1500 ), .Q(n7328) );
  MUX21X1 U7318 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1499 ), .Q(n7327) );
  XOR2X1 U7319 ( .IN1(n7252), .IN2(n7329), .Q(n7308) );
  NAND2X0 U7320 ( .IN1(n7255), .IN2(n7256), .QN(n7329) );
  AO22X1 U7321 ( .IN1(n7330), .IN2(n7331), .IN3(n7332), .IN4(n7333), .Q(n7252)
         );
  OR2X1 U7322 ( .IN1(n7331), .IN2(n7330), .Q(n7332) );
  AO22X1 U7323 ( .IN1(n7334), .IN2(n7335), .IN3(n7336), .IN4(n6168), .Q(
        \i_m4stg_frac/a0cout[44] ) );
  AO22X1 U7324 ( .IN1(n7337), .IN2(n7338), .IN3(n7339), .IN4(n7340), .Q(n6168)
         );
  OR2X1 U7325 ( .IN1(n7337), .IN2(n7338), .Q(n7340) );
  AND2X1 U7326 ( .IN1(n7341), .IN2(n7342), .Q(n7339) );
  NAND2X0 U7327 ( .IN1(n6169), .IN2(n6167), .QN(n7336) );
  INVX0 U7328 ( .INP(n7334), .ZN(n6167) );
  INVX0 U7329 ( .INP(n6169), .ZN(n7335) );
  MUX21X1 U7330 ( .IN1(n7343), .IN2(n7344), .S(n7345), .Q(n6169) );
  INVX0 U7331 ( .INP(n7346), .ZN(n7345) );
  XOR2X1 U7332 ( .IN1(n7303), .IN2(n7301), .Q(n7334) );
  OA22X1 U7333 ( .IN1(n7347), .IN2(n7348), .IN3(n7349), .IN4(n7350), .Q(n7301)
         );
  AND2X1 U7334 ( .IN1(n7348), .IN2(n7347), .Q(n7350) );
  XNOR3X1 U7335 ( .IN1(n7351), .IN2(n7294), .IN3(n7300), .Q(n7303) );
  XOR3X1 U7336 ( .IN1(n7306), .IN2(n7305), .IN3(n7304), .Q(n7300) );
  XNOR3X1 U7337 ( .IN1(n7315), .IN2(n7316), .IN3(n7318), .Q(n7304) );
  NAND2X0 U7338 ( .IN1(n7352), .IN2(n7353), .QN(n7318) );
  MUX21X1 U7339 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1506 ), .Q(n7353) );
  MUX21X1 U7340 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1507 ), .Q(n7352) );
  NAND2X0 U7341 ( .IN1(n7354), .IN2(n7355), .QN(n7316) );
  MUX21X1 U7342 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1511 ), .Q(n7355) );
  MUX21X1 U7343 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1510 ), .Q(n7354) );
  NAND2X0 U7344 ( .IN1(n7356), .IN2(n7357), .QN(n7315) );
  MUX21X1 U7345 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1509 ), .Q(n7357) );
  MUX21X1 U7346 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1508 ), .Q(n7356) );
  AOI22X1 U7347 ( .IN1(n7358), .IN2(n7359), .IN3(n7360), .IN4(n7361), .QN(
        n7305) );
  OR2X1 U7348 ( .IN1(n7359), .IN2(n7358), .Q(n7360) );
  XNOR3X1 U7349 ( .IN1(n7330), .IN2(n7331), .IN3(n7333), .Q(n7306) );
  NAND2X0 U7350 ( .IN1(n7362), .IN2(n7363), .QN(n7333) );
  MUX21X1 U7351 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1500 ), .Q(n7363) );
  MUX21X1 U7352 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1501 ), .Q(n7362) );
  NAND2X0 U7353 ( .IN1(n7364), .IN2(n7365), .QN(n7331) );
  MUX21X1 U7354 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1505 ), .Q(n7365) );
  MUX21X1 U7355 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1504 ), .Q(n7364) );
  NAND2X0 U7356 ( .IN1(n7366), .IN2(n7367), .QN(n7330) );
  MUX21X1 U7357 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1502 ), .Q(n7367) );
  MUX21X1 U7358 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1503 ), .Q(n7366) );
  XOR2X1 U7359 ( .IN1(n7256), .IN2(n7255), .Q(n7294) );
  NAND2X0 U7360 ( .IN1(n7368), .IN2(n7369), .QN(n7255) );
  MUX21X1 U7361 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1497 ), .Q(n7369) );
  MUX21X1 U7362 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1496 ), .Q(n7368) );
  NAND2X0 U7363 ( .IN1(n7370), .IN2(n7371), .QN(n7256) );
  MUX21X1 U7364 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1499 ), .Q(n7371) );
  MUX21X1 U7365 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1498 ), .Q(n7370) );
  XOR2X1 U7366 ( .IN1(n7295), .IN2(n7372), .Q(n7351) );
  NAND2X0 U7367 ( .IN1(n7298), .IN2(n7299), .QN(n7372) );
  AO22X1 U7368 ( .IN1(n7373), .IN2(n7374), .IN3(n7375), .IN4(n7376), .Q(n7295)
         );
  OR2X1 U7369 ( .IN1(n7374), .IN2(n7373), .Q(n7375) );
  AO22X1 U7370 ( .IN1(n7377), .IN2(n7378), .IN3(n7379), .IN4(n6171), .Q(
        \i_m4stg_frac/a0cout[43] ) );
  AO22X1 U7371 ( .IN1(n7380), .IN2(n7381), .IN3(n7382), .IN4(n7383), .Q(n6171)
         );
  OR2X1 U7372 ( .IN1(n7380), .IN2(n7381), .Q(n7383) );
  AND2X1 U7373 ( .IN1(n7384), .IN2(n7385), .Q(n7382) );
  NAND2X0 U7374 ( .IN1(n6172), .IN2(n6170), .QN(n7379) );
  INVX0 U7375 ( .INP(n7377), .ZN(n6170) );
  INVX0 U7376 ( .INP(n6172), .ZN(n7378) );
  MUX21X1 U7377 ( .IN1(n7386), .IN2(n7387), .S(n7388), .Q(n6172) );
  INVX0 U7378 ( .INP(n7389), .ZN(n7388) );
  XOR2X1 U7379 ( .IN1(n7346), .IN2(n7344), .Q(n7377) );
  OA22X1 U7380 ( .IN1(n7390), .IN2(n7391), .IN3(n7392), .IN4(n7393), .Q(n7344)
         );
  AND2X1 U7381 ( .IN1(n7391), .IN2(n7390), .Q(n7393) );
  XNOR3X1 U7382 ( .IN1(n7394), .IN2(n7337), .IN3(n7343), .Q(n7346) );
  XOR3X1 U7383 ( .IN1(n7349), .IN2(n7348), .IN3(n7347), .Q(n7343) );
  XNOR3X1 U7384 ( .IN1(n7358), .IN2(n7359), .IN3(n7361), .Q(n7347) );
  NAND2X0 U7385 ( .IN1(n7395), .IN2(n7396), .QN(n7361) );
  MUX21X1 U7386 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1505 ), .Q(n7396) );
  MUX21X1 U7387 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1506 ), .Q(n7395) );
  NAND2X0 U7388 ( .IN1(n7397), .IN2(n7398), .QN(n7359) );
  MUX21X1 U7389 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1510 ), .Q(n7398) );
  MUX21X1 U7390 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1509 ), .Q(n7397) );
  NAND2X0 U7391 ( .IN1(n7399), .IN2(n7400), .QN(n7358) );
  MUX21X1 U7392 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1508 ), .Q(n7400) );
  MUX21X1 U7393 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1507 ), .Q(n7399) );
  AOI22X1 U7394 ( .IN1(n7401), .IN2(n7402), .IN3(n7403), .IN4(n7404), .QN(
        n7348) );
  OR2X1 U7395 ( .IN1(n7402), .IN2(n7401), .Q(n7403) );
  XNOR3X1 U7396 ( .IN1(n7373), .IN2(n7374), .IN3(n7376), .Q(n7349) );
  NAND2X0 U7397 ( .IN1(n7405), .IN2(n7406), .QN(n7376) );
  MUX21X1 U7398 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1499 ), .Q(n7406) );
  MUX21X1 U7399 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1500 ), .Q(n7405) );
  NAND2X0 U7400 ( .IN1(n7407), .IN2(n7408), .QN(n7374) );
  MUX21X1 U7401 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1504 ), .Q(n7408) );
  MUX21X1 U7402 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1503 ), .Q(n7407) );
  NAND2X0 U7403 ( .IN1(n7409), .IN2(n7410), .QN(n7373) );
  MUX21X1 U7404 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1501 ), .Q(n7410) );
  MUX21X1 U7405 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1502 ), .Q(n7409) );
  XOR2X1 U7406 ( .IN1(n7299), .IN2(n7298), .Q(n7337) );
  NAND2X0 U7407 ( .IN1(n7411), .IN2(n7412), .QN(n7298) );
  MUX21X1 U7408 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1496 ), .Q(n7412) );
  MUX21X1 U7409 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1495 ), .Q(n7411) );
  NAND2X0 U7410 ( .IN1(n7413), .IN2(n7414), .QN(n7299) );
  MUX21X1 U7411 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1498 ), .Q(n7414) );
  MUX21X1 U7412 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1497 ), .Q(n7413) );
  XOR2X1 U7413 ( .IN1(n7338), .IN2(n7415), .Q(n7394) );
  NAND2X0 U7414 ( .IN1(n7341), .IN2(n7342), .QN(n7415) );
  AO22X1 U7415 ( .IN1(n7416), .IN2(n7417), .IN3(n7418), .IN4(n7419), .Q(n7338)
         );
  OR2X1 U7416 ( .IN1(n7417), .IN2(n7416), .Q(n7418) );
  AO22X1 U7417 ( .IN1(n7420), .IN2(n7421), .IN3(n7422), .IN4(n6174), .Q(
        \i_m4stg_frac/a0cout[42] ) );
  AO22X1 U7418 ( .IN1(n7423), .IN2(n7424), .IN3(n7425), .IN4(n7426), .Q(n6174)
         );
  OR2X1 U7419 ( .IN1(n7423), .IN2(n7424), .Q(n7426) );
  AND2X1 U7420 ( .IN1(n7427), .IN2(n7428), .Q(n7425) );
  NAND2X0 U7421 ( .IN1(n6175), .IN2(n6173), .QN(n7422) );
  INVX0 U7422 ( .INP(n7420), .ZN(n6173) );
  INVX0 U7423 ( .INP(n6175), .ZN(n7421) );
  MUX21X1 U7424 ( .IN1(n7429), .IN2(n7430), .S(n7431), .Q(n6175) );
  INVX0 U7425 ( .INP(n7432), .ZN(n7431) );
  XOR2X1 U7426 ( .IN1(n7389), .IN2(n7387), .Q(n7420) );
  OA22X1 U7427 ( .IN1(n7433), .IN2(n7434), .IN3(n7435), .IN4(n7436), .Q(n7387)
         );
  AND2X1 U7428 ( .IN1(n7434), .IN2(n7433), .Q(n7436) );
  XNOR3X1 U7429 ( .IN1(n7437), .IN2(n7380), .IN3(n7386), .Q(n7389) );
  XOR3X1 U7430 ( .IN1(n7392), .IN2(n7391), .IN3(n7390), .Q(n7386) );
  XNOR3X1 U7431 ( .IN1(n7401), .IN2(n7402), .IN3(n7404), .Q(n7390) );
  NAND2X0 U7432 ( .IN1(n7438), .IN2(n7439), .QN(n7404) );
  MUX21X1 U7433 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1504 ), .Q(n7439) );
  MUX21X1 U7434 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1505 ), .Q(n7438) );
  NAND2X0 U7435 ( .IN1(n7440), .IN2(n7441), .QN(n7402) );
  MUX21X1 U7436 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1509 ), .Q(n7441) );
  MUX21X1 U7437 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1508 ), .Q(n7440) );
  NAND2X0 U7438 ( .IN1(n7442), .IN2(n7443), .QN(n7401) );
  MUX21X1 U7439 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1507 ), .Q(n7443) );
  MUX21X1 U7440 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1506 ), .Q(n7442) );
  AOI22X1 U7441 ( .IN1(n7444), .IN2(n7445), .IN3(n7446), .IN4(n7447), .QN(
        n7391) );
  OR2X1 U7442 ( .IN1(n7445), .IN2(n7444), .Q(n7446) );
  XNOR3X1 U7443 ( .IN1(n7416), .IN2(n7417), .IN3(n7419), .Q(n7392) );
  NAND2X0 U7444 ( .IN1(n7448), .IN2(n7449), .QN(n7419) );
  MUX21X1 U7445 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1498 ), .Q(n7449) );
  MUX21X1 U7446 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1499 ), .Q(n7448) );
  NAND2X0 U7447 ( .IN1(n7450), .IN2(n7451), .QN(n7417) );
  MUX21X1 U7448 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1503 ), .Q(n7451) );
  MUX21X1 U7449 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1502 ), .Q(n7450) );
  NAND2X0 U7450 ( .IN1(n7452), .IN2(n7453), .QN(n7416) );
  MUX21X1 U7451 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1500 ), .Q(n7453) );
  MUX21X1 U7452 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1501 ), .Q(n7452) );
  XOR2X1 U7453 ( .IN1(n7342), .IN2(n7341), .Q(n7380) );
  NAND2X0 U7454 ( .IN1(n7454), .IN2(n7455), .QN(n7341) );
  MUX21X1 U7455 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1495 ), .Q(n7455) );
  MUX21X1 U7456 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1494 ), .Q(n7454) );
  NAND2X0 U7457 ( .IN1(n7456), .IN2(n7457), .QN(n7342) );
  MUX21X1 U7458 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1497 ), .Q(n7457) );
  MUX21X1 U7459 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1496 ), .Q(n7456) );
  XOR2X1 U7460 ( .IN1(n7381), .IN2(n7458), .Q(n7437) );
  NAND2X0 U7461 ( .IN1(n7384), .IN2(n7385), .QN(n7458) );
  AO22X1 U7462 ( .IN1(n7459), .IN2(n7460), .IN3(n7461), .IN4(n7462), .Q(n7381)
         );
  OR2X1 U7463 ( .IN1(n7460), .IN2(n7459), .Q(n7461) );
  AO22X1 U7464 ( .IN1(n7463), .IN2(n7464), .IN3(n7465), .IN4(n6177), .Q(
        \i_m4stg_frac/a0cout[41] ) );
  AO22X1 U7465 ( .IN1(n7466), .IN2(n7467), .IN3(n7468), .IN4(n7469), .Q(n6177)
         );
  OR2X1 U7466 ( .IN1(n7466), .IN2(n7467), .Q(n7469) );
  AND2X1 U7467 ( .IN1(n7470), .IN2(n7471), .Q(n7468) );
  NAND2X0 U7468 ( .IN1(n6178), .IN2(n6176), .QN(n7465) );
  INVX0 U7469 ( .INP(n7463), .ZN(n6176) );
  INVX0 U7470 ( .INP(n6178), .ZN(n7464) );
  MUX21X1 U7471 ( .IN1(n7472), .IN2(n7473), .S(n7474), .Q(n6178) );
  INVX0 U7472 ( .INP(n7475), .ZN(n7474) );
  XOR2X1 U7473 ( .IN1(n7432), .IN2(n7430), .Q(n7463) );
  OA22X1 U7474 ( .IN1(n7476), .IN2(n7477), .IN3(n7478), .IN4(n7479), .Q(n7430)
         );
  AND2X1 U7475 ( .IN1(n7477), .IN2(n7476), .Q(n7479) );
  XNOR3X1 U7476 ( .IN1(n7480), .IN2(n7423), .IN3(n7429), .Q(n7432) );
  XOR3X1 U7477 ( .IN1(n7435), .IN2(n7434), .IN3(n7433), .Q(n7429) );
  XNOR3X1 U7478 ( .IN1(n7444), .IN2(n7445), .IN3(n7447), .Q(n7433) );
  NAND2X0 U7479 ( .IN1(n7481), .IN2(n7482), .QN(n7447) );
  MUX21X1 U7480 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1503 ), .Q(n7482) );
  MUX21X1 U7481 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1504 ), .Q(n7481) );
  NAND2X0 U7482 ( .IN1(n7483), .IN2(n7484), .QN(n7445) );
  MUX21X1 U7483 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1508 ), .Q(n7484) );
  MUX21X1 U7484 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1507 ), .Q(n7483) );
  NAND2X0 U7485 ( .IN1(n7485), .IN2(n7486), .QN(n7444) );
  MUX21X1 U7486 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1506 ), .Q(n7486) );
  MUX21X1 U7487 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1505 ), .Q(n7485) );
  AOI22X1 U7488 ( .IN1(n7487), .IN2(n7488), .IN3(n7489), .IN4(n7490), .QN(
        n7434) );
  OR2X1 U7489 ( .IN1(n7488), .IN2(n7487), .Q(n7489) );
  XNOR3X1 U7490 ( .IN1(n7459), .IN2(n7460), .IN3(n7462), .Q(n7435) );
  NAND2X0 U7491 ( .IN1(n7491), .IN2(n7492), .QN(n7462) );
  MUX21X1 U7492 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1497 ), .Q(n7492) );
  MUX21X1 U7493 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1498 ), .Q(n7491) );
  NAND2X0 U7494 ( .IN1(n7493), .IN2(n7494), .QN(n7460) );
  MUX21X1 U7495 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1502 ), .Q(n7494) );
  MUX21X1 U7496 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1501 ), .Q(n7493) );
  NAND2X0 U7497 ( .IN1(n7495), .IN2(n7496), .QN(n7459) );
  MUX21X1 U7498 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1499 ), .Q(n7496) );
  MUX21X1 U7499 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1500 ), .Q(n7495) );
  XOR2X1 U7500 ( .IN1(n7385), .IN2(n7384), .Q(n7423) );
  NAND2X0 U7501 ( .IN1(n7497), .IN2(n7498), .QN(n7384) );
  MUX21X1 U7502 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1494 ), .Q(n7498) );
  MUX21X1 U7503 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1493 ), .Q(n7497) );
  NAND2X0 U7504 ( .IN1(n7499), .IN2(n7500), .QN(n7385) );
  MUX21X1 U7505 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1496 ), .Q(n7500) );
  MUX21X1 U7506 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1495 ), .Q(n7499) );
  XOR2X1 U7507 ( .IN1(n7424), .IN2(n7501), .Q(n7480) );
  NAND2X0 U7508 ( .IN1(n7427), .IN2(n7428), .QN(n7501) );
  AO22X1 U7509 ( .IN1(n7502), .IN2(n7503), .IN3(n7504), .IN4(n7505), .Q(n7424)
         );
  OR2X1 U7510 ( .IN1(n7503), .IN2(n7502), .Q(n7504) );
  AO22X1 U7511 ( .IN1(n7506), .IN2(n7507), .IN3(n7508), .IN4(n6180), .Q(
        \i_m4stg_frac/a0cout[40] ) );
  AO22X1 U7512 ( .IN1(n7509), .IN2(n7510), .IN3(n7511), .IN4(n7512), .Q(n6180)
         );
  OR2X1 U7513 ( .IN1(n7509), .IN2(n7510), .Q(n7512) );
  AND2X1 U7514 ( .IN1(n7513), .IN2(n7514), .Q(n7511) );
  NAND2X0 U7515 ( .IN1(n6181), .IN2(n6179), .QN(n7508) );
  INVX0 U7516 ( .INP(n7506), .ZN(n6179) );
  INVX0 U7517 ( .INP(n6181), .ZN(n7507) );
  MUX21X1 U7518 ( .IN1(n7515), .IN2(n7516), .S(n7517), .Q(n6181) );
  INVX0 U7519 ( .INP(n7518), .ZN(n7517) );
  XOR2X1 U7520 ( .IN1(n7475), .IN2(n7473), .Q(n7506) );
  OA22X1 U7521 ( .IN1(n7519), .IN2(n7520), .IN3(n7521), .IN4(n7522), .Q(n7473)
         );
  AND2X1 U7522 ( .IN1(n7520), .IN2(n7519), .Q(n7522) );
  XNOR3X1 U7523 ( .IN1(n7523), .IN2(n7466), .IN3(n7472), .Q(n7475) );
  XOR3X1 U7524 ( .IN1(n7478), .IN2(n7477), .IN3(n7476), .Q(n7472) );
  XNOR3X1 U7525 ( .IN1(n7487), .IN2(n7488), .IN3(n7490), .Q(n7476) );
  NAND2X0 U7526 ( .IN1(n7524), .IN2(n7525), .QN(n7490) );
  MUX21X1 U7527 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1502 ), .Q(n7525) );
  MUX21X1 U7528 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1503 ), .Q(n7524) );
  NAND2X0 U7529 ( .IN1(n7526), .IN2(n7527), .QN(n7488) );
  MUX21X1 U7530 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1507 ), .Q(n7527) );
  MUX21X1 U7531 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1506 ), .Q(n7526) );
  NAND2X0 U7532 ( .IN1(n7528), .IN2(n7529), .QN(n7487) );
  MUX21X1 U7533 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1505 ), .Q(n7529) );
  MUX21X1 U7534 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1504 ), .Q(n7528) );
  AOI22X1 U7535 ( .IN1(n7530), .IN2(n7531), .IN3(n7532), .IN4(n7533), .QN(
        n7477) );
  OR2X1 U7536 ( .IN1(n7531), .IN2(n7530), .Q(n7532) );
  XNOR3X1 U7537 ( .IN1(n7502), .IN2(n7503), .IN3(n7505), .Q(n7478) );
  NAND2X0 U7538 ( .IN1(n7534), .IN2(n7535), .QN(n7505) );
  MUX21X1 U7539 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1496 ), .Q(n7535) );
  MUX21X1 U7540 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1497 ), .Q(n7534) );
  NAND2X0 U7541 ( .IN1(n7536), .IN2(n7537), .QN(n7503) );
  MUX21X1 U7542 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1501 ), .Q(n7537) );
  MUX21X1 U7543 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1500 ), .Q(n7536) );
  NAND2X0 U7544 ( .IN1(n7538), .IN2(n7539), .QN(n7502) );
  MUX21X1 U7545 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1498 ), .Q(n7539) );
  MUX21X1 U7546 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1499 ), .Q(n7538) );
  XOR2X1 U7547 ( .IN1(n7428), .IN2(n7427), .Q(n7466) );
  NAND2X0 U7548 ( .IN1(n7540), .IN2(n7541), .QN(n7427) );
  MUX21X1 U7549 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1493 ), .Q(n7541) );
  MUX21X1 U7550 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1492 ), .Q(n7540) );
  NAND2X0 U7551 ( .IN1(n7542), .IN2(n7543), .QN(n7428) );
  MUX21X1 U7552 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1495 ), .Q(n7543) );
  MUX21X1 U7553 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1494 ), .Q(n7542) );
  XOR2X1 U7554 ( .IN1(n7467), .IN2(n7544), .Q(n7523) );
  NAND2X0 U7555 ( .IN1(n7470), .IN2(n7471), .QN(n7544) );
  AO22X1 U7556 ( .IN1(n7545), .IN2(n7546), .IN3(n7547), .IN4(n7548), .Q(n7467)
         );
  OR2X1 U7557 ( .IN1(n7546), .IN2(n7545), .Q(n7547) );
  AO22X1 U7558 ( .IN1(n7549), .IN2(n7550), .IN3(n7551), .IN4(n6186), .Q(
        \i_m4stg_frac/a0cout[39] ) );
  AO22X1 U7559 ( .IN1(n7552), .IN2(n7553), .IN3(n7554), .IN4(n7555), .Q(n6186)
         );
  OR2X1 U7560 ( .IN1(n7552), .IN2(n7553), .Q(n7555) );
  AND2X1 U7561 ( .IN1(n7556), .IN2(n7557), .Q(n7554) );
  NAND2X0 U7562 ( .IN1(n6187), .IN2(n6185), .QN(n7551) );
  INVX0 U7563 ( .INP(n7549), .ZN(n6185) );
  INVX0 U7564 ( .INP(n6187), .ZN(n7550) );
  MUX21X1 U7565 ( .IN1(n7558), .IN2(n7559), .S(n7560), .Q(n6187) );
  INVX0 U7566 ( .INP(n7561), .ZN(n7560) );
  XOR2X1 U7567 ( .IN1(n7518), .IN2(n7516), .Q(n7549) );
  OA22X1 U7568 ( .IN1(n7562), .IN2(n7563), .IN3(n7564), .IN4(n7565), .Q(n7516)
         );
  AND2X1 U7569 ( .IN1(n7563), .IN2(n7562), .Q(n7565) );
  XNOR3X1 U7570 ( .IN1(n7566), .IN2(n7509), .IN3(n7515), .Q(n7518) );
  XOR3X1 U7571 ( .IN1(n7521), .IN2(n7520), .IN3(n7519), .Q(n7515) );
  XNOR3X1 U7572 ( .IN1(n7530), .IN2(n7531), .IN3(n7533), .Q(n7519) );
  NAND2X0 U7573 ( .IN1(n7567), .IN2(n7568), .QN(n7533) );
  MUX21X1 U7574 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1501 ), .Q(n7568) );
  MUX21X1 U7575 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1502 ), .Q(n7567) );
  NAND2X0 U7576 ( .IN1(n7569), .IN2(n7570), .QN(n7531) );
  MUX21X1 U7577 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1506 ), .Q(n7570) );
  MUX21X1 U7578 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1505 ), .Q(n7569) );
  NAND2X0 U7579 ( .IN1(n7571), .IN2(n7572), .QN(n7530) );
  MUX21X1 U7580 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1504 ), .Q(n7572) );
  MUX21X1 U7581 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1503 ), .Q(n7571) );
  AOI22X1 U7582 ( .IN1(n7573), .IN2(n7574), .IN3(n7575), .IN4(n7576), .QN(
        n7520) );
  OR2X1 U7583 ( .IN1(n7574), .IN2(n7573), .Q(n7575) );
  XNOR3X1 U7584 ( .IN1(n7545), .IN2(n7546), .IN3(n7548), .Q(n7521) );
  NAND2X0 U7585 ( .IN1(n7577), .IN2(n7578), .QN(n7548) );
  MUX21X1 U7586 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1495 ), .Q(n7578) );
  MUX21X1 U7587 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1496 ), .Q(n7577) );
  NAND2X0 U7588 ( .IN1(n7579), .IN2(n7580), .QN(n7546) );
  MUX21X1 U7589 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1500 ), .Q(n7580) );
  MUX21X1 U7590 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1499 ), .Q(n7579) );
  NAND2X0 U7591 ( .IN1(n7581), .IN2(n7582), .QN(n7545) );
  MUX21X1 U7592 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1497 ), .Q(n7582) );
  MUX21X1 U7593 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1498 ), .Q(n7581) );
  XOR2X1 U7594 ( .IN1(n7471), .IN2(n7470), .Q(n7509) );
  NAND2X0 U7595 ( .IN1(n7583), .IN2(n7584), .QN(n7470) );
  MUX21X1 U7596 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1492 ), .Q(n7584) );
  MUX21X1 U7597 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1491 ), .Q(n7583) );
  NAND2X0 U7598 ( .IN1(n7585), .IN2(n7586), .QN(n7471) );
  MUX21X1 U7599 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1494 ), .Q(n7586) );
  MUX21X1 U7600 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1493 ), .Q(n7585) );
  XOR2X1 U7601 ( .IN1(n7510), .IN2(n7587), .Q(n7566) );
  NAND2X0 U7602 ( .IN1(n7513), .IN2(n7514), .QN(n7587) );
  AO22X1 U7603 ( .IN1(n7588), .IN2(n7589), .IN3(n7590), .IN4(n7591), .Q(n7510)
         );
  OR2X1 U7604 ( .IN1(n7589), .IN2(n7588), .Q(n7590) );
  AO22X1 U7605 ( .IN1(n7592), .IN2(n7593), .IN3(n7594), .IN4(n6189), .Q(
        \i_m4stg_frac/a0cout[38] ) );
  AO22X1 U7606 ( .IN1(n7595), .IN2(n7596), .IN3(n7597), .IN4(n7598), .Q(n6189)
         );
  OR2X1 U7607 ( .IN1(n7595), .IN2(n7596), .Q(n7598) );
  AND2X1 U7608 ( .IN1(n7599), .IN2(n7600), .Q(n7597) );
  NAND2X0 U7609 ( .IN1(n6190), .IN2(n6188), .QN(n7594) );
  INVX0 U7610 ( .INP(n7592), .ZN(n6188) );
  INVX0 U7611 ( .INP(n6190), .ZN(n7593) );
  MUX21X1 U7612 ( .IN1(n7601), .IN2(n7602), .S(n7603), .Q(n6190) );
  INVX0 U7613 ( .INP(n7604), .ZN(n7603) );
  XOR2X1 U7614 ( .IN1(n7561), .IN2(n7559), .Q(n7592) );
  OA22X1 U7615 ( .IN1(n7605), .IN2(n7606), .IN3(n7607), .IN4(n7608), .Q(n7559)
         );
  AND2X1 U7616 ( .IN1(n7606), .IN2(n7605), .Q(n7608) );
  XNOR3X1 U7617 ( .IN1(n7609), .IN2(n7552), .IN3(n7558), .Q(n7561) );
  XOR3X1 U7618 ( .IN1(n7564), .IN2(n7563), .IN3(n7562), .Q(n7558) );
  XNOR3X1 U7619 ( .IN1(n7573), .IN2(n7574), .IN3(n7576), .Q(n7562) );
  NAND2X0 U7620 ( .IN1(n7610), .IN2(n7611), .QN(n7576) );
  MUX21X1 U7621 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1500 ), .Q(n7611) );
  MUX21X1 U7622 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1501 ), .Q(n7610) );
  NAND2X0 U7623 ( .IN1(n7612), .IN2(n7613), .QN(n7574) );
  MUX21X1 U7624 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1505 ), .Q(n7613) );
  MUX21X1 U7625 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1504 ), .Q(n7612) );
  NAND2X0 U7626 ( .IN1(n7614), .IN2(n7615), .QN(n7573) );
  MUX21X1 U7627 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1503 ), .Q(n7615) );
  MUX21X1 U7628 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1502 ), .Q(n7614) );
  AOI22X1 U7629 ( .IN1(n7616), .IN2(n7617), .IN3(n7618), .IN4(n7619), .QN(
        n7563) );
  OR2X1 U7630 ( .IN1(n7617), .IN2(n7616), .Q(n7618) );
  XNOR3X1 U7631 ( .IN1(n7588), .IN2(n7589), .IN3(n7591), .Q(n7564) );
  NAND2X0 U7632 ( .IN1(n7620), .IN2(n7621), .QN(n7591) );
  MUX21X1 U7633 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1494 ), .Q(n7621) );
  MUX21X1 U7634 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1495 ), .Q(n7620) );
  NAND2X0 U7635 ( .IN1(n7622), .IN2(n7623), .QN(n7589) );
  MUX21X1 U7636 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1499 ), .Q(n7623) );
  MUX21X1 U7637 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1498 ), .Q(n7622) );
  NAND2X0 U7638 ( .IN1(n7624), .IN2(n7625), .QN(n7588) );
  MUX21X1 U7639 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1496 ), .Q(n7625) );
  MUX21X1 U7640 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1497 ), .Q(n7624) );
  XOR2X1 U7641 ( .IN1(n7514), .IN2(n7513), .Q(n7552) );
  NAND2X0 U7642 ( .IN1(n7626), .IN2(n7627), .QN(n7513) );
  MUX21X1 U7643 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1491 ), .Q(n7627) );
  MUX21X1 U7644 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1490 ), .Q(n7626) );
  NAND2X0 U7645 ( .IN1(n7628), .IN2(n7629), .QN(n7514) );
  MUX21X1 U7646 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1493 ), .Q(n7629) );
  MUX21X1 U7647 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1492 ), .Q(n7628) );
  XOR2X1 U7648 ( .IN1(n7553), .IN2(n7630), .Q(n7609) );
  NAND2X0 U7649 ( .IN1(n7556), .IN2(n7557), .QN(n7630) );
  AO22X1 U7650 ( .IN1(n7631), .IN2(n7632), .IN3(n7633), .IN4(n7634), .Q(n7553)
         );
  OR2X1 U7651 ( .IN1(n7632), .IN2(n7631), .Q(n7633) );
  AO22X1 U7652 ( .IN1(n7635), .IN2(n7636), .IN3(n7637), .IN4(n6192), .Q(
        \i_m4stg_frac/a0cout[37] ) );
  AO22X1 U7653 ( .IN1(n7638), .IN2(n7639), .IN3(n7640), .IN4(n7641), .Q(n6192)
         );
  OR2X1 U7654 ( .IN1(n7638), .IN2(n7639), .Q(n7641) );
  AND2X1 U7655 ( .IN1(n7642), .IN2(n7643), .Q(n7640) );
  NAND2X0 U7656 ( .IN1(n6193), .IN2(n6191), .QN(n7637) );
  INVX0 U7657 ( .INP(n7635), .ZN(n6191) );
  INVX0 U7658 ( .INP(n6193), .ZN(n7636) );
  MUX21X1 U7659 ( .IN1(n7644), .IN2(n7645), .S(n7646), .Q(n6193) );
  INVX0 U7660 ( .INP(n7647), .ZN(n7646) );
  XOR2X1 U7661 ( .IN1(n7604), .IN2(n7602), .Q(n7635) );
  OA22X1 U7662 ( .IN1(n7648), .IN2(n7649), .IN3(n7650), .IN4(n7651), .Q(n7602)
         );
  AND2X1 U7663 ( .IN1(n7649), .IN2(n7648), .Q(n7651) );
  XNOR3X1 U7664 ( .IN1(n7652), .IN2(n7595), .IN3(n7601), .Q(n7604) );
  XOR3X1 U7665 ( .IN1(n7607), .IN2(n7606), .IN3(n7605), .Q(n7601) );
  XNOR3X1 U7666 ( .IN1(n7616), .IN2(n7617), .IN3(n7619), .Q(n7605) );
  NAND2X0 U7667 ( .IN1(n7653), .IN2(n7654), .QN(n7619) );
  MUX21X1 U7668 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1499 ), .Q(n7654) );
  MUX21X1 U7669 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1500 ), .Q(n7653) );
  NAND2X0 U7670 ( .IN1(n7655), .IN2(n7656), .QN(n7617) );
  MUX21X1 U7671 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1504 ), .Q(n7656) );
  MUX21X1 U7672 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1503 ), .Q(n7655) );
  NAND2X0 U7673 ( .IN1(n7657), .IN2(n7658), .QN(n7616) );
  MUX21X1 U7674 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1502 ), .Q(n7658) );
  MUX21X1 U7675 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1501 ), .Q(n7657) );
  AOI22X1 U7676 ( .IN1(n7659), .IN2(n7660), .IN3(n7661), .IN4(n7662), .QN(
        n7606) );
  OR2X1 U7677 ( .IN1(n7660), .IN2(n7659), .Q(n7661) );
  XNOR3X1 U7678 ( .IN1(n7631), .IN2(n7632), .IN3(n7634), .Q(n7607) );
  NAND2X0 U7679 ( .IN1(n7663), .IN2(n7664), .QN(n7634) );
  MUX21X1 U7680 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1493 ), .Q(n7664) );
  MUX21X1 U7681 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1494 ), .Q(n7663) );
  NAND2X0 U7682 ( .IN1(n7665), .IN2(n7666), .QN(n7632) );
  MUX21X1 U7683 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1498 ), .Q(n7666) );
  MUX21X1 U7684 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1497 ), .Q(n7665) );
  NAND2X0 U7685 ( .IN1(n7667), .IN2(n7668), .QN(n7631) );
  MUX21X1 U7686 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1495 ), .Q(n7668) );
  MUX21X1 U7687 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1496 ), .Q(n7667) );
  XOR2X1 U7688 ( .IN1(n7557), .IN2(n7556), .Q(n7595) );
  NAND2X0 U7689 ( .IN1(n7669), .IN2(n7670), .QN(n7556) );
  MUX21X1 U7690 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1490 ), .Q(n7670) );
  MUX21X1 U7691 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1489 ), .Q(n7669) );
  NAND2X0 U7692 ( .IN1(n7671), .IN2(n7672), .QN(n7557) );
  MUX21X1 U7693 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1492 ), .Q(n7672) );
  MUX21X1 U7694 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1491 ), .Q(n7671) );
  XOR2X1 U7695 ( .IN1(n7596), .IN2(n7673), .Q(n7652) );
  NAND2X0 U7696 ( .IN1(n7599), .IN2(n7600), .QN(n7673) );
  AO22X1 U7697 ( .IN1(n7674), .IN2(n7675), .IN3(n7676), .IN4(n7677), .Q(n7596)
         );
  OR2X1 U7698 ( .IN1(n7675), .IN2(n7674), .Q(n7676) );
  AO22X1 U7699 ( .IN1(n7678), .IN2(n7679), .IN3(n7680), .IN4(n6195), .Q(
        \i_m4stg_frac/a0cout[36] ) );
  AO22X1 U7700 ( .IN1(n7681), .IN2(n7682), .IN3(n7683), .IN4(n7684), .Q(n6195)
         );
  OR2X1 U7701 ( .IN1(n7681), .IN2(n7682), .Q(n7684) );
  AND2X1 U7702 ( .IN1(n7685), .IN2(n7686), .Q(n7683) );
  NAND2X0 U7703 ( .IN1(n6196), .IN2(n6194), .QN(n7680) );
  INVX0 U7704 ( .INP(n7678), .ZN(n6194) );
  INVX0 U7705 ( .INP(n6196), .ZN(n7679) );
  MUX21X1 U7706 ( .IN1(n7687), .IN2(n7688), .S(n7689), .Q(n6196) );
  INVX0 U7707 ( .INP(n7690), .ZN(n7689) );
  XOR2X1 U7708 ( .IN1(n7647), .IN2(n7645), .Q(n7678) );
  OA22X1 U7709 ( .IN1(n7691), .IN2(n7692), .IN3(n7693), .IN4(n7694), .Q(n7645)
         );
  AND2X1 U7710 ( .IN1(n7692), .IN2(n7691), .Q(n7694) );
  XNOR3X1 U7711 ( .IN1(n7695), .IN2(n7638), .IN3(n7644), .Q(n7647) );
  XOR3X1 U7712 ( .IN1(n7650), .IN2(n7649), .IN3(n7648), .Q(n7644) );
  XNOR3X1 U7713 ( .IN1(n7659), .IN2(n7660), .IN3(n7662), .Q(n7648) );
  NAND2X0 U7714 ( .IN1(n7696), .IN2(n7697), .QN(n7662) );
  MUX21X1 U7715 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1498 ), .Q(n7697) );
  MUX21X1 U7716 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1499 ), .Q(n7696) );
  NAND2X0 U7717 ( .IN1(n7698), .IN2(n7699), .QN(n7660) );
  MUX21X1 U7718 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1503 ), .Q(n7699) );
  MUX21X1 U7719 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1502 ), .Q(n7698) );
  NAND2X0 U7720 ( .IN1(n7700), .IN2(n7701), .QN(n7659) );
  MUX21X1 U7721 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1501 ), .Q(n7701) );
  MUX21X1 U7722 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1500 ), .Q(n7700) );
  AOI22X1 U7723 ( .IN1(n7702), .IN2(n7703), .IN3(n7704), .IN4(n7705), .QN(
        n7649) );
  OR2X1 U7724 ( .IN1(n7703), .IN2(n7702), .Q(n7704) );
  XNOR3X1 U7725 ( .IN1(n7674), .IN2(n7675), .IN3(n7677), .Q(n7650) );
  NAND2X0 U7726 ( .IN1(n7706), .IN2(n7707), .QN(n7677) );
  MUX21X1 U7727 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1492 ), .Q(n7707) );
  MUX21X1 U7728 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1493 ), .Q(n7706) );
  NAND2X0 U7729 ( .IN1(n7708), .IN2(n7709), .QN(n7675) );
  MUX21X1 U7730 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1497 ), .Q(n7709) );
  MUX21X1 U7731 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1496 ), .Q(n7708) );
  NAND2X0 U7732 ( .IN1(n7710), .IN2(n7711), .QN(n7674) );
  MUX21X1 U7733 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1494 ), .Q(n7711) );
  MUX21X1 U7734 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1495 ), .Q(n7710) );
  XOR2X1 U7735 ( .IN1(n7600), .IN2(n7599), .Q(n7638) );
  NAND2X0 U7736 ( .IN1(n7712), .IN2(n7713), .QN(n7599) );
  MUX21X1 U7737 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1489 ), .Q(n7713) );
  MUX21X1 U7738 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1488 ), .Q(n7712) );
  NAND2X0 U7739 ( .IN1(n7714), .IN2(n7715), .QN(n7600) );
  MUX21X1 U7740 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1491 ), .Q(n7715) );
  MUX21X1 U7741 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1490 ), .Q(n7714) );
  XOR2X1 U7742 ( .IN1(n7639), .IN2(n7716), .Q(n7695) );
  NAND2X0 U7743 ( .IN1(n7642), .IN2(n7643), .QN(n7716) );
  AO22X1 U7744 ( .IN1(n7717), .IN2(n7718), .IN3(n7719), .IN4(n7720), .Q(n7639)
         );
  OR2X1 U7745 ( .IN1(n7718), .IN2(n7717), .Q(n7719) );
  AO22X1 U7746 ( .IN1(n7721), .IN2(n7722), .IN3(n7723), .IN4(n6198), .Q(
        \i_m4stg_frac/a0cout[35] ) );
  AO22X1 U7747 ( .IN1(n7724), .IN2(n7725), .IN3(n7726), .IN4(n7727), .Q(n6198)
         );
  OR2X1 U7748 ( .IN1(n7724), .IN2(n7725), .Q(n7727) );
  AND2X1 U7749 ( .IN1(n7728), .IN2(n7729), .Q(n7726) );
  NAND2X0 U7750 ( .IN1(n6199), .IN2(n6197), .QN(n7723) );
  INVX0 U7751 ( .INP(n7721), .ZN(n6197) );
  INVX0 U7752 ( .INP(n6199), .ZN(n7722) );
  MUX21X1 U7753 ( .IN1(n7730), .IN2(n7731), .S(n7732), .Q(n6199) );
  INVX0 U7754 ( .INP(n7733), .ZN(n7732) );
  XOR2X1 U7755 ( .IN1(n7690), .IN2(n7688), .Q(n7721) );
  OA22X1 U7756 ( .IN1(n7734), .IN2(n7735), .IN3(n7736), .IN4(n7737), .Q(n7688)
         );
  AND2X1 U7757 ( .IN1(n7735), .IN2(n7734), .Q(n7737) );
  XNOR3X1 U7758 ( .IN1(n7738), .IN2(n7681), .IN3(n7687), .Q(n7690) );
  XOR3X1 U7759 ( .IN1(n7693), .IN2(n7692), .IN3(n7691), .Q(n7687) );
  XNOR3X1 U7760 ( .IN1(n7702), .IN2(n7703), .IN3(n7705), .Q(n7691) );
  NAND2X0 U7761 ( .IN1(n7739), .IN2(n7740), .QN(n7705) );
  MUX21X1 U7762 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1497 ), .Q(n7740) );
  MUX21X1 U7763 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1498 ), .Q(n7739) );
  NAND2X0 U7764 ( .IN1(n7741), .IN2(n7742), .QN(n7703) );
  MUX21X1 U7765 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1502 ), .Q(n7742) );
  MUX21X1 U7766 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1501 ), .Q(n7741) );
  NAND2X0 U7767 ( .IN1(n7743), .IN2(n7744), .QN(n7702) );
  MUX21X1 U7768 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1500 ), .Q(n7744) );
  MUX21X1 U7769 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1499 ), .Q(n7743) );
  AOI22X1 U7770 ( .IN1(n7745), .IN2(n7746), .IN3(n7747), .IN4(n7748), .QN(
        n7692) );
  OR2X1 U7771 ( .IN1(n7746), .IN2(n7745), .Q(n7747) );
  XNOR3X1 U7772 ( .IN1(n7717), .IN2(n7718), .IN3(n7720), .Q(n7693) );
  NAND2X0 U7773 ( .IN1(n7749), .IN2(n7750), .QN(n7720) );
  MUX21X1 U7774 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1491 ), .Q(n7750) );
  MUX21X1 U7775 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1492 ), .Q(n7749) );
  NAND2X0 U7776 ( .IN1(n7751), .IN2(n7752), .QN(n7718) );
  MUX21X1 U7777 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1496 ), .Q(n7752) );
  MUX21X1 U7778 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1495 ), .Q(n7751) );
  NAND2X0 U7779 ( .IN1(n7753), .IN2(n7754), .QN(n7717) );
  MUX21X1 U7780 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1493 ), .Q(n7754) );
  MUX21X1 U7781 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1494 ), .Q(n7753) );
  XOR2X1 U7782 ( .IN1(n7643), .IN2(n7642), .Q(n7681) );
  NAND2X0 U7783 ( .IN1(n7755), .IN2(n7756), .QN(n7642) );
  MUX21X1 U7784 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1488 ), .Q(n7756) );
  MUX21X1 U7785 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1487 ), .Q(n7755) );
  NAND2X0 U7786 ( .IN1(n7757), .IN2(n7758), .QN(n7643) );
  MUX21X1 U7787 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1490 ), .Q(n7758) );
  MUX21X1 U7788 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1489 ), .Q(n7757) );
  XOR2X1 U7789 ( .IN1(n7682), .IN2(n7759), .Q(n7738) );
  NAND2X0 U7790 ( .IN1(n7685), .IN2(n7686), .QN(n7759) );
  AO22X1 U7791 ( .IN1(n7760), .IN2(n7761), .IN3(n7762), .IN4(n7763), .Q(n7682)
         );
  OR2X1 U7792 ( .IN1(n7761), .IN2(n7760), .Q(n7762) );
  AO22X1 U7793 ( .IN1(n7764), .IN2(n7765), .IN3(n7766), .IN4(n6201), .Q(
        \i_m4stg_frac/a0cout[34] ) );
  AO22X1 U7794 ( .IN1(n7767), .IN2(n7768), .IN3(n7769), .IN4(n7770), .Q(n6201)
         );
  OR2X1 U7795 ( .IN1(n7767), .IN2(n7768), .Q(n7770) );
  AND2X1 U7796 ( .IN1(n7771), .IN2(n7772), .Q(n7769) );
  NAND2X0 U7797 ( .IN1(n6202), .IN2(n6200), .QN(n7766) );
  INVX0 U7798 ( .INP(n7764), .ZN(n6200) );
  INVX0 U7799 ( .INP(n6202), .ZN(n7765) );
  MUX21X1 U7800 ( .IN1(n7773), .IN2(n7774), .S(n7775), .Q(n6202) );
  INVX0 U7801 ( .INP(n7776), .ZN(n7775) );
  XOR2X1 U7802 ( .IN1(n7733), .IN2(n7731), .Q(n7764) );
  OA22X1 U7803 ( .IN1(n7777), .IN2(n7778), .IN3(n7779), .IN4(n7780), .Q(n7731)
         );
  AND2X1 U7804 ( .IN1(n7778), .IN2(n7777), .Q(n7780) );
  XNOR3X1 U7805 ( .IN1(n7781), .IN2(n7724), .IN3(n7730), .Q(n7733) );
  XOR3X1 U7806 ( .IN1(n7736), .IN2(n7735), .IN3(n7734), .Q(n7730) );
  XNOR3X1 U7807 ( .IN1(n7745), .IN2(n7746), .IN3(n7748), .Q(n7734) );
  NAND2X0 U7808 ( .IN1(n7782), .IN2(n7783), .QN(n7748) );
  MUX21X1 U7809 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1496 ), .Q(n7783) );
  MUX21X1 U7810 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1497 ), .Q(n7782) );
  NAND2X0 U7811 ( .IN1(n7784), .IN2(n7785), .QN(n7746) );
  MUX21X1 U7812 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1501 ), .Q(n7785) );
  MUX21X1 U7813 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1500 ), .Q(n7784) );
  NAND2X0 U7814 ( .IN1(n7786), .IN2(n7787), .QN(n7745) );
  MUX21X1 U7815 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1499 ), .Q(n7787) );
  MUX21X1 U7816 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1498 ), .Q(n7786) );
  AOI22X1 U7817 ( .IN1(n7788), .IN2(n7789), .IN3(n7790), .IN4(n7791), .QN(
        n7735) );
  OR2X1 U7818 ( .IN1(n7789), .IN2(n7788), .Q(n7790) );
  XNOR3X1 U7819 ( .IN1(n7760), .IN2(n7761), .IN3(n7763), .Q(n7736) );
  NAND2X0 U7820 ( .IN1(n7792), .IN2(n7793), .QN(n7763) );
  MUX21X1 U7821 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1490 ), .Q(n7793) );
  MUX21X1 U7822 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1491 ), .Q(n7792) );
  NAND2X0 U7823 ( .IN1(n7794), .IN2(n7795), .QN(n7761) );
  MUX21X1 U7824 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1495 ), .Q(n7795) );
  MUX21X1 U7825 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1494 ), .Q(n7794) );
  NAND2X0 U7826 ( .IN1(n7796), .IN2(n7797), .QN(n7760) );
  MUX21X1 U7827 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1492 ), .Q(n7797) );
  MUX21X1 U7828 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1493 ), .Q(n7796) );
  XOR2X1 U7829 ( .IN1(n7686), .IN2(n7685), .Q(n7724) );
  NAND2X0 U7830 ( .IN1(n7798), .IN2(n7799), .QN(n7685) );
  MUX21X1 U7831 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1487 ), .Q(n7799) );
  MUX21X1 U7832 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1486 ), .Q(n7798) );
  NAND2X0 U7833 ( .IN1(n7800), .IN2(n7801), .QN(n7686) );
  MUX21X1 U7834 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1489 ), .Q(n7801) );
  MUX21X1 U7835 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1488 ), .Q(n7800) );
  XOR2X1 U7836 ( .IN1(n7725), .IN2(n7802), .Q(n7781) );
  NAND2X0 U7837 ( .IN1(n7728), .IN2(n7729), .QN(n7802) );
  AO22X1 U7838 ( .IN1(n7803), .IN2(n7804), .IN3(n7805), .IN4(n7806), .Q(n7725)
         );
  OR2X1 U7839 ( .IN1(n7804), .IN2(n7803), .Q(n7805) );
  AO22X1 U7840 ( .IN1(n7807), .IN2(n7808), .IN3(n7809), .IN4(n6204), .Q(
        \i_m4stg_frac/a0cout[33] ) );
  AO22X1 U7841 ( .IN1(n7810), .IN2(n7811), .IN3(n7812), .IN4(n7813), .Q(n6204)
         );
  OR2X1 U7842 ( .IN1(n7810), .IN2(n7811), .Q(n7813) );
  AND2X1 U7843 ( .IN1(n7814), .IN2(n7815), .Q(n7812) );
  NAND2X0 U7844 ( .IN1(n6205), .IN2(n6203), .QN(n7809) );
  INVX0 U7845 ( .INP(n7807), .ZN(n6203) );
  INVX0 U7846 ( .INP(n6205), .ZN(n7808) );
  MUX21X1 U7847 ( .IN1(n7816), .IN2(n7817), .S(n7818), .Q(n6205) );
  INVX0 U7848 ( .INP(n7819), .ZN(n7818) );
  XOR2X1 U7849 ( .IN1(n7776), .IN2(n7774), .Q(n7807) );
  OA22X1 U7850 ( .IN1(n7820), .IN2(n7821), .IN3(n7822), .IN4(n7823), .Q(n7774)
         );
  AND2X1 U7851 ( .IN1(n7821), .IN2(n7820), .Q(n7823) );
  XNOR3X1 U7852 ( .IN1(n7824), .IN2(n7767), .IN3(n7773), .Q(n7776) );
  XOR3X1 U7853 ( .IN1(n7779), .IN2(n7778), .IN3(n7777), .Q(n7773) );
  XNOR3X1 U7854 ( .IN1(n7788), .IN2(n7789), .IN3(n7791), .Q(n7777) );
  NAND2X0 U7855 ( .IN1(n7825), .IN2(n7826), .QN(n7791) );
  MUX21X1 U7856 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1495 ), .Q(n7826) );
  MUX21X1 U7857 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1496 ), .Q(n7825) );
  NAND2X0 U7858 ( .IN1(n7827), .IN2(n7828), .QN(n7789) );
  MUX21X1 U7859 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1500 ), .Q(n7828) );
  MUX21X1 U7860 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1499 ), .Q(n7827) );
  NAND2X0 U7861 ( .IN1(n7829), .IN2(n7830), .QN(n7788) );
  MUX21X1 U7862 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1498 ), .Q(n7830) );
  MUX21X1 U7863 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1497 ), .Q(n7829) );
  AOI22X1 U7864 ( .IN1(n7831), .IN2(n7832), .IN3(n7833), .IN4(n7834), .QN(
        n7778) );
  OR2X1 U7865 ( .IN1(n7832), .IN2(n7831), .Q(n7833) );
  XNOR3X1 U7866 ( .IN1(n7803), .IN2(n7804), .IN3(n7806), .Q(n7779) );
  NAND2X0 U7867 ( .IN1(n7835), .IN2(n7836), .QN(n7806) );
  MUX21X1 U7868 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1489 ), .Q(n7836) );
  MUX21X1 U7869 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1490 ), .Q(n7835) );
  NAND2X0 U7870 ( .IN1(n7837), .IN2(n7838), .QN(n7804) );
  MUX21X1 U7871 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1494 ), .Q(n7838) );
  MUX21X1 U7872 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1493 ), .Q(n7837) );
  NAND2X0 U7873 ( .IN1(n7839), .IN2(n7840), .QN(n7803) );
  MUX21X1 U7874 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1491 ), .Q(n7840) );
  MUX21X1 U7875 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1492 ), .Q(n7839) );
  XOR2X1 U7876 ( .IN1(n7729), .IN2(n7728), .Q(n7767) );
  NAND2X0 U7877 ( .IN1(n7841), .IN2(n7842), .QN(n7728) );
  MUX21X1 U7878 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1486 ), .Q(n7842) );
  MUX21X1 U7879 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1485 ), .Q(n7841) );
  NAND2X0 U7880 ( .IN1(n7843), .IN2(n7844), .QN(n7729) );
  MUX21X1 U7881 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1488 ), .Q(n7844) );
  MUX21X1 U7882 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1487 ), .Q(n7843) );
  XOR2X1 U7883 ( .IN1(n7768), .IN2(n7845), .Q(n7824) );
  NAND2X0 U7884 ( .IN1(n7771), .IN2(n7772), .QN(n7845) );
  AO22X1 U7885 ( .IN1(n7846), .IN2(n7847), .IN3(n7848), .IN4(n7849), .Q(n7768)
         );
  OR2X1 U7886 ( .IN1(n7847), .IN2(n7846), .Q(n7848) );
  AO22X1 U7887 ( .IN1(n7850), .IN2(n7851), .IN3(n7852), .IN4(n6207), .Q(
        \i_m4stg_frac/a0cout[32] ) );
  AO22X1 U7888 ( .IN1(n7853), .IN2(n7854), .IN3(n7855), .IN4(n7856), .Q(n6207)
         );
  OR2X1 U7889 ( .IN1(n7853), .IN2(n7854), .Q(n7856) );
  AND2X1 U7890 ( .IN1(n7857), .IN2(n7858), .Q(n7855) );
  NAND2X0 U7891 ( .IN1(n6208), .IN2(n6206), .QN(n7852) );
  INVX0 U7892 ( .INP(n7850), .ZN(n6206) );
  INVX0 U7893 ( .INP(n6208), .ZN(n7851) );
  MUX21X1 U7894 ( .IN1(n7859), .IN2(n7860), .S(n7861), .Q(n6208) );
  INVX0 U7895 ( .INP(n7862), .ZN(n7861) );
  XOR2X1 U7896 ( .IN1(n7819), .IN2(n7817), .Q(n7850) );
  OA22X1 U7897 ( .IN1(n7863), .IN2(n7864), .IN3(n7865), .IN4(n7866), .Q(n7817)
         );
  AND2X1 U7898 ( .IN1(n7864), .IN2(n7863), .Q(n7866) );
  XNOR3X1 U7899 ( .IN1(n7867), .IN2(n7810), .IN3(n7816), .Q(n7819) );
  XOR3X1 U7900 ( .IN1(n7822), .IN2(n7821), .IN3(n7820), .Q(n7816) );
  XNOR3X1 U7901 ( .IN1(n7831), .IN2(n7832), .IN3(n7834), .Q(n7820) );
  NAND2X0 U7902 ( .IN1(n7868), .IN2(n7869), .QN(n7834) );
  MUX21X1 U7903 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1494 ), .Q(n7869) );
  MUX21X1 U7904 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1495 ), .Q(n7868) );
  NAND2X0 U7905 ( .IN1(n7870), .IN2(n7871), .QN(n7832) );
  MUX21X1 U7906 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1499 ), .Q(n7871) );
  MUX21X1 U7907 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1498 ), .Q(n7870) );
  NAND2X0 U7908 ( .IN1(n7872), .IN2(n7873), .QN(n7831) );
  MUX21X1 U7909 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1497 ), .Q(n7873) );
  MUX21X1 U7910 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1496 ), .Q(n7872) );
  AOI22X1 U7911 ( .IN1(n7874), .IN2(n7875), .IN3(n7876), .IN4(n7877), .QN(
        n7821) );
  OR2X1 U7912 ( .IN1(n7875), .IN2(n7874), .Q(n7876) );
  XNOR3X1 U7913 ( .IN1(n7846), .IN2(n7847), .IN3(n7849), .Q(n7822) );
  NAND2X0 U7914 ( .IN1(n7878), .IN2(n7879), .QN(n7849) );
  MUX21X1 U7915 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1488 ), .Q(n7879) );
  MUX21X1 U7916 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1489 ), .Q(n7878) );
  NAND2X0 U7917 ( .IN1(n7880), .IN2(n7881), .QN(n7847) );
  MUX21X1 U7918 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1493 ), .Q(n7881) );
  MUX21X1 U7919 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1492 ), .Q(n7880) );
  NAND2X0 U7920 ( .IN1(n7882), .IN2(n7883), .QN(n7846) );
  MUX21X1 U7921 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1490 ), .Q(n7883) );
  MUX21X1 U7922 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1491 ), .Q(n7882) );
  XOR2X1 U7923 ( .IN1(n7772), .IN2(n7771), .Q(n7810) );
  NAND2X0 U7924 ( .IN1(n7884), .IN2(n7885), .QN(n7771) );
  MUX21X1 U7925 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1485 ), .Q(n7885) );
  MUX21X1 U7926 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1484 ), .Q(n7884) );
  NAND2X0 U7927 ( .IN1(n7886), .IN2(n7887), .QN(n7772) );
  MUX21X1 U7928 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1487 ), .Q(n7887) );
  MUX21X1 U7929 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1486 ), .Q(n7886) );
  XOR2X1 U7930 ( .IN1(n7811), .IN2(n7888), .Q(n7867) );
  NAND2X0 U7931 ( .IN1(n7814), .IN2(n7815), .QN(n7888) );
  AO22X1 U7932 ( .IN1(n7889), .IN2(n7890), .IN3(n7891), .IN4(n7892), .Q(n7811)
         );
  OR2X1 U7933 ( .IN1(n7890), .IN2(n7889), .Q(n7891) );
  AO22X1 U7934 ( .IN1(n7893), .IN2(n7894), .IN3(n7895), .IN4(n6210), .Q(
        \i_m4stg_frac/a0cout[31] ) );
  AO22X1 U7935 ( .IN1(n7896), .IN2(n7897), .IN3(n7898), .IN4(n7899), .Q(n6210)
         );
  OR2X1 U7936 ( .IN1(n7896), .IN2(n7897), .Q(n7899) );
  AND2X1 U7937 ( .IN1(n7900), .IN2(n7901), .Q(n7898) );
  NAND2X0 U7938 ( .IN1(n6211), .IN2(n6209), .QN(n7895) );
  INVX0 U7939 ( .INP(n7893), .ZN(n6209) );
  INVX0 U7940 ( .INP(n6211), .ZN(n7894) );
  MUX21X1 U7941 ( .IN1(n7902), .IN2(n7903), .S(n7904), .Q(n6211) );
  INVX0 U7942 ( .INP(n7905), .ZN(n7904) );
  XOR2X1 U7943 ( .IN1(n7862), .IN2(n7860), .Q(n7893) );
  OA22X1 U7944 ( .IN1(n7906), .IN2(n7907), .IN3(n7908), .IN4(n7909), .Q(n7860)
         );
  AND2X1 U7945 ( .IN1(n7907), .IN2(n7906), .Q(n7909) );
  XNOR3X1 U7946 ( .IN1(n7910), .IN2(n7853), .IN3(n7859), .Q(n7862) );
  XOR3X1 U7947 ( .IN1(n7865), .IN2(n7864), .IN3(n7863), .Q(n7859) );
  XNOR3X1 U7948 ( .IN1(n7874), .IN2(n7875), .IN3(n7877), .Q(n7863) );
  NAND2X0 U7949 ( .IN1(n7911), .IN2(n7912), .QN(n7877) );
  MUX21X1 U7950 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1493 ), .Q(n7912) );
  MUX21X1 U7951 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1494 ), .Q(n7911) );
  NAND2X0 U7952 ( .IN1(n7913), .IN2(n7914), .QN(n7875) );
  MUX21X1 U7953 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1498 ), .Q(n7914) );
  MUX21X1 U7954 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1497 ), .Q(n7913) );
  NAND2X0 U7955 ( .IN1(n7915), .IN2(n7916), .QN(n7874) );
  MUX21X1 U7956 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1496 ), .Q(n7916) );
  MUX21X1 U7957 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1495 ), .Q(n7915) );
  AOI22X1 U7958 ( .IN1(n7917), .IN2(n7918), .IN3(n7919), .IN4(n7920), .QN(
        n7864) );
  OR2X1 U7959 ( .IN1(n7918), .IN2(n7917), .Q(n7919) );
  XNOR3X1 U7960 ( .IN1(n7889), .IN2(n7890), .IN3(n7892), .Q(n7865) );
  NAND2X0 U7961 ( .IN1(n7921), .IN2(n7922), .QN(n7892) );
  MUX21X1 U7962 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1487 ), .Q(n7922) );
  MUX21X1 U7963 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1488 ), .Q(n7921) );
  NAND2X0 U7964 ( .IN1(n7923), .IN2(n7924), .QN(n7890) );
  MUX21X1 U7965 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1492 ), .Q(n7924) );
  MUX21X1 U7966 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1491 ), .Q(n7923) );
  NAND2X0 U7967 ( .IN1(n7925), .IN2(n7926), .QN(n7889) );
  MUX21X1 U7968 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1489 ), .Q(n7926) );
  MUX21X1 U7969 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1490 ), .Q(n7925) );
  XOR2X1 U7970 ( .IN1(n7815), .IN2(n7814), .Q(n7853) );
  NAND2X0 U7971 ( .IN1(n7927), .IN2(n7928), .QN(n7814) );
  MUX21X1 U7972 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1484 ), .Q(n7928) );
  MUX21X1 U7973 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1483 ), .Q(n7927) );
  NAND2X0 U7974 ( .IN1(n7929), .IN2(n7930), .QN(n7815) );
  MUX21X1 U7975 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1486 ), .Q(n7930) );
  MUX21X1 U7976 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1485 ), .Q(n7929) );
  XOR2X1 U7977 ( .IN1(n7854), .IN2(n7931), .Q(n7910) );
  NAND2X0 U7978 ( .IN1(n7857), .IN2(n7858), .QN(n7931) );
  AO22X1 U7979 ( .IN1(n7932), .IN2(n7933), .IN3(n7934), .IN4(n7935), .Q(n7854)
         );
  OR2X1 U7980 ( .IN1(n7933), .IN2(n7932), .Q(n7934) );
  AO22X1 U7981 ( .IN1(n7936), .IN2(n7937), .IN3(n7938), .IN4(n6213), .Q(
        \i_m4stg_frac/a0cout[30] ) );
  AO22X1 U7982 ( .IN1(n7939), .IN2(n7940), .IN3(n7941), .IN4(n7942), .Q(n6213)
         );
  OR2X1 U7983 ( .IN1(n7939), .IN2(n7940), .Q(n7942) );
  AND2X1 U7984 ( .IN1(n7943), .IN2(n7944), .Q(n7941) );
  NAND2X0 U7985 ( .IN1(n6214), .IN2(n6212), .QN(n7938) );
  INVX0 U7986 ( .INP(n7936), .ZN(n6212) );
  INVX0 U7987 ( .INP(n6214), .ZN(n7937) );
  MUX21X1 U7988 ( .IN1(n7945), .IN2(n7946), .S(n7947), .Q(n6214) );
  INVX0 U7989 ( .INP(n7948), .ZN(n7947) );
  XOR2X1 U7990 ( .IN1(n7905), .IN2(n7903), .Q(n7936) );
  OA22X1 U7991 ( .IN1(n7949), .IN2(n7950), .IN3(n7951), .IN4(n7952), .Q(n7903)
         );
  AND2X1 U7992 ( .IN1(n7950), .IN2(n7949), .Q(n7952) );
  XNOR3X1 U7993 ( .IN1(n7953), .IN2(n7896), .IN3(n7902), .Q(n7905) );
  XOR3X1 U7994 ( .IN1(n7908), .IN2(n7907), .IN3(n7906), .Q(n7902) );
  XNOR3X1 U7995 ( .IN1(n7917), .IN2(n7918), .IN3(n7920), .Q(n7906) );
  NAND2X0 U7996 ( .IN1(n7954), .IN2(n7955), .QN(n7920) );
  MUX21X1 U7997 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1492 ), .Q(n7955) );
  MUX21X1 U7998 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1493 ), .Q(n7954) );
  NAND2X0 U7999 ( .IN1(n7956), .IN2(n7957), .QN(n7918) );
  MUX21X1 U8000 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1497 ), .Q(n7957) );
  MUX21X1 U8001 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1496 ), .Q(n7956) );
  NAND2X0 U8002 ( .IN1(n7958), .IN2(n7959), .QN(n7917) );
  MUX21X1 U8003 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1495 ), .Q(n7959) );
  MUX21X1 U8004 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1494 ), .Q(n7958) );
  AOI22X1 U8005 ( .IN1(n7960), .IN2(n7961), .IN3(n7962), .IN4(n7963), .QN(
        n7907) );
  OR2X1 U8006 ( .IN1(n7961), .IN2(n7960), .Q(n7962) );
  XNOR3X1 U8007 ( .IN1(n7932), .IN2(n7933), .IN3(n7935), .Q(n7908) );
  NAND2X0 U8008 ( .IN1(n7964), .IN2(n7965), .QN(n7935) );
  MUX21X1 U8009 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1486 ), .Q(n7965) );
  MUX21X1 U8010 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1487 ), .Q(n7964) );
  NAND2X0 U8011 ( .IN1(n7966), .IN2(n7967), .QN(n7933) );
  MUX21X1 U8012 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1491 ), .Q(n7967) );
  MUX21X1 U8013 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1490 ), .Q(n7966) );
  NAND2X0 U8014 ( .IN1(n7968), .IN2(n7969), .QN(n7932) );
  MUX21X1 U8015 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1488 ), .Q(n7969) );
  MUX21X1 U8016 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1489 ), .Q(n7968) );
  XOR2X1 U8017 ( .IN1(n7858), .IN2(n7857), .Q(n7896) );
  NAND2X0 U8018 ( .IN1(n7970), .IN2(n7971), .QN(n7857) );
  MUX21X1 U8019 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1483 ), .Q(n7971) );
  MUX21X1 U8020 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1482 ), .Q(n7970) );
  NAND2X0 U8021 ( .IN1(n7972), .IN2(n7973), .QN(n7858) );
  MUX21X1 U8022 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1485 ), .Q(n7973) );
  MUX21X1 U8023 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1484 ), .Q(n7972) );
  XOR2X1 U8024 ( .IN1(n7897), .IN2(n7974), .Q(n7953) );
  NAND2X0 U8025 ( .IN1(n7900), .IN2(n7901), .QN(n7974) );
  AO22X1 U8026 ( .IN1(n7975), .IN2(n7976), .IN3(n7977), .IN4(n7978), .Q(n7897)
         );
  OR2X1 U8027 ( .IN1(n7976), .IN2(n7975), .Q(n7977) );
  AO22X1 U8028 ( .IN1(n7979), .IN2(n7980), .IN3(n7981), .IN4(n6218), .Q(
        \i_m4stg_frac/a0cout[29] ) );
  AO22X1 U8029 ( .IN1(n7982), .IN2(n7983), .IN3(n7984), .IN4(n7985), .Q(n6218)
         );
  OR2X1 U8030 ( .IN1(n7982), .IN2(n7983), .Q(n7985) );
  AND2X1 U8031 ( .IN1(n7986), .IN2(n7987), .Q(n7984) );
  NAND2X0 U8032 ( .IN1(n6219), .IN2(n6217), .QN(n7981) );
  INVX0 U8033 ( .INP(n7979), .ZN(n6217) );
  INVX0 U8034 ( .INP(n6219), .ZN(n7980) );
  MUX21X1 U8035 ( .IN1(n7988), .IN2(n7989), .S(n7990), .Q(n6219) );
  INVX0 U8036 ( .INP(n7991), .ZN(n7990) );
  XOR2X1 U8037 ( .IN1(n7948), .IN2(n7946), .Q(n7979) );
  OA22X1 U8038 ( .IN1(n7992), .IN2(n7993), .IN3(n7994), .IN4(n7995), .Q(n7946)
         );
  AND2X1 U8039 ( .IN1(n7993), .IN2(n7992), .Q(n7995) );
  XNOR3X1 U8040 ( .IN1(n7996), .IN2(n7939), .IN3(n7945), .Q(n7948) );
  XOR3X1 U8041 ( .IN1(n7951), .IN2(n7950), .IN3(n7949), .Q(n7945) );
  XNOR3X1 U8042 ( .IN1(n7960), .IN2(n7961), .IN3(n7963), .Q(n7949) );
  NAND2X0 U8043 ( .IN1(n7997), .IN2(n7998), .QN(n7963) );
  MUX21X1 U8044 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1491 ), .Q(n7998) );
  MUX21X1 U8045 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1492 ), .Q(n7997) );
  NAND2X0 U8046 ( .IN1(n7999), .IN2(n8000), .QN(n7961) );
  MUX21X1 U8047 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1496 ), .Q(n8000) );
  MUX21X1 U8048 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1495 ), .Q(n7999) );
  NAND2X0 U8049 ( .IN1(n8001), .IN2(n8002), .QN(n7960) );
  MUX21X1 U8050 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1494 ), .Q(n8002) );
  MUX21X1 U8051 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1493 ), .Q(n8001) );
  AOI22X1 U8052 ( .IN1(n8003), .IN2(n8004), .IN3(n8005), .IN4(n8006), .QN(
        n7950) );
  OR2X1 U8053 ( .IN1(n8004), .IN2(n8003), .Q(n8005) );
  XNOR3X1 U8054 ( .IN1(n7975), .IN2(n7976), .IN3(n7978), .Q(n7951) );
  NAND2X0 U8055 ( .IN1(n8007), .IN2(n8008), .QN(n7978) );
  MUX21X1 U8056 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1485 ), .Q(n8008) );
  MUX21X1 U8057 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1486 ), .Q(n8007) );
  NAND2X0 U8058 ( .IN1(n8009), .IN2(n8010), .QN(n7976) );
  MUX21X1 U8059 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1490 ), .Q(n8010) );
  MUX21X1 U8060 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1489 ), .Q(n8009) );
  NAND2X0 U8061 ( .IN1(n8011), .IN2(n8012), .QN(n7975) );
  MUX21X1 U8062 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1487 ), .Q(n8012) );
  MUX21X1 U8063 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1488 ), .Q(n8011) );
  XOR2X1 U8064 ( .IN1(n7901), .IN2(n7900), .Q(n7939) );
  NAND2X0 U8065 ( .IN1(n8013), .IN2(n8014), .QN(n7900) );
  MUX21X1 U8066 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1482 ), .Q(n8014) );
  MUX21X1 U8067 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1481 ), .Q(n8013) );
  NAND2X0 U8068 ( .IN1(n8015), .IN2(n8016), .QN(n7901) );
  MUX21X1 U8069 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1484 ), .Q(n8016) );
  MUX21X1 U8070 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1483 ), .Q(n8015) );
  XOR2X1 U8071 ( .IN1(n7940), .IN2(n8017), .Q(n7996) );
  NAND2X0 U8072 ( .IN1(n7943), .IN2(n7944), .QN(n8017) );
  AO22X1 U8073 ( .IN1(n8018), .IN2(n8019), .IN3(n8020), .IN4(n8021), .Q(n7940)
         );
  OR2X1 U8074 ( .IN1(n8019), .IN2(n8018), .Q(n8020) );
  AO22X1 U8075 ( .IN1(n8022), .IN2(n8023), .IN3(n8024), .IN4(n6221), .Q(
        \i_m4stg_frac/a0cout[28] ) );
  AO22X1 U8076 ( .IN1(n8025), .IN2(n8026), .IN3(n8027), .IN4(n8028), .Q(n6221)
         );
  OR2X1 U8077 ( .IN1(n8025), .IN2(n8026), .Q(n8028) );
  AND2X1 U8078 ( .IN1(n8029), .IN2(n8030), .Q(n8027) );
  NAND2X0 U8079 ( .IN1(n6222), .IN2(n6220), .QN(n8024) );
  INVX0 U8080 ( .INP(n8022), .ZN(n6220) );
  INVX0 U8081 ( .INP(n6222), .ZN(n8023) );
  MUX21X1 U8082 ( .IN1(n8031), .IN2(n8032), .S(n8033), .Q(n6222) );
  INVX0 U8083 ( .INP(n8034), .ZN(n8033) );
  XOR2X1 U8084 ( .IN1(n7991), .IN2(n7989), .Q(n8022) );
  OA22X1 U8085 ( .IN1(n8035), .IN2(n8036), .IN3(n8037), .IN4(n8038), .Q(n7989)
         );
  AND2X1 U8086 ( .IN1(n8036), .IN2(n8035), .Q(n8038) );
  XNOR3X1 U8087 ( .IN1(n8039), .IN2(n7982), .IN3(n7988), .Q(n7991) );
  XOR3X1 U8088 ( .IN1(n7994), .IN2(n7993), .IN3(n7992), .Q(n7988) );
  XNOR3X1 U8089 ( .IN1(n8003), .IN2(n8004), .IN3(n8006), .Q(n7992) );
  NAND2X0 U8090 ( .IN1(n8040), .IN2(n8041), .QN(n8006) );
  MUX21X1 U8091 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1490 ), .Q(n8041) );
  MUX21X1 U8092 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1491 ), .Q(n8040) );
  NAND2X0 U8093 ( .IN1(n8042), .IN2(n8043), .QN(n8004) );
  MUX21X1 U8094 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1495 ), .Q(n8043) );
  MUX21X1 U8095 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1494 ), .Q(n8042) );
  NAND2X0 U8096 ( .IN1(n8044), .IN2(n8045), .QN(n8003) );
  MUX21X1 U8097 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1493 ), .Q(n8045) );
  MUX21X1 U8098 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1492 ), .Q(n8044) );
  AOI22X1 U8099 ( .IN1(n8046), .IN2(n8047), .IN3(n8048), .IN4(n8049), .QN(
        n7993) );
  OR2X1 U8100 ( .IN1(n8047), .IN2(n8046), .Q(n8048) );
  XNOR3X1 U8101 ( .IN1(n8018), .IN2(n8019), .IN3(n8021), .Q(n7994) );
  NAND2X0 U8102 ( .IN1(n8050), .IN2(n8051), .QN(n8021) );
  MUX21X1 U8103 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1484 ), .Q(n8051) );
  MUX21X1 U8104 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1485 ), .Q(n8050) );
  NAND2X0 U8105 ( .IN1(n8052), .IN2(n8053), .QN(n8019) );
  MUX21X1 U8106 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1489 ), .Q(n8053) );
  MUX21X1 U8107 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1488 ), .Q(n8052) );
  NAND2X0 U8108 ( .IN1(n8054), .IN2(n8055), .QN(n8018) );
  MUX21X1 U8109 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1486 ), .Q(n8055) );
  MUX21X1 U8110 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1487 ), .Q(n8054) );
  XOR2X1 U8111 ( .IN1(n7944), .IN2(n7943), .Q(n7982) );
  NAND2X0 U8112 ( .IN1(n8056), .IN2(n8057), .QN(n7943) );
  MUX21X1 U8113 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1481 ), .Q(n8057) );
  MUX21X1 U8114 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1480 ), .Q(n8056) );
  NAND2X0 U8115 ( .IN1(n8058), .IN2(n8059), .QN(n7944) );
  MUX21X1 U8116 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1483 ), .Q(n8059) );
  MUX21X1 U8117 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1482 ), .Q(n8058) );
  XOR2X1 U8118 ( .IN1(n7983), .IN2(n8060), .Q(n8039) );
  NAND2X0 U8119 ( .IN1(n7986), .IN2(n7987), .QN(n8060) );
  AO22X1 U8120 ( .IN1(n8061), .IN2(n8062), .IN3(n8063), .IN4(n8064), .Q(n7983)
         );
  OR2X1 U8121 ( .IN1(n8062), .IN2(n8061), .Q(n8063) );
  AO22X1 U8122 ( .IN1(n8065), .IN2(n8066), .IN3(n8067), .IN4(n6224), .Q(
        \i_m4stg_frac/a0cout[27] ) );
  AO22X1 U8123 ( .IN1(n8068), .IN2(n8069), .IN3(n8070), .IN4(n8071), .Q(n6224)
         );
  OR2X1 U8124 ( .IN1(n8068), .IN2(n8069), .Q(n8071) );
  AND2X1 U8125 ( .IN1(n8072), .IN2(n8073), .Q(n8070) );
  NAND2X0 U8126 ( .IN1(n6225), .IN2(n6223), .QN(n8067) );
  INVX0 U8127 ( .INP(n8065), .ZN(n6223) );
  INVX0 U8128 ( .INP(n6225), .ZN(n8066) );
  MUX21X1 U8129 ( .IN1(n8074), .IN2(n8075), .S(n8076), .Q(n6225) );
  INVX0 U8130 ( .INP(n8077), .ZN(n8076) );
  XOR2X1 U8131 ( .IN1(n8034), .IN2(n8032), .Q(n8065) );
  OA22X1 U8132 ( .IN1(n8078), .IN2(n8079), .IN3(n8080), .IN4(n8081), .Q(n8032)
         );
  AND2X1 U8133 ( .IN1(n8079), .IN2(n8078), .Q(n8081) );
  XNOR3X1 U8134 ( .IN1(n8082), .IN2(n8025), .IN3(n8031), .Q(n8034) );
  XOR3X1 U8135 ( .IN1(n8037), .IN2(n8036), .IN3(n8035), .Q(n8031) );
  XNOR3X1 U8136 ( .IN1(n8046), .IN2(n8047), .IN3(n8049), .Q(n8035) );
  NAND2X0 U8137 ( .IN1(n8083), .IN2(n8084), .QN(n8049) );
  MUX21X1 U8138 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1489 ), .Q(n8084) );
  MUX21X1 U8139 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1490 ), .Q(n8083) );
  NAND2X0 U8140 ( .IN1(n8085), .IN2(n8086), .QN(n8047) );
  MUX21X1 U8141 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1494 ), .Q(n8086) );
  MUX21X1 U8142 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1493 ), .Q(n8085) );
  NAND2X0 U8143 ( .IN1(n8087), .IN2(n8088), .QN(n8046) );
  MUX21X1 U8144 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1492 ), .Q(n8088) );
  MUX21X1 U8145 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1491 ), .Q(n8087) );
  AOI22X1 U8146 ( .IN1(n8089), .IN2(n8090), .IN3(n8091), .IN4(n8092), .QN(
        n8036) );
  OR2X1 U8147 ( .IN1(n8090), .IN2(n8089), .Q(n8091) );
  XNOR3X1 U8148 ( .IN1(n8061), .IN2(n8062), .IN3(n8064), .Q(n8037) );
  NAND2X0 U8149 ( .IN1(n8093), .IN2(n8094), .QN(n8064) );
  MUX21X1 U8150 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1483 ), .Q(n8094) );
  MUX21X1 U8151 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1484 ), .Q(n8093) );
  NAND2X0 U8152 ( .IN1(n8095), .IN2(n8096), .QN(n8062) );
  MUX21X1 U8153 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1488 ), .Q(n8096) );
  MUX21X1 U8154 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1487 ), .Q(n8095) );
  NAND2X0 U8155 ( .IN1(n8097), .IN2(n8098), .QN(n8061) );
  MUX21X1 U8156 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1485 ), .Q(n8098) );
  MUX21X1 U8157 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1486 ), .Q(n8097) );
  XOR2X1 U8158 ( .IN1(n7987), .IN2(n7986), .Q(n8025) );
  NAND2X0 U8159 ( .IN1(n8099), .IN2(n8100), .QN(n7986) );
  MUX21X1 U8160 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1480 ), .Q(n8100) );
  MUX21X1 U8161 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1479 ), .Q(n8099) );
  NAND2X0 U8162 ( .IN1(n8101), .IN2(n8102), .QN(n7987) );
  MUX21X1 U8163 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1482 ), .Q(n8102) );
  MUX21X1 U8164 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1481 ), .Q(n8101) );
  XOR2X1 U8165 ( .IN1(n8026), .IN2(n8103), .Q(n8082) );
  NAND2X0 U8166 ( .IN1(n8029), .IN2(n8030), .QN(n8103) );
  AO22X1 U8167 ( .IN1(n8104), .IN2(n8105), .IN3(n8106), .IN4(n8107), .Q(n8026)
         );
  OR2X1 U8168 ( .IN1(n8105), .IN2(n8104), .Q(n8106) );
  AO22X1 U8169 ( .IN1(n8108), .IN2(n8109), .IN3(n8110), .IN4(n6227), .Q(
        \i_m4stg_frac/a0cout[26] ) );
  AO22X1 U8170 ( .IN1(n8111), .IN2(n8112), .IN3(n8113), .IN4(n8114), .Q(n6227)
         );
  OR2X1 U8171 ( .IN1(n8111), .IN2(n8112), .Q(n8114) );
  AND2X1 U8172 ( .IN1(n8115), .IN2(n8116), .Q(n8113) );
  NAND2X0 U8173 ( .IN1(n6228), .IN2(n6226), .QN(n8110) );
  INVX0 U8174 ( .INP(n8108), .ZN(n6226) );
  INVX0 U8175 ( .INP(n6228), .ZN(n8109) );
  MUX21X1 U8176 ( .IN1(n8117), .IN2(n8118), .S(n8119), .Q(n6228) );
  INVX0 U8177 ( .INP(n8120), .ZN(n8119) );
  XOR2X1 U8178 ( .IN1(n8077), .IN2(n8075), .Q(n8108) );
  OA22X1 U8179 ( .IN1(n8121), .IN2(n8122), .IN3(n8123), .IN4(n8124), .Q(n8075)
         );
  AND2X1 U8180 ( .IN1(n8122), .IN2(n8121), .Q(n8124) );
  XNOR3X1 U8181 ( .IN1(n8125), .IN2(n8068), .IN3(n8074), .Q(n8077) );
  XOR3X1 U8182 ( .IN1(n8080), .IN2(n8079), .IN3(n8078), .Q(n8074) );
  XNOR3X1 U8183 ( .IN1(n8089), .IN2(n8090), .IN3(n8092), .Q(n8078) );
  NAND2X0 U8184 ( .IN1(n8126), .IN2(n8127), .QN(n8092) );
  MUX21X1 U8185 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1488 ), .Q(n8127) );
  MUX21X1 U8186 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1489 ), .Q(n8126) );
  NAND2X0 U8187 ( .IN1(n8128), .IN2(n8129), .QN(n8090) );
  MUX21X1 U8188 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1493 ), .Q(n8129) );
  MUX21X1 U8189 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1492 ), .Q(n8128) );
  NAND2X0 U8190 ( .IN1(n8130), .IN2(n8131), .QN(n8089) );
  MUX21X1 U8191 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1491 ), .Q(n8131) );
  MUX21X1 U8192 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1490 ), .Q(n8130) );
  AOI22X1 U8193 ( .IN1(n8132), .IN2(n8133), .IN3(n8134), .IN4(n8135), .QN(
        n8079) );
  OR2X1 U8194 ( .IN1(n8133), .IN2(n8132), .Q(n8134) );
  XNOR3X1 U8195 ( .IN1(n8104), .IN2(n8105), .IN3(n8107), .Q(n8080) );
  NAND2X0 U8196 ( .IN1(n8136), .IN2(n8137), .QN(n8107) );
  MUX21X1 U8197 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1482 ), .Q(n8137) );
  MUX21X1 U8198 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1483 ), .Q(n8136) );
  NAND2X0 U8199 ( .IN1(n8138), .IN2(n8139), .QN(n8105) );
  MUX21X1 U8200 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1487 ), .Q(n8139) );
  MUX21X1 U8201 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1486 ), .Q(n8138) );
  NAND2X0 U8202 ( .IN1(n8140), .IN2(n8141), .QN(n8104) );
  MUX21X1 U8203 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1484 ), .Q(n8141) );
  MUX21X1 U8204 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1485 ), .Q(n8140) );
  XOR2X1 U8205 ( .IN1(n8030), .IN2(n8029), .Q(n8068) );
  NAND2X0 U8206 ( .IN1(n8142), .IN2(n8143), .QN(n8029) );
  MUX21X1 U8207 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1479 ), .Q(n8143) );
  MUX21X1 U8208 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1478 ), .Q(n8142) );
  NAND2X0 U8209 ( .IN1(n8144), .IN2(n8145), .QN(n8030) );
  MUX21X1 U8210 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1481 ), .Q(n8145) );
  MUX21X1 U8211 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1480 ), .Q(n8144) );
  XOR2X1 U8212 ( .IN1(n8069), .IN2(n8146), .Q(n8125) );
  NAND2X0 U8213 ( .IN1(n8072), .IN2(n8073), .QN(n8146) );
  AO22X1 U8214 ( .IN1(n8147), .IN2(n8148), .IN3(n8149), .IN4(n8150), .Q(n8069)
         );
  OR2X1 U8215 ( .IN1(n8148), .IN2(n8147), .Q(n8149) );
  AO22X1 U8216 ( .IN1(n8151), .IN2(n8152), .IN3(n8153), .IN4(n6230), .Q(
        \i_m4stg_frac/a0cout[25] ) );
  AO22X1 U8217 ( .IN1(n8154), .IN2(n8155), .IN3(n8156), .IN4(n8157), .Q(n6230)
         );
  OR2X1 U8218 ( .IN1(n8154), .IN2(n8155), .Q(n8157) );
  AND2X1 U8219 ( .IN1(n8158), .IN2(n8159), .Q(n8156) );
  NAND2X0 U8220 ( .IN1(n6231), .IN2(n6229), .QN(n8153) );
  INVX0 U8221 ( .INP(n8151), .ZN(n6229) );
  INVX0 U8222 ( .INP(n6231), .ZN(n8152) );
  MUX21X1 U8223 ( .IN1(n8160), .IN2(n8161), .S(n8162), .Q(n6231) );
  INVX0 U8224 ( .INP(n8163), .ZN(n8162) );
  XOR2X1 U8225 ( .IN1(n8120), .IN2(n8118), .Q(n8151) );
  OA22X1 U8226 ( .IN1(n8164), .IN2(n8165), .IN3(n8166), .IN4(n8167), .Q(n8118)
         );
  AND2X1 U8227 ( .IN1(n8165), .IN2(n8164), .Q(n8167) );
  XNOR3X1 U8228 ( .IN1(n8168), .IN2(n8111), .IN3(n8117), .Q(n8120) );
  XOR3X1 U8229 ( .IN1(n8123), .IN2(n8122), .IN3(n8121), .Q(n8117) );
  XNOR3X1 U8230 ( .IN1(n8132), .IN2(n8133), .IN3(n8135), .Q(n8121) );
  NAND2X0 U8231 ( .IN1(n8169), .IN2(n8170), .QN(n8135) );
  MUX21X1 U8232 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1487 ), .Q(n8170) );
  MUX21X1 U8233 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1488 ), .Q(n8169) );
  NAND2X0 U8234 ( .IN1(n8171), .IN2(n8172), .QN(n8133) );
  MUX21X1 U8235 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1492 ), .Q(n8172) );
  MUX21X1 U8236 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1491 ), .Q(n8171) );
  NAND2X0 U8237 ( .IN1(n8173), .IN2(n8174), .QN(n8132) );
  MUX21X1 U8238 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1490 ), .Q(n8174) );
  MUX21X1 U8239 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1489 ), .Q(n8173) );
  AOI22X1 U8240 ( .IN1(n8175), .IN2(n8176), .IN3(n8177), .IN4(n8178), .QN(
        n8122) );
  OR2X1 U8241 ( .IN1(n8176), .IN2(n8175), .Q(n8177) );
  XNOR3X1 U8242 ( .IN1(n8147), .IN2(n8148), .IN3(n8150), .Q(n8123) );
  NAND2X0 U8243 ( .IN1(n8179), .IN2(n8180), .QN(n8150) );
  MUX21X1 U8244 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1481 ), .Q(n8180) );
  MUX21X1 U8245 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1482 ), .Q(n8179) );
  NAND2X0 U8246 ( .IN1(n8181), .IN2(n8182), .QN(n8148) );
  MUX21X1 U8247 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1486 ), .Q(n8182) );
  MUX21X1 U8248 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1485 ), .Q(n8181) );
  NAND2X0 U8249 ( .IN1(n8183), .IN2(n8184), .QN(n8147) );
  MUX21X1 U8250 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1483 ), .Q(n8184) );
  MUX21X1 U8251 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1484 ), .Q(n8183) );
  XOR2X1 U8252 ( .IN1(n8073), .IN2(n8072), .Q(n8111) );
  NAND2X0 U8253 ( .IN1(n8185), .IN2(n8186), .QN(n8072) );
  MUX21X1 U8254 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1478 ), .Q(n8186) );
  MUX21X1 U8255 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1477 ), .Q(n8185) );
  NAND2X0 U8256 ( .IN1(n8187), .IN2(n8188), .QN(n8073) );
  MUX21X1 U8257 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1480 ), .Q(n8188) );
  MUX21X1 U8258 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1479 ), .Q(n8187) );
  XOR2X1 U8259 ( .IN1(n8112), .IN2(n8189), .Q(n8168) );
  NAND2X0 U8260 ( .IN1(n8115), .IN2(n8116), .QN(n8189) );
  AO22X1 U8261 ( .IN1(n8190), .IN2(n8191), .IN3(n8192), .IN4(n8193), .Q(n8112)
         );
  OR2X1 U8262 ( .IN1(n8191), .IN2(n8190), .Q(n8192) );
  AO22X1 U8263 ( .IN1(n8194), .IN2(n8195), .IN3(n8196), .IN4(n6233), .Q(
        \i_m4stg_frac/a0cout[24] ) );
  AO22X1 U8264 ( .IN1(n8197), .IN2(n8198), .IN3(n8199), .IN4(n8200), .Q(n6233)
         );
  OR2X1 U8265 ( .IN1(n8197), .IN2(n8198), .Q(n8200) );
  AND2X1 U8266 ( .IN1(n8201), .IN2(n8202), .Q(n8199) );
  NAND2X0 U8267 ( .IN1(n6234), .IN2(n6232), .QN(n8196) );
  INVX0 U8268 ( .INP(n8194), .ZN(n6232) );
  INVX0 U8269 ( .INP(n6234), .ZN(n8195) );
  MUX21X1 U8270 ( .IN1(n8203), .IN2(n8204), .S(n8205), .Q(n6234) );
  INVX0 U8271 ( .INP(n8206), .ZN(n8205) );
  XOR2X1 U8272 ( .IN1(n8163), .IN2(n8161), .Q(n8194) );
  OA22X1 U8273 ( .IN1(n8207), .IN2(n8208), .IN3(n8209), .IN4(n8210), .Q(n8161)
         );
  AND2X1 U8274 ( .IN1(n8208), .IN2(n8207), .Q(n8210) );
  XNOR3X1 U8275 ( .IN1(n8211), .IN2(n8154), .IN3(n8160), .Q(n8163) );
  XOR3X1 U8276 ( .IN1(n8166), .IN2(n8165), .IN3(n8164), .Q(n8160) );
  XNOR3X1 U8277 ( .IN1(n8175), .IN2(n8176), .IN3(n8178), .Q(n8164) );
  NAND2X0 U8278 ( .IN1(n8212), .IN2(n8213), .QN(n8178) );
  MUX21X1 U8279 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1486 ), .Q(n8213) );
  MUX21X1 U8280 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1487 ), .Q(n8212) );
  NAND2X0 U8281 ( .IN1(n8214), .IN2(n8215), .QN(n8176) );
  MUX21X1 U8282 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1491 ), .Q(n8215) );
  MUX21X1 U8283 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1490 ), .Q(n8214) );
  NAND2X0 U8284 ( .IN1(n8216), .IN2(n8217), .QN(n8175) );
  MUX21X1 U8285 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1489 ), .Q(n8217) );
  MUX21X1 U8286 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1488 ), .Q(n8216) );
  AOI22X1 U8287 ( .IN1(n8218), .IN2(n8219), .IN3(n8220), .IN4(n8221), .QN(
        n8165) );
  OR2X1 U8288 ( .IN1(n8219), .IN2(n8218), .Q(n8220) );
  XNOR3X1 U8289 ( .IN1(n8190), .IN2(n8191), .IN3(n8193), .Q(n8166) );
  NAND2X0 U8290 ( .IN1(n8222), .IN2(n8223), .QN(n8193) );
  MUX21X1 U8291 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1480 ), .Q(n8223) );
  MUX21X1 U8292 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1481 ), .Q(n8222) );
  NAND2X0 U8293 ( .IN1(n8224), .IN2(n8225), .QN(n8191) );
  MUX21X1 U8294 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1485 ), .Q(n8225) );
  MUX21X1 U8295 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1484 ), .Q(n8224) );
  NAND2X0 U8296 ( .IN1(n8226), .IN2(n8227), .QN(n8190) );
  MUX21X1 U8297 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1482 ), .Q(n8227) );
  MUX21X1 U8298 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1483 ), .Q(n8226) );
  XOR2X1 U8299 ( .IN1(n8116), .IN2(n8115), .Q(n8154) );
  NAND2X0 U8300 ( .IN1(n8228), .IN2(n8229), .QN(n8115) );
  MUX21X1 U8301 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1477 ), .Q(n8229) );
  MUX21X1 U8302 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1476 ), .Q(n8228) );
  NAND2X0 U8303 ( .IN1(n8230), .IN2(n8231), .QN(n8116) );
  MUX21X1 U8304 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1479 ), .Q(n8231) );
  MUX21X1 U8305 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1478 ), .Q(n8230) );
  XOR2X1 U8306 ( .IN1(n8155), .IN2(n8232), .Q(n8211) );
  NAND2X0 U8307 ( .IN1(n8158), .IN2(n8159), .QN(n8232) );
  AO22X1 U8308 ( .IN1(n8233), .IN2(n8234), .IN3(n8235), .IN4(n8236), .Q(n8155)
         );
  OR2X1 U8309 ( .IN1(n8234), .IN2(n8233), .Q(n8235) );
  AO22X1 U8310 ( .IN1(n8237), .IN2(n8238), .IN3(n8239), .IN4(n6236), .Q(
        \i_m4stg_frac/a0cout[23] ) );
  AO22X1 U8311 ( .IN1(n8240), .IN2(n8241), .IN3(n8242), .IN4(n8243), .Q(n6236)
         );
  OR2X1 U8312 ( .IN1(n8240), .IN2(n8241), .Q(n8243) );
  AND2X1 U8313 ( .IN1(n8244), .IN2(n8245), .Q(n8242) );
  NAND2X0 U8314 ( .IN1(n6237), .IN2(n6235), .QN(n8239) );
  INVX0 U8315 ( .INP(n8237), .ZN(n6235) );
  INVX0 U8316 ( .INP(n6237), .ZN(n8238) );
  MUX21X1 U8317 ( .IN1(n8246), .IN2(n8247), .S(n8248), .Q(n6237) );
  INVX0 U8318 ( .INP(n8249), .ZN(n8248) );
  XOR2X1 U8319 ( .IN1(n8206), .IN2(n8204), .Q(n8237) );
  OA22X1 U8320 ( .IN1(n8250), .IN2(n8251), .IN3(n8252), .IN4(n8253), .Q(n8204)
         );
  AND2X1 U8321 ( .IN1(n8251), .IN2(n8250), .Q(n8253) );
  XNOR3X1 U8322 ( .IN1(n8254), .IN2(n8197), .IN3(n8203), .Q(n8206) );
  XOR3X1 U8323 ( .IN1(n8209), .IN2(n8208), .IN3(n8207), .Q(n8203) );
  XNOR3X1 U8324 ( .IN1(n8218), .IN2(n8219), .IN3(n8221), .Q(n8207) );
  NAND2X0 U8325 ( .IN1(n8255), .IN2(n8256), .QN(n8221) );
  MUX21X1 U8326 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1485 ), .Q(n8256) );
  MUX21X1 U8327 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1486 ), .Q(n8255) );
  NAND2X0 U8328 ( .IN1(n8257), .IN2(n8258), .QN(n8219) );
  MUX21X1 U8329 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1490 ), .Q(n8258) );
  MUX21X1 U8330 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1489 ), .Q(n8257) );
  NAND2X0 U8331 ( .IN1(n8259), .IN2(n8260), .QN(n8218) );
  MUX21X1 U8332 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1488 ), .Q(n8260) );
  MUX21X1 U8333 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1487 ), .Q(n8259) );
  AOI22X1 U8334 ( .IN1(n8261), .IN2(n8262), .IN3(n8263), .IN4(n8264), .QN(
        n8208) );
  OR2X1 U8335 ( .IN1(n8262), .IN2(n8261), .Q(n8263) );
  XNOR3X1 U8336 ( .IN1(n8233), .IN2(n8234), .IN3(n8236), .Q(n8209) );
  NAND2X0 U8337 ( .IN1(n8265), .IN2(n8266), .QN(n8236) );
  MUX21X1 U8338 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1479 ), .Q(n8266) );
  MUX21X1 U8339 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1480 ), .Q(n8265) );
  NAND2X0 U8340 ( .IN1(n8267), .IN2(n8268), .QN(n8234) );
  MUX21X1 U8341 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1484 ), .Q(n8268) );
  MUX21X1 U8342 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1483 ), .Q(n8267) );
  NAND2X0 U8343 ( .IN1(n8269), .IN2(n8270), .QN(n8233) );
  MUX21X1 U8344 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1481 ), .Q(n8270) );
  MUX21X1 U8345 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1482 ), .Q(n8269) );
  XOR2X1 U8346 ( .IN1(n8159), .IN2(n8158), .Q(n8197) );
  NAND2X0 U8347 ( .IN1(n8271), .IN2(n8272), .QN(n8158) );
  MUX21X1 U8348 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1475 ), .Q(n8272) );
  MUX21X1 U8349 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1476 ), .Q(n8271) );
  NAND2X0 U8350 ( .IN1(n8273), .IN2(n8274), .QN(n8159) );
  MUX21X1 U8351 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1478 ), .Q(n8274) );
  MUX21X1 U8352 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1477 ), .Q(n8273) );
  XOR2X1 U8353 ( .IN1(n8198), .IN2(n8275), .Q(n8254) );
  NAND2X0 U8354 ( .IN1(n8201), .IN2(n8202), .QN(n8275) );
  AO22X1 U8355 ( .IN1(n8276), .IN2(n8277), .IN3(n8278), .IN4(n8279), .Q(n8198)
         );
  OR2X1 U8356 ( .IN1(n8277), .IN2(n8276), .Q(n8278) );
  AO22X1 U8357 ( .IN1(n8280), .IN2(n8281), .IN3(n8282), .IN4(n6239), .Q(
        \i_m4stg_frac/a0cout[22] ) );
  AO22X1 U8358 ( .IN1(n8283), .IN2(n8284), .IN3(n8285), .IN4(n8286), .Q(n6239)
         );
  OR2X1 U8359 ( .IN1(n8283), .IN2(n8284), .Q(n8286) );
  AND2X1 U8360 ( .IN1(n8287), .IN2(n8288), .Q(n8285) );
  NAND2X0 U8361 ( .IN1(n6240), .IN2(n6238), .QN(n8282) );
  INVX0 U8362 ( .INP(n8280), .ZN(n6238) );
  INVX0 U8363 ( .INP(n6240), .ZN(n8281) );
  MUX21X1 U8364 ( .IN1(n8289), .IN2(n8290), .S(n8291), .Q(n6240) );
  INVX0 U8365 ( .INP(n8292), .ZN(n8291) );
  XOR2X1 U8366 ( .IN1(n8249), .IN2(n8247), .Q(n8280) );
  OA22X1 U8367 ( .IN1(n8293), .IN2(n8294), .IN3(n8295), .IN4(n8296), .Q(n8247)
         );
  AND2X1 U8368 ( .IN1(n8294), .IN2(n8293), .Q(n8296) );
  XNOR3X1 U8369 ( .IN1(n8297), .IN2(n8240), .IN3(n8246), .Q(n8249) );
  XOR3X1 U8370 ( .IN1(n8252), .IN2(n8251), .IN3(n8250), .Q(n8246) );
  XNOR3X1 U8371 ( .IN1(n8261), .IN2(n8262), .IN3(n8264), .Q(n8250) );
  NAND2X0 U8372 ( .IN1(n8298), .IN2(n8299), .QN(n8264) );
  MUX21X1 U8373 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1484 ), .Q(n8299) );
  MUX21X1 U8374 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1485 ), .Q(n8298) );
  NAND2X0 U8375 ( .IN1(n8300), .IN2(n8301), .QN(n8262) );
  MUX21X1 U8376 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1489 ), .Q(n8301) );
  MUX21X1 U8377 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1488 ), .Q(n8300) );
  NAND2X0 U8378 ( .IN1(n8302), .IN2(n8303), .QN(n8261) );
  MUX21X1 U8379 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1487 ), .Q(n8303) );
  MUX21X1 U8380 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1486 ), .Q(n8302) );
  AOI22X1 U8381 ( .IN1(n8304), .IN2(n8305), .IN3(n8306), .IN4(n8307), .QN(
        n8251) );
  OR2X1 U8382 ( .IN1(n8305), .IN2(n8304), .Q(n8306) );
  XNOR3X1 U8383 ( .IN1(n8276), .IN2(n8277), .IN3(n8279), .Q(n8252) );
  NAND2X0 U8384 ( .IN1(n8308), .IN2(n8309), .QN(n8279) );
  MUX21X1 U8385 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1478 ), .Q(n8309) );
  MUX21X1 U8386 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1479 ), .Q(n8308) );
  NAND2X0 U8387 ( .IN1(n8310), .IN2(n8311), .QN(n8277) );
  MUX21X1 U8388 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1483 ), .Q(n8311) );
  MUX21X1 U8389 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1482 ), .Q(n8310) );
  NAND2X0 U8390 ( .IN1(n8312), .IN2(n8313), .QN(n8276) );
  MUX21X1 U8391 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1480 ), .Q(n8313) );
  MUX21X1 U8392 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1481 ), .Q(n8312) );
  XOR2X1 U8393 ( .IN1(n8202), .IN2(n8201), .Q(n8240) );
  NAND2X0 U8394 ( .IN1(n8314), .IN2(n8315), .QN(n8201) );
  MUX21X1 U8395 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1475 ), .Q(n8315) );
  MUX21X1 U8396 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1474 ), .Q(n8314) );
  NAND2X0 U8397 ( .IN1(n8316), .IN2(n8317), .QN(n8202) );
  MUX21X1 U8398 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1477 ), .Q(n8317) );
  MUX21X1 U8399 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1476 ), .Q(n8316) );
  XOR2X1 U8400 ( .IN1(n8241), .IN2(n8318), .Q(n8297) );
  NAND2X0 U8401 ( .IN1(n8244), .IN2(n8245), .QN(n8318) );
  AO22X1 U8402 ( .IN1(n8319), .IN2(n8320), .IN3(n8321), .IN4(n8322), .Q(n8241)
         );
  OR2X1 U8403 ( .IN1(n8320), .IN2(n8319), .Q(n8321) );
  AO22X1 U8404 ( .IN1(n8323), .IN2(n8324), .IN3(n8325), .IN4(n6242), .Q(
        \i_m4stg_frac/a0cout[21] ) );
  AO22X1 U8405 ( .IN1(n8326), .IN2(n8327), .IN3(n8328), .IN4(n8329), .Q(n6242)
         );
  OR2X1 U8406 ( .IN1(n8326), .IN2(n8327), .Q(n8329) );
  AND2X1 U8407 ( .IN1(n8330), .IN2(n8331), .Q(n8328) );
  NAND2X0 U8408 ( .IN1(n6243), .IN2(n6241), .QN(n8325) );
  INVX0 U8409 ( .INP(n8323), .ZN(n6241) );
  INVX0 U8410 ( .INP(n6243), .ZN(n8324) );
  MUX21X1 U8411 ( .IN1(n8332), .IN2(n8333), .S(n8334), .Q(n6243) );
  INVX0 U8412 ( .INP(n8335), .ZN(n8334) );
  XOR2X1 U8413 ( .IN1(n8292), .IN2(n8290), .Q(n8323) );
  OA22X1 U8414 ( .IN1(n8336), .IN2(n8337), .IN3(n8338), .IN4(n8339), .Q(n8290)
         );
  AND2X1 U8415 ( .IN1(n8337), .IN2(n8336), .Q(n8339) );
  XNOR3X1 U8416 ( .IN1(n8340), .IN2(n8283), .IN3(n8289), .Q(n8292) );
  XOR3X1 U8417 ( .IN1(n8295), .IN2(n8294), .IN3(n8293), .Q(n8289) );
  XNOR3X1 U8418 ( .IN1(n8304), .IN2(n8305), .IN3(n8307), .Q(n8293) );
  NAND2X0 U8419 ( .IN1(n8341), .IN2(n8342), .QN(n8307) );
  MUX21X1 U8420 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1483 ), .Q(n8342) );
  MUX21X1 U8421 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1484 ), .Q(n8341) );
  NAND2X0 U8422 ( .IN1(n8343), .IN2(n8344), .QN(n8305) );
  MUX21X1 U8423 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1488 ), .Q(n8344) );
  MUX21X1 U8424 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1487 ), .Q(n8343) );
  NAND2X0 U8425 ( .IN1(n8345), .IN2(n8346), .QN(n8304) );
  MUX21X1 U8426 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1486 ), .Q(n8346) );
  MUX21X1 U8427 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1485 ), .Q(n8345) );
  AOI22X1 U8428 ( .IN1(n8347), .IN2(n8348), .IN3(n8349), .IN4(n8350), .QN(
        n8294) );
  OR2X1 U8429 ( .IN1(n8348), .IN2(n8347), .Q(n8349) );
  XNOR3X1 U8430 ( .IN1(n8319), .IN2(n8320), .IN3(n8322), .Q(n8295) );
  NAND2X0 U8431 ( .IN1(n8351), .IN2(n8352), .QN(n8322) );
  MUX21X1 U8432 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1477 ), .Q(n8352) );
  MUX21X1 U8433 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1478 ), .Q(n8351) );
  NAND2X0 U8434 ( .IN1(n8353), .IN2(n8354), .QN(n8320) );
  MUX21X1 U8435 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1482 ), .Q(n8354) );
  MUX21X1 U8436 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1481 ), .Q(n8353) );
  NAND2X0 U8437 ( .IN1(n8355), .IN2(n8356), .QN(n8319) );
  MUX21X1 U8438 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1479 ), .Q(n8356) );
  MUX21X1 U8439 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1480 ), .Q(n8355) );
  XOR2X1 U8440 ( .IN1(n8245), .IN2(n8244), .Q(n8283) );
  NAND2X0 U8441 ( .IN1(n8357), .IN2(n8358), .QN(n8244) );
  MUX21X1 U8442 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1473 ), .Q(n8358) );
  MUX21X1 U8443 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1474 ), .Q(n8357) );
  NAND2X0 U8444 ( .IN1(n8359), .IN2(n8360), .QN(n8245) );
  MUX21X1 U8445 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1475 ), .Q(n8360) );
  MUX21X1 U8446 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1476 ), .Q(n8359) );
  XOR2X1 U8447 ( .IN1(n8284), .IN2(n8361), .Q(n8340) );
  NAND2X0 U8448 ( .IN1(n8287), .IN2(n8288), .QN(n8361) );
  AO22X1 U8449 ( .IN1(n8362), .IN2(n8363), .IN3(n8364), .IN4(n8365), .Q(n8284)
         );
  OR2X1 U8450 ( .IN1(n8363), .IN2(n8362), .Q(n8364) );
  AO22X1 U8451 ( .IN1(n8366), .IN2(n8367), .IN3(n8368), .IN4(n6245), .Q(
        \i_m4stg_frac/a0cout[20] ) );
  AO22X1 U8452 ( .IN1(n8369), .IN2(n8370), .IN3(n8371), .IN4(n8372), .Q(n6245)
         );
  OR2X1 U8453 ( .IN1(n8369), .IN2(n8370), .Q(n8372) );
  AND2X1 U8454 ( .IN1(n8373), .IN2(n8374), .Q(n8371) );
  NAND2X0 U8455 ( .IN1(n6246), .IN2(n6244), .QN(n8368) );
  INVX0 U8456 ( .INP(n8366), .ZN(n6244) );
  INVX0 U8457 ( .INP(n6246), .ZN(n8367) );
  MUX21X1 U8458 ( .IN1(n8375), .IN2(n8376), .S(n8377), .Q(n6246) );
  INVX0 U8459 ( .INP(n8378), .ZN(n8377) );
  XOR2X1 U8460 ( .IN1(n8335), .IN2(n8333), .Q(n8366) );
  OA22X1 U8461 ( .IN1(n8379), .IN2(n8380), .IN3(n8381), .IN4(n8382), .Q(n8333)
         );
  AND2X1 U8462 ( .IN1(n8380), .IN2(n8379), .Q(n8382) );
  XNOR3X1 U8463 ( .IN1(n8383), .IN2(n8326), .IN3(n8332), .Q(n8335) );
  XOR3X1 U8464 ( .IN1(n8338), .IN2(n8337), .IN3(n8336), .Q(n8332) );
  XNOR3X1 U8465 ( .IN1(n8347), .IN2(n8348), .IN3(n8350), .Q(n8336) );
  NAND2X0 U8466 ( .IN1(n8384), .IN2(n8385), .QN(n8350) );
  MUX21X1 U8467 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1482 ), .Q(n8385) );
  MUX21X1 U8468 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1483 ), .Q(n8384) );
  NAND2X0 U8469 ( .IN1(n8386), .IN2(n8387), .QN(n8348) );
  MUX21X1 U8470 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1487 ), .Q(n8387) );
  MUX21X1 U8471 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1486 ), .Q(n8386) );
  NAND2X0 U8472 ( .IN1(n8388), .IN2(n8389), .QN(n8347) );
  MUX21X1 U8473 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1485 ), .Q(n8389) );
  MUX21X1 U8474 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1484 ), .Q(n8388) );
  AOI22X1 U8475 ( .IN1(n8390), .IN2(n8391), .IN3(n8392), .IN4(n8393), .QN(
        n8337) );
  OR2X1 U8476 ( .IN1(n8391), .IN2(n8390), .Q(n8392) );
  XNOR3X1 U8477 ( .IN1(n8362), .IN2(n8363), .IN3(n8365), .Q(n8338) );
  NAND2X0 U8478 ( .IN1(n8394), .IN2(n8395), .QN(n8365) );
  MUX21X1 U8479 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1476 ), .Q(n8395) );
  MUX21X1 U8480 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1477 ), .Q(n8394) );
  NAND2X0 U8481 ( .IN1(n8396), .IN2(n8397), .QN(n8363) );
  MUX21X1 U8482 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1481 ), .Q(n8397) );
  MUX21X1 U8483 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1480 ), .Q(n8396) );
  NAND2X0 U8484 ( .IN1(n8398), .IN2(n8399), .QN(n8362) );
  MUX21X1 U8485 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1478 ), .Q(n8399) );
  MUX21X1 U8486 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1479 ), .Q(n8398) );
  XOR2X1 U8487 ( .IN1(n8288), .IN2(n8287), .Q(n8326) );
  NAND2X0 U8488 ( .IN1(n8400), .IN2(n8401), .QN(n8287) );
  MUX21X1 U8489 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1473 ), .Q(n8401) );
  MUX21X1 U8490 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1472 ), .Q(n8400) );
  NAND2X0 U8491 ( .IN1(n8402), .IN2(n8403), .QN(n8288) );
  MUX21X1 U8492 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1475 ), .Q(n8403) );
  MUX21X1 U8493 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1474 ), .Q(n8402) );
  XOR2X1 U8494 ( .IN1(n8327), .IN2(n8404), .Q(n8383) );
  NAND2X0 U8495 ( .IN1(n8330), .IN2(n8331), .QN(n8404) );
  AO22X1 U8496 ( .IN1(n8405), .IN2(n8406), .IN3(n8407), .IN4(n8408), .Q(n8327)
         );
  OR2X1 U8497 ( .IN1(n8406), .IN2(n8405), .Q(n8407) );
  AO22X1 U8498 ( .IN1(n8409), .IN2(n8410), .IN3(n8411), .IN4(n6251), .Q(
        \i_m4stg_frac/a0cout[19] ) );
  AO22X1 U8499 ( .IN1(n8412), .IN2(n8413), .IN3(n8414), .IN4(n8415), .Q(n6251)
         );
  OR2X1 U8500 ( .IN1(n8412), .IN2(n8413), .Q(n8415) );
  AND2X1 U8501 ( .IN1(n8416), .IN2(n8417), .Q(n8414) );
  NAND2X0 U8502 ( .IN1(n6252), .IN2(n6250), .QN(n8411) );
  INVX0 U8503 ( .INP(n8409), .ZN(n6250) );
  INVX0 U8504 ( .INP(n6252), .ZN(n8410) );
  MUX21X1 U8505 ( .IN1(n8418), .IN2(n8419), .S(n8420), .Q(n6252) );
  INVX0 U8506 ( .INP(n8421), .ZN(n8420) );
  XOR2X1 U8507 ( .IN1(n8378), .IN2(n8376), .Q(n8409) );
  OA22X1 U8508 ( .IN1(n8422), .IN2(n8423), .IN3(n8424), .IN4(n8425), .Q(n8376)
         );
  AND2X1 U8509 ( .IN1(n8423), .IN2(n8422), .Q(n8425) );
  XNOR3X1 U8510 ( .IN1(n8426), .IN2(n8369), .IN3(n8375), .Q(n8378) );
  XOR3X1 U8511 ( .IN1(n8381), .IN2(n8380), .IN3(n8379), .Q(n8375) );
  XNOR3X1 U8512 ( .IN1(n8390), .IN2(n8391), .IN3(n8393), .Q(n8379) );
  NAND2X0 U8513 ( .IN1(n8427), .IN2(n8428), .QN(n8393) );
  MUX21X1 U8514 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1481 ), .Q(n8428) );
  MUX21X1 U8515 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1482 ), .Q(n8427) );
  NAND2X0 U8516 ( .IN1(n8429), .IN2(n8430), .QN(n8391) );
  MUX21X1 U8517 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1486 ), .Q(n8430) );
  MUX21X1 U8518 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1485 ), .Q(n8429) );
  NAND2X0 U8519 ( .IN1(n8431), .IN2(n8432), .QN(n8390) );
  MUX21X1 U8520 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1484 ), .Q(n8432) );
  MUX21X1 U8521 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1483 ), .Q(n8431) );
  AOI22X1 U8522 ( .IN1(n8433), .IN2(n8434), .IN3(n8435), .IN4(n8436), .QN(
        n8380) );
  OR2X1 U8523 ( .IN1(n8434), .IN2(n8433), .Q(n8435) );
  XNOR3X1 U8524 ( .IN1(n8405), .IN2(n8406), .IN3(n8408), .Q(n8381) );
  NAND2X0 U8525 ( .IN1(n8437), .IN2(n8438), .QN(n8408) );
  MUX21X1 U8526 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1475 ), .Q(n8438) );
  MUX21X1 U8527 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1476 ), .Q(n8437) );
  NAND2X0 U8528 ( .IN1(n8439), .IN2(n8440), .QN(n8406) );
  MUX21X1 U8529 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1480 ), .Q(n8440) );
  MUX21X1 U8530 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1479 ), .Q(n8439) );
  NAND2X0 U8531 ( .IN1(n8441), .IN2(n8442), .QN(n8405) );
  MUX21X1 U8532 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1477 ), .Q(n8442) );
  MUX21X1 U8533 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1478 ), .Q(n8441) );
  XOR2X1 U8534 ( .IN1(n8331), .IN2(n8330), .Q(n8369) );
  NAND2X0 U8535 ( .IN1(n8443), .IN2(n8444), .QN(n8330) );
  MUX21X1 U8536 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1472 ), .Q(n8444) );
  MUX21X1 U8537 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1471 ), .Q(n8443) );
  NAND2X0 U8538 ( .IN1(n8445), .IN2(n8446), .QN(n8331) );
  MUX21X1 U8539 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1473 ), .Q(n8446) );
  MUX21X1 U8540 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1474 ), .Q(n8445) );
  XOR2X1 U8541 ( .IN1(n8370), .IN2(n8447), .Q(n8426) );
  NAND2X0 U8542 ( .IN1(n8373), .IN2(n8374), .QN(n8447) );
  AO22X1 U8543 ( .IN1(n8448), .IN2(n8449), .IN3(n8450), .IN4(n8451), .Q(n8370)
         );
  OR2X1 U8544 ( .IN1(n8449), .IN2(n8448), .Q(n8450) );
  AO22X1 U8545 ( .IN1(n8452), .IN2(n8453), .IN3(n8454), .IN4(n6254), .Q(
        \i_m4stg_frac/a0cout[18] ) );
  AO22X1 U8546 ( .IN1(n8455), .IN2(n8456), .IN3(n8457), .IN4(n8458), .Q(n6254)
         );
  OR2X1 U8547 ( .IN1(n8455), .IN2(n8456), .Q(n8458) );
  AND2X1 U8548 ( .IN1(n8459), .IN2(n8460), .Q(n8457) );
  NAND2X0 U8549 ( .IN1(n6255), .IN2(n6253), .QN(n8454) );
  INVX0 U8550 ( .INP(n8452), .ZN(n6253) );
  INVX0 U8551 ( .INP(n6255), .ZN(n8453) );
  MUX21X1 U8552 ( .IN1(n8461), .IN2(n8462), .S(n8463), .Q(n6255) );
  INVX0 U8553 ( .INP(n8464), .ZN(n8463) );
  XOR2X1 U8554 ( .IN1(n8421), .IN2(n8419), .Q(n8452) );
  OA22X1 U8555 ( .IN1(n8465), .IN2(n8466), .IN3(n8467), .IN4(n8468), .Q(n8419)
         );
  AND2X1 U8556 ( .IN1(n8466), .IN2(n8465), .Q(n8468) );
  XNOR3X1 U8557 ( .IN1(n8469), .IN2(n8412), .IN3(n8418), .Q(n8421) );
  XOR3X1 U8558 ( .IN1(n8424), .IN2(n8423), .IN3(n8422), .Q(n8418) );
  XNOR3X1 U8559 ( .IN1(n8433), .IN2(n8434), .IN3(n8436), .Q(n8422) );
  NAND2X0 U8560 ( .IN1(n8470), .IN2(n8471), .QN(n8436) );
  MUX21X1 U8561 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1480 ), .Q(n8471) );
  MUX21X1 U8562 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1481 ), .Q(n8470) );
  NAND2X0 U8563 ( .IN1(n8472), .IN2(n8473), .QN(n8434) );
  MUX21X1 U8564 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1485 ), .Q(n8473) );
  MUX21X1 U8565 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1484 ), .Q(n8472) );
  NAND2X0 U8566 ( .IN1(n8474), .IN2(n8475), .QN(n8433) );
  MUX21X1 U8567 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1483 ), .Q(n8475) );
  MUX21X1 U8568 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1482 ), .Q(n8474) );
  AOI22X1 U8569 ( .IN1(n8476), .IN2(n8477), .IN3(n8478), .IN4(n8479), .QN(
        n8423) );
  OR2X1 U8570 ( .IN1(n8477), .IN2(n8476), .Q(n8478) );
  XNOR3X1 U8571 ( .IN1(n8448), .IN2(n8449), .IN3(n8451), .Q(n8424) );
  NAND2X0 U8572 ( .IN1(n8480), .IN2(n8481), .QN(n8451) );
  MUX21X1 U8573 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1474 ), .Q(n8481) );
  MUX21X1 U8574 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1475 ), .Q(n8480) );
  NAND2X0 U8575 ( .IN1(n8482), .IN2(n8483), .QN(n8449) );
  MUX21X1 U8576 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1479 ), .Q(n8483) );
  MUX21X1 U8577 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1478 ), .Q(n8482) );
  NAND2X0 U8578 ( .IN1(n8484), .IN2(n8485), .QN(n8448) );
  MUX21X1 U8579 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1476 ), .Q(n8485) );
  MUX21X1 U8580 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1477 ), .Q(n8484) );
  XOR2X1 U8581 ( .IN1(n8374), .IN2(n8373), .Q(n8412) );
  NAND2X0 U8582 ( .IN1(n8486), .IN2(n8487), .QN(n8373) );
  MUX21X1 U8583 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1471 ), .Q(n8487) );
  MUX21X1 U8584 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1470 ), .Q(n8486) );
  NAND2X0 U8585 ( .IN1(n8488), .IN2(n8489), .QN(n8374) );
  MUX21X1 U8586 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1473 ), .Q(n8489) );
  MUX21X1 U8587 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1472 ), .Q(n8488) );
  XOR2X1 U8588 ( .IN1(n8413), .IN2(n8490), .Q(n8469) );
  NAND2X0 U8589 ( .IN1(n8416), .IN2(n8417), .QN(n8490) );
  AO22X1 U8590 ( .IN1(n8491), .IN2(n8492), .IN3(n8493), .IN4(n8494), .Q(n8413)
         );
  OR2X1 U8591 ( .IN1(n8492), .IN2(n8491), .Q(n8493) );
  AO22X1 U8592 ( .IN1(n8495), .IN2(n8496), .IN3(n8497), .IN4(n6257), .Q(
        \i_m4stg_frac/a0cout[17] ) );
  AO22X1 U8593 ( .IN1(n8498), .IN2(n8499), .IN3(n8500), .IN4(n8501), .Q(n6257)
         );
  OR2X1 U8594 ( .IN1(n8498), .IN2(n8499), .Q(n8501) );
  NAND2X0 U8595 ( .IN1(n6258), .IN2(n6256), .QN(n8497) );
  INVX0 U8596 ( .INP(n8495), .ZN(n6256) );
  INVX0 U8597 ( .INP(n6258), .ZN(n8496) );
  MUX21X1 U8598 ( .IN1(n8502), .IN2(n8503), .S(n8504), .Q(n6258) );
  INVX0 U8599 ( .INP(n8505), .ZN(n8504) );
  XOR2X1 U8600 ( .IN1(n8464), .IN2(n8462), .Q(n8495) );
  OA22X1 U8601 ( .IN1(n8506), .IN2(n8507), .IN3(n8508), .IN4(n8509), .Q(n8462)
         );
  AND2X1 U8602 ( .IN1(n8507), .IN2(n8506), .Q(n8509) );
  XNOR3X1 U8603 ( .IN1(n8510), .IN2(n8455), .IN3(n8461), .Q(n8464) );
  XOR3X1 U8604 ( .IN1(n8467), .IN2(n8466), .IN3(n8465), .Q(n8461) );
  XNOR3X1 U8605 ( .IN1(n8476), .IN2(n8477), .IN3(n8479), .Q(n8465) );
  NAND2X0 U8606 ( .IN1(n8511), .IN2(n8512), .QN(n8479) );
  MUX21X1 U8607 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1479 ), .Q(n8512) );
  MUX21X1 U8608 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1480 ), .Q(n8511) );
  NAND2X0 U8609 ( .IN1(n8513), .IN2(n8514), .QN(n8477) );
  MUX21X1 U8610 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1484 ), .Q(n8514) );
  MUX21X1 U8611 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1483 ), .Q(n8513) );
  NAND2X0 U8612 ( .IN1(n8515), .IN2(n8516), .QN(n8476) );
  MUX21X1 U8613 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1482 ), .Q(n8516) );
  MUX21X1 U8614 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1481 ), .Q(n8515) );
  AOI22X1 U8615 ( .IN1(n8517), .IN2(n8518), .IN3(n8519), .IN4(n8520), .QN(
        n8466) );
  OR2X1 U8616 ( .IN1(n8518), .IN2(n8517), .Q(n8519) );
  XNOR3X1 U8617 ( .IN1(n8491), .IN2(n8492), .IN3(n8494), .Q(n8467) );
  NAND2X0 U8618 ( .IN1(n8521), .IN2(n8522), .QN(n8494) );
  MUX21X1 U8619 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1474 ), .Q(n8522) );
  MUX21X1 U8620 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1473 ), .Q(n8521) );
  NAND2X0 U8621 ( .IN1(n8523), .IN2(n8524), .QN(n8492) );
  MUX21X1 U8622 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1478 ), .Q(n8524) );
  MUX21X1 U8623 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1477 ), .Q(n8523) );
  NAND2X0 U8624 ( .IN1(n8525), .IN2(n8526), .QN(n8491) );
  MUX21X1 U8625 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1475 ), .Q(n8526) );
  MUX21X1 U8626 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1476 ), .Q(n8525) );
  XOR2X1 U8627 ( .IN1(n8417), .IN2(n8416), .Q(n8455) );
  NAND2X0 U8628 ( .IN1(n8527), .IN2(n8528), .QN(n8416) );
  MUX21X1 U8629 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1470 ), .Q(n8528) );
  MUX21X1 U8630 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1469 ), .Q(n8527) );
  NAND2X0 U8631 ( .IN1(n8529), .IN2(n8530), .QN(n8417) );
  MUX21X1 U8632 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1472 ), .Q(n8530) );
  MUX21X1 U8633 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1471 ), .Q(n8529) );
  XOR2X1 U8634 ( .IN1(n8456), .IN2(n8531), .Q(n8510) );
  NAND2X0 U8635 ( .IN1(n8459), .IN2(n8460), .QN(n8531) );
  AO22X1 U8636 ( .IN1(n8532), .IN2(n8533), .IN3(n8534), .IN4(n8535), .Q(n8456)
         );
  OR2X1 U8637 ( .IN1(n8533), .IN2(n8532), .Q(n8534) );
  AO22X1 U8638 ( .IN1(n6260), .IN2(n6261), .IN3(n8536), .IN4(n6259), .Q(
        \i_m4stg_frac/a0cout[16] ) );
  AO22X1 U8639 ( .IN1(n8537), .IN2(n8538), .IN3(n8539), .IN4(n8540), .Q(n6259)
         );
  OR2X1 U8640 ( .IN1(n8537), .IN2(n8538), .Q(n8540) );
  OR2X1 U8641 ( .IN1(n6261), .IN2(n6260), .Q(n8536) );
  INVX0 U8642 ( .INP(n8541), .ZN(n6261) );
  MUX21X1 U8643 ( .IN1(n8542), .IN2(n8543), .S(n8544), .Q(n8541) );
  INVX0 U8644 ( .INP(n8545), .ZN(n8544) );
  XNOR2X1 U8645 ( .IN1(n8505), .IN2(n8502), .Q(n6260) );
  OA22X1 U8646 ( .IN1(n8546), .IN2(n8547), .IN3(n8548), .IN4(n8549), .Q(n8502)
         );
  AND2X1 U8647 ( .IN1(n8547), .IN2(n8546), .Q(n8549) );
  XNOR3X1 U8648 ( .IN1(n8550), .IN2(n8500), .IN3(n8503), .Q(n8505) );
  XOR3X1 U8649 ( .IN1(n8508), .IN2(n8507), .IN3(n8506), .Q(n8503) );
  XNOR3X1 U8650 ( .IN1(n8517), .IN2(n8518), .IN3(n8520), .Q(n8506) );
  NAND2X0 U8651 ( .IN1(n8551), .IN2(n8552), .QN(n8520) );
  MUX21X1 U8652 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1478 ), .Q(n8552) );
  MUX21X1 U8653 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1479 ), .Q(n8551) );
  NAND2X0 U8654 ( .IN1(n8553), .IN2(n8554), .QN(n8518) );
  MUX21X1 U8655 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1483 ), .Q(n8554) );
  MUX21X1 U8656 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1482 ), .Q(n8553) );
  NAND2X0 U8657 ( .IN1(n8555), .IN2(n8556), .QN(n8517) );
  MUX21X1 U8658 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1481 ), .Q(n8556) );
  MUX21X1 U8659 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1480 ), .Q(n8555) );
  AOI22X1 U8660 ( .IN1(n8557), .IN2(n8558), .IN3(n8559), .IN4(n8560), .QN(
        n8507) );
  OR2X1 U8661 ( .IN1(n8558), .IN2(n8557), .Q(n8559) );
  XNOR3X1 U8662 ( .IN1(n8532), .IN2(n8533), .IN3(n8535), .Q(n8508) );
  NAND2X0 U8663 ( .IN1(n8561), .IN2(n8562), .QN(n8535) );
  MUX21X1 U8664 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1472 ), .Q(n8562) );
  MUX21X1 U8665 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1473 ), .Q(n8561) );
  NAND2X0 U8666 ( .IN1(n8563), .IN2(n8564), .QN(n8533) );
  MUX21X1 U8667 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1477 ), .Q(n8564) );
  MUX21X1 U8668 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1476 ), .Q(n8563) );
  NAND2X0 U8669 ( .IN1(n8565), .IN2(n8566), .QN(n8532) );
  MUX21X1 U8670 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1474 ), .Q(n8566) );
  MUX21X1 U8671 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1475 ), .Q(n8565) );
  XOR2X1 U8672 ( .IN1(n8459), .IN2(n8460), .Q(n8500) );
  NAND2X0 U8673 ( .IN1(n8567), .IN2(n8568), .QN(n8460) );
  MUX21X1 U8674 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1468 ), .Q(n8568) );
  MUX21X1 U8675 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1469 ), .Q(n8567) );
  NAND2X0 U8676 ( .IN1(n8569), .IN2(n8570), .QN(n8459) );
  MUX21X1 U8677 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1471 ), .Q(n8570) );
  MUX21X1 U8678 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1470 ), .Q(n8569) );
  XOR2X1 U8679 ( .IN1(n8499), .IN2(n8498), .Q(n8550) );
  AO22X1 U8680 ( .IN1(n8571), .IN2(n8572), .IN3(n8573), .IN4(n8574), .Q(n8498)
         );
  OR2X1 U8681 ( .IN1(n8571), .IN2(n8572), .Q(n8573) );
  AO22X1 U8682 ( .IN1(n8575), .IN2(n8576), .IN3(n8577), .IN4(n8578), .Q(n8499)
         );
  OR2X1 U8683 ( .IN1(n8576), .IN2(n8575), .Q(n8578) );
  AO22X1 U8684 ( .IN1(n8579), .IN2(n8580), .IN3(n8581), .IN4(n6263), .Q(
        \i_m4stg_frac/a0cout[15] ) );
  AO22X1 U8685 ( .IN1(n8582), .IN2(n8583), .IN3(n8584), .IN4(n8585), .Q(n6263)
         );
  OR2X1 U8686 ( .IN1(n8583), .IN2(n8582), .Q(n8585) );
  INVX0 U8687 ( .INP(n8586), .ZN(n8584) );
  NAND2X0 U8688 ( .IN1(n6264), .IN2(n6262), .QN(n8581) );
  INVX0 U8689 ( .INP(n8579), .ZN(n6262) );
  INVX0 U8690 ( .INP(n6264), .ZN(n8580) );
  MUX21X1 U8691 ( .IN1(n8587), .IN2(n8588), .S(n8589), .Q(n6264) );
  INVX0 U8692 ( .INP(n8590), .ZN(n8589) );
  INVX0 U8693 ( .INP(n8591), .ZN(n8587) );
  XOR2X1 U8694 ( .IN1(n8545), .IN2(n8543), .Q(n8579) );
  AOI22X1 U8695 ( .IN1(n8592), .IN2(n8593), .IN3(n8594), .IN4(n8595), .QN(
        n8543) );
  OR2X1 U8696 ( .IN1(n8593), .IN2(n8592), .Q(n8595) );
  XOR3X1 U8697 ( .IN1(n8596), .IN2(n8538), .IN3(n8542), .Q(n8545) );
  XOR3X1 U8698 ( .IN1(n8548), .IN2(n8547), .IN3(n8546), .Q(n8542) );
  XNOR3X1 U8699 ( .IN1(n8557), .IN2(n8558), .IN3(n8560), .Q(n8546) );
  NAND2X0 U8700 ( .IN1(n8597), .IN2(n8598), .QN(n8560) );
  MUX21X1 U8701 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1477 ), .Q(n8598) );
  MUX21X1 U8702 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1478 ), .Q(n8597) );
  NAND2X0 U8703 ( .IN1(n8599), .IN2(n8600), .QN(n8558) );
  MUX21X1 U8704 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1482 ), .Q(n8600) );
  MUX21X1 U8705 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1481 ), .Q(n8599) );
  NAND2X0 U8706 ( .IN1(n8601), .IN2(n8602), .QN(n8557) );
  MUX21X1 U8707 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1480 ), .Q(n8602) );
  MUX21X1 U8708 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1479 ), .Q(n8601) );
  AOI22X1 U8709 ( .IN1(n8603), .IN2(n8604), .IN3(n8605), .IN4(n8606), .QN(
        n8547) );
  OR2X1 U8710 ( .IN1(n8604), .IN2(n8603), .Q(n8605) );
  XNOR3X1 U8711 ( .IN1(n8571), .IN2(n8572), .IN3(n8574), .Q(n8548) );
  NAND2X0 U8712 ( .IN1(n8607), .IN2(n8608), .QN(n8574) );
  MUX21X1 U8713 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1472 ), .Q(n8608) );
  MUX21X1 U8714 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1471 ), .Q(n8607) );
  NAND2X0 U8715 ( .IN1(n8609), .IN2(n8610), .QN(n8572) );
  MUX21X1 U8716 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1476 ), .Q(n8610) );
  MUX21X1 U8717 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1475 ), .Q(n8609) );
  NAND2X0 U8718 ( .IN1(n8611), .IN2(n8612), .QN(n8571) );
  MUX21X1 U8719 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1474 ), .Q(n8612) );
  MUX21X1 U8720 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1473 ), .Q(n8611) );
  AO22X1 U8721 ( .IN1(n8613), .IN2(n8614), .IN3(n8615), .IN4(n8616), .Q(n8538)
         );
  OR2X1 U8722 ( .IN1(n8614), .IN2(n8613), .Q(n8615) );
  XOR2X1 U8723 ( .IN1(n8539), .IN2(n8537), .Q(n8596) );
  INVX0 U8724 ( .INP(n8617), .ZN(n8537) );
  MUX21X1 U8725 ( .IN1(n6353), .IN2(n8618), .S(\i_m4stg_frac/n1467 ), .Q(n8617) );
  NAND2X0 U8726 ( .IN1(n8619), .IN2(n8620), .QN(n8618) );
  XOR3X1 U8727 ( .IN1(n8575), .IN2(n8577), .IN3(n8576), .Q(n8539) );
  NAND2X0 U8728 ( .IN1(n8621), .IN2(n8622), .QN(n8576) );
  MUX21X1 U8729 ( .IN1(n6353), .IN2(n6493), .S(\i_m4stg_frac/n1468 ), .Q(n8622) );
  INVX0 U8730 ( .INP(n8623), .ZN(n8619) );
  OR2X1 U8731 ( .IN1(n8623), .IN2(\i_m4stg_frac/n998 ), .Q(n6353) );
  MUX21X1 U8732 ( .IN1(n6491), .IN2(n6492), .S(\i_m4stg_frac/n1467 ), .Q(n8621) );
  INVX0 U8733 ( .INP(n6491), .ZN(n8577) );
  NOR2X0 U8734 ( .IN1(\i_m4stg_frac/n999 ), .IN2(\i_m4stg_frac/n998 ), .QN(
        n6054) );
  NAND2X0 U8735 ( .IN1(n8624), .IN2(n8625), .QN(n8575) );
  MUX21X1 U8736 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1470 ), .Q(n8625) );
  MUX21X1 U8737 ( .IN1(n6566), .IN2(n6567), .S(\i_m4stg_frac/n1469 ), .Q(n8624) );
  AO22X1 U8738 ( .IN1(n8626), .IN2(n8627), .IN3(n8628), .IN4(n6266), .Q(
        \i_m4stg_frac/a0cout[14] ) );
  AO22X1 U8739 ( .IN1(n8629), .IN2(n8630), .IN3(n8631), .IN4(n8632), .Q(n6266)
         );
  OR2X1 U8740 ( .IN1(n8630), .IN2(n8629), .Q(n8632) );
  NAND2X0 U8741 ( .IN1(n6267), .IN2(n6265), .QN(n8628) );
  INVX0 U8742 ( .INP(n6267), .ZN(n8627) );
  MUX21X1 U8743 ( .IN1(n8633), .IN2(n8634), .S(n8635), .Q(n6267) );
  INVX0 U8744 ( .INP(n8636), .ZN(n8635) );
  INVX0 U8745 ( .INP(n6265), .ZN(n8626) );
  XNOR2X1 U8746 ( .IN1(n8590), .IN2(n8591), .Q(n6265) );
  XOR3X1 U8747 ( .IN1(n8637), .IN2(n8582), .IN3(n8588), .Q(n8590) );
  XNOR3X1 U8748 ( .IN1(n8593), .IN2(n8592), .IN3(n8594), .Q(n8588) );
  XOR3X1 U8749 ( .IN1(n8613), .IN2(n8614), .IN3(n8616), .Q(n8594) );
  NAND2X0 U8750 ( .IN1(n8638), .IN2(n8639), .QN(n8616) );
  MUX21X1 U8751 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1470 ), .Q(n8639) );
  MUX21X1 U8752 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1471 ), .Q(n8638) );
  NAND2X0 U8753 ( .IN1(n8640), .IN2(n8641), .QN(n8614) );
  MUX21X1 U8754 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1474 ), .Q(n8641) );
  MUX21X1 U8755 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1475 ), .Q(n8640) );
  NAND2X0 U8756 ( .IN1(n8642), .IN2(n8643), .QN(n8613) );
  MUX21X1 U8757 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1472 ), .Q(n8643) );
  MUX21X1 U8758 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1473 ), .Q(n8642) );
  XOR3X1 U8759 ( .IN1(n8603), .IN2(n8604), .IN3(n8606), .Q(n8592) );
  NAND2X0 U8760 ( .IN1(n8644), .IN2(n8645), .QN(n8606) );
  MUX21X1 U8761 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1476 ), .Q(n8645) );
  MUX21X1 U8762 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1477 ), .Q(n8644) );
  NAND2X0 U8763 ( .IN1(n8646), .IN2(n8647), .QN(n8604) );
  MUX21X1 U8764 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1481 ), .Q(n8647) );
  MUX21X1 U8765 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1480 ), .Q(n8646) );
  NAND2X0 U8766 ( .IN1(n8648), .IN2(n8649), .QN(n8603) );
  MUX21X1 U8767 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1479 ), .Q(n8649) );
  MUX21X1 U8768 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1478 ), .Q(n8648) );
  AO22X1 U8769 ( .IN1(n8650), .IN2(n8651), .IN3(n8652), .IN4(n8653), .Q(n8593)
         );
  OR2X1 U8770 ( .IN1(n8651), .IN2(n8650), .Q(n8652) );
  XOR2X1 U8771 ( .IN1(n8620), .IN2(n8654), .Q(n8582) );
  NOR2X0 U8772 ( .IN1(n1034), .IN2(n8623), .QN(n8654) );
  NAND2X0 U8773 ( .IN1(\i_m4stg_frac/n1000 ), .IN2(n976), .QN(n8623) );
  AO21X1 U8774 ( .IN1(n8655), .IN2(n6362), .IN3(n8656), .Q(n8620) );
  INVX0 U8775 ( .INP(n8657), .ZN(n8656) );
  MUX21X1 U8776 ( .IN1(n6361), .IN2(n6565), .S(\i_m4stg_frac/n1469 ), .Q(n8657) );
  XOR2X1 U8777 ( .IN1(n8586), .IN2(n8583), .Q(n8637) );
  AO22X1 U8778 ( .IN1(n8658), .IN2(n8659), .IN3(n8660), .IN4(n8661), .Q(n8583)
         );
  OR2X1 U8779 ( .IN1(n8659), .IN2(n8658), .Q(n8660) );
  AO22X1 U8780 ( .IN1(n6269), .IN2(n6270), .IN3(n8662), .IN4(n6268), .Q(
        \i_m4stg_frac/a0cout[13] ) );
  AO22X1 U8781 ( .IN1(n8663), .IN2(n8664), .IN3(n8665), .IN4(n6541), .Q(n6268)
         );
  OA21X1 U8782 ( .IN1(n8663), .IN2(n8664), .IN3(\i_m4stg_frac/n1467 ), .Q(
        n8665) );
  OR2X1 U8783 ( .IN1(n6270), .IN2(n6269), .Q(n8662) );
  INVX0 U8784 ( .INP(n8666), .ZN(n6270) );
  MUX21X1 U8785 ( .IN1(n8667), .IN2(n8668), .S(n8669), .Q(n8666) );
  INVX0 U8786 ( .INP(n8670), .ZN(n8669) );
  XOR2X1 U8787 ( .IN1(n8636), .IN2(n8634), .Q(n6269) );
  INVX0 U8788 ( .INP(n8671), .ZN(n8634) );
  XNOR3X1 U8789 ( .IN1(n8672), .IN2(n8629), .IN3(n8633), .Q(n8636) );
  AO21X1 U8790 ( .IN1(n8673), .IN2(n8674), .IN3(n8591), .Q(n8633) );
  NOR2X0 U8791 ( .IN1(n8674), .IN2(n8673), .QN(n8591) );
  XNOR3X1 U8792 ( .IN1(n8650), .IN2(n8651), .IN3(n8653), .Q(n8674) );
  NAND2X0 U8793 ( .IN1(n8675), .IN2(n8676), .QN(n8653) );
  MUX21X1 U8794 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1475 ), .Q(n8676) );
  MUX21X1 U8795 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1476 ), .Q(n8675) );
  NAND2X0 U8796 ( .IN1(n8677), .IN2(n8678), .QN(n8651) );
  MUX21X1 U8797 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1480 ), .Q(n8678) );
  MUX21X1 U8798 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1479 ), .Q(n8677) );
  NAND2X0 U8799 ( .IN1(n8679), .IN2(n8680), .QN(n8650) );
  MUX21X1 U8800 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1478 ), .Q(n8680) );
  MUX21X1 U8801 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1477 ), .Q(n8679) );
  AOI22X1 U8802 ( .IN1(n8681), .IN2(n8682), .IN3(n8683), .IN4(n8684), .QN(
        n8673) );
  OR2X1 U8803 ( .IN1(n8682), .IN2(n8681), .Q(n8683) );
  XOR3X1 U8804 ( .IN1(n8658), .IN2(n8659), .IN3(n8661), .Q(n8629) );
  NAND2X0 U8805 ( .IN1(n8685), .IN2(n8686), .QN(n8661) );
  MUX21X1 U8806 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1469 ), .Q(n8686) );
  MUX21X1 U8807 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1470 ), .Q(n8685) );
  NAND2X0 U8808 ( .IN1(n8687), .IN2(n8688), .QN(n8659) );
  MUX21X1 U8809 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1474 ), .Q(n8688) );
  MUX21X1 U8810 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1473 ), .Q(n8687) );
  NAND2X0 U8811 ( .IN1(n8689), .IN2(n8690), .QN(n8658) );
  MUX21X1 U8812 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1472 ), .Q(n8690) );
  MUX21X1 U8813 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1471 ), .Q(n8689) );
  XNOR2X1 U8814 ( .IN1(n8631), .IN2(n8630), .Q(n8672) );
  AO22X1 U8815 ( .IN1(n8691), .IN2(n8692), .IN3(n8693), .IN4(n8694), .Q(n8630)
         );
  OR2X1 U8816 ( .IN1(n8692), .IN2(n8691), .Q(n8693) );
  OA21X1 U8817 ( .IN1(n8695), .IN2(n8696), .IN3(n8586), .Q(n8631) );
  NAND3X0 U8818 ( .IN1(n8697), .IN2(n8695), .IN3(n6355), .QN(n8586) );
  AND2X1 U8819 ( .IN1(n6355), .IN2(n8697), .Q(n8696) );
  NAND2X0 U8820 ( .IN1(\i_m4stg_frac/n1003 ), .IN2(\i_m4stg_frac/n1467 ), .QN(
        n8697) );
  NOR2X0 U8821 ( .IN1(\i_m4stg_frac/n1001 ), .IN2(\i_m4stg_frac/n1002 ), .QN(
        n6355) );
  AO21X1 U8822 ( .IN1(n8655), .IN2(n6541), .IN3(n8698), .Q(n8695) );
  MUX21X1 U8823 ( .IN1(n6543), .IN2(n6544), .S(\i_m4stg_frac/n1467 ), .Q(n8698) );
  INVX0 U8824 ( .INP(n6567), .ZN(n6544) );
  INVX0 U8825 ( .INP(n6566), .ZN(n6543) );
  NOR2X0 U8826 ( .IN1(\i_m4stg_frac/n1002 ), .IN2(\i_m4stg_frac/n1003 ), .QN(
        n6362) );
  INVX0 U8827 ( .INP(n8699), .ZN(n6541) );
  XOR2X1 U8828 ( .IN1(n1038), .IN2(\i_m4stg_frac/n1468 ), .Q(n8655) );
  AO22X1 U8829 ( .IN1(n6272), .IN2(n6273), .IN3(n8700), .IN4(n6271), .Q(
        \i_m4stg_frac/a0cout[12] ) );
  AO22X1 U8830 ( .IN1(n8701), .IN2(n8702), .IN3(n8703), .IN4(n8704), .Q(n6271)
         );
  NAND2X0 U8831 ( .IN1(n8705), .IN2(n6597), .QN(n8704) );
  OR2X1 U8832 ( .IN1(n6273), .IN2(n6272), .Q(n8700) );
  INVX0 U8833 ( .INP(n8706), .ZN(n6273) );
  MUX21X1 U8834 ( .IN1(n8707), .IN2(n8708), .S(n8709), .Q(n8706) );
  INVX0 U8835 ( .INP(n8710), .ZN(n8709) );
  XOR2X1 U8836 ( .IN1(n8670), .IN2(n8668), .Q(n6272) );
  INVX0 U8837 ( .INP(n8711), .ZN(n8668) );
  XNOR3X1 U8838 ( .IN1(n8712), .IN2(n8664), .IN3(n8667), .Q(n8670) );
  AO21X1 U8839 ( .IN1(n8713), .IN2(n8714), .IN3(n8671), .Q(n8667) );
  NOR2X0 U8840 ( .IN1(n8714), .IN2(n8713), .QN(n8671) );
  XNOR3X1 U8841 ( .IN1(n8681), .IN2(n8682), .IN3(n8684), .Q(n8714) );
  NAND2X0 U8842 ( .IN1(n8715), .IN2(n8716), .QN(n8684) );
  MUX21X1 U8843 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1475 ), .Q(n8716) );
  MUX21X1 U8844 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1474 ), .Q(n8715) );
  NAND2X0 U8845 ( .IN1(n8717), .IN2(n8718), .QN(n8682) );
  MUX21X1 U8846 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1479 ), .Q(n8718) );
  MUX21X1 U8847 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1478 ), .Q(n8717) );
  NAND2X0 U8848 ( .IN1(n8719), .IN2(n8720), .QN(n8681) );
  MUX21X1 U8849 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1477 ), .Q(n8720) );
  MUX21X1 U8850 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1476 ), .Q(n8719) );
  AOI22X1 U8851 ( .IN1(n8721), .IN2(n8722), .IN3(n8723), .IN4(n8724), .QN(
        n8713) );
  OR2X1 U8852 ( .IN1(n8722), .IN2(n8721), .Q(n8723) );
  AO22X1 U8853 ( .IN1(n8725), .IN2(n8726), .IN3(n8727), .IN4(n8728), .Q(n8664)
         );
  OR2X1 U8854 ( .IN1(n8726), .IN2(n8725), .Q(n8727) );
  XNOR2X1 U8855 ( .IN1(n8729), .IN2(n8663), .Q(n8712) );
  XOR3X1 U8856 ( .IN1(n8691), .IN2(n8692), .IN3(n8694), .Q(n8663) );
  NAND2X0 U8857 ( .IN1(n8730), .IN2(n8731), .QN(n8694) );
  MUX21X1 U8858 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1468 ), .Q(n8731) );
  MUX21X1 U8859 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1469 ), .Q(n8730) );
  NAND2X0 U8860 ( .IN1(n8732), .IN2(n8733), .QN(n8692) );
  MUX21X1 U8861 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1472 ), .Q(n8733) );
  MUX21X1 U8862 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1473 ), .Q(n8732) );
  NAND2X0 U8863 ( .IN1(n8734), .IN2(n8735), .QN(n8691) );
  MUX21X1 U8864 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1470 ), .Q(n8735) );
  MUX21X1 U8865 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1471 ), .Q(n8734) );
  NOR2X0 U8866 ( .IN1(n1034), .IN2(n8699), .QN(n8729) );
  NAND2X0 U8867 ( .IN1(\i_m4stg_frac/n1003 ), .IN2(n1229), .QN(n8699) );
  NOR2X0 U8868 ( .IN1(n6274), .IN2(n6275), .QN(\i_m4stg_frac/a0cout[11] ) );
  OAI22X1 U8869 ( .IN1(n8736), .IN2(n8737), .IN3(n8738), .IN4(n8739), .QN(
        n6275) );
  AND2X1 U8870 ( .IN1(n8737), .IN2(n8736), .Q(n8739) );
  XOR2X1 U8871 ( .IN1(n8710), .IN2(n8707), .Q(n6274) );
  INVX0 U8872 ( .INP(n8740), .ZN(n8707) );
  XNOR3X1 U8873 ( .IN1(n8741), .IN2(n8703), .IN3(n8708), .Q(n8710) );
  AO21X1 U8874 ( .IN1(n8742), .IN2(n8743), .IN3(n8711), .Q(n8708) );
  NOR2X0 U8875 ( .IN1(n8743), .IN2(n8742), .QN(n8711) );
  XNOR3X1 U8876 ( .IN1(n8721), .IN2(n8722), .IN3(n8724), .Q(n8743) );
  NAND2X0 U8877 ( .IN1(n8744), .IN2(n8745), .QN(n8724) );
  MUX21X1 U8878 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1473 ), .Q(n8745) );
  MUX21X1 U8879 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1474 ), .Q(n8744) );
  NAND2X0 U8880 ( .IN1(n8746), .IN2(n8747), .QN(n8722) );
  MUX21X1 U8881 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1478 ), .Q(n8747) );
  MUX21X1 U8882 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1477 ), .Q(n8746) );
  NAND2X0 U8883 ( .IN1(n8748), .IN2(n8749), .QN(n8721) );
  MUX21X1 U8884 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1475 ), .Q(n8749) );
  MUX21X1 U8885 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1476 ), .Q(n8748) );
  AOI22X1 U8886 ( .IN1(n8750), .IN2(n8751), .IN3(n8752), .IN4(n8753), .QN(
        n8742) );
  OR2X1 U8887 ( .IN1(n8751), .IN2(n8750), .Q(n8752) );
  XOR3X1 U8888 ( .IN1(n8725), .IN2(n8726), .IN3(n8728), .Q(n8703) );
  NAND2X0 U8889 ( .IN1(n8754), .IN2(n8755), .QN(n8728) );
  MUX21X1 U8890 ( .IN1(n6597), .IN2(n6598), .S(\i_m4stg_frac/n1467 ), .Q(n8755) );
  MUX21X1 U8891 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1468 ), .Q(n8754) );
  NAND2X0 U8892 ( .IN1(n8756), .IN2(n8757), .QN(n8726) );
  MUX21X1 U8893 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1472 ), .Q(n8757) );
  MUX21X1 U8894 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1471 ), .Q(n8756) );
  NAND2X0 U8895 ( .IN1(n8758), .IN2(n8759), .QN(n8725) );
  MUX21X1 U8896 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1469 ), .Q(n8759) );
  MUX21X1 U8897 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1470 ), .Q(n8758) );
  XOR2X1 U8898 ( .IN1(n8702), .IN2(n8701), .Q(n8741) );
  INVX0 U8899 ( .INP(n8705), .ZN(n8701) );
  AO22X1 U8900 ( .IN1(n8760), .IN2(n8761), .IN3(n8762), .IN4(n8763), .Q(n8705)
         );
  OR2X1 U8901 ( .IN1(n8761), .IN2(n8760), .Q(n8763) );
  NOR2X0 U8902 ( .IN1(n6356), .IN2(\i_m4stg_frac/n1006 ), .QN(n8702) );
  AO22X1 U8903 ( .IN1(n6278), .IN2(n6277), .IN3(n6276), .IN4(n8764), .Q(
        \i_m4stg_frac/a0cout[10] ) );
  OR2X1 U8904 ( .IN1(n6278), .IN2(n6277), .Q(n8764) );
  AOI21X1 U8905 ( .IN1(n8765), .IN2(n8766), .IN3(n8740), .QN(n6276) );
  NOR2X0 U8906 ( .IN1(n8766), .IN2(n8765), .QN(n8740) );
  XNOR3X1 U8907 ( .IN1(n8750), .IN2(n8751), .IN3(n8753), .Q(n8766) );
  NAND2X0 U8908 ( .IN1(n8767), .IN2(n8768), .QN(n8753) );
  MUX21X1 U8909 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1472 ), .Q(n8768) );
  MUX21X1 U8910 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1473 ), .Q(n8767) );
  NAND2X0 U8911 ( .IN1(n8769), .IN2(n8770), .QN(n8751) );
  MUX21X1 U8912 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1477 ), .Q(n8770) );
  MUX21X1 U8913 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1476 ), .Q(n8769) );
  NAND2X0 U8914 ( .IN1(n8771), .IN2(n8772), .QN(n8750) );
  MUX21X1 U8915 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1475 ), .Q(n8772) );
  MUX21X1 U8916 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1474 ), .Q(n8771) );
  AOI22X1 U8917 ( .IN1(n8773), .IN2(n8774), .IN3(n8775), .IN4(n8776), .QN(
        n8765) );
  OR2X1 U8918 ( .IN1(n8773), .IN2(n8774), .Q(n8775) );
  AO22X1 U8919 ( .IN1(n8777), .IN2(n6284), .IN3(n8778), .IN4(n6283), .Q(n6277)
         );
  AO22X1 U8920 ( .IN1(n6304), .IN2(n6303), .IN3(n8779), .IN4(n6302), .Q(n6283)
         );
  NAND2X0 U8921 ( .IN1(n8780), .IN2(n8781), .QN(n6302) );
  MUX21X1 U8922 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1472 ), .Q(n8781) );
  MUX21X1 U8923 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1473 ), .Q(n8780) );
  OR2X1 U8924 ( .IN1(n6303), .IN2(n6304), .Q(n8779) );
  NAND2X0 U8925 ( .IN1(n8782), .IN2(n8783), .QN(n6303) );
  MUX21X1 U8926 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1475 ), .Q(n8783) );
  MUX21X1 U8927 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1474 ), .Q(n8782) );
  NAND2X0 U8928 ( .IN1(n8784), .IN2(n8785), .QN(n6304) );
  MUX21X1 U8929 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1470 ), .Q(n8785) );
  MUX21X1 U8930 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1471 ), .Q(n8784) );
  NAND2X0 U8931 ( .IN1(n8786), .IN2(n6285), .QN(n8778) );
  INVX0 U8932 ( .INP(n8777), .ZN(n6285) );
  INVX0 U8933 ( .INP(n8786), .ZN(n6284) );
  XOR3X1 U8934 ( .IN1(n6643), .IN2(n8787), .IN3(n8788), .Q(n8786) );
  XOR3X1 U8935 ( .IN1(n8776), .IN2(n8774), .IN3(n8773), .Q(n8777) );
  NAND2X0 U8936 ( .IN1(n8789), .IN2(n8790), .QN(n8773) );
  MUX21X1 U8937 ( .IN1(n6326), .IN2(n6327), .S(\i_m4stg_frac/n1472 ), .Q(n8790) );
  NOR2X0 U8938 ( .IN1(n950), .IN2(n6413), .QN(n6694) );
  MUX21X1 U8939 ( .IN1(n6324), .IN2(n6325), .S(\i_m4stg_frac/n1471 ), .Q(n8789) );
  NOR2X0 U8940 ( .IN1(n6413), .IN2(\i_m4stg_frac/n1015 ), .QN(n6434) );
  NAND2X0 U8941 ( .IN1(n1144), .IN2(n935), .QN(n6413) );
  NAND2X0 U8942 ( .IN1(n8791), .IN2(n8792), .QN(n8774) );
  MUX21X1 U8943 ( .IN1(n6332), .IN2(n6333), .S(\i_m4stg_frac/n1475 ), .Q(n8792) );
  NOR2X0 U8944 ( .IN1(\i_m4stg_frac/n1020 ), .IN2(\i_m4stg_frac/n1021 ), .QN(
        n6569) );
  MUX21X1 U8945 ( .IN1(n6330), .IN2(n6331), .S(\i_m4stg_frac/n1476 ), .Q(n8791) );
  OR2X1 U8946 ( .IN1(n1053), .IN2(n6279), .Q(n6331) );
  NOR2X0 U8947 ( .IN1(n6279), .IN2(\i_m4stg_frac/n1019 ), .QN(n6570) );
  NAND2X0 U8948 ( .IN1(\i_m4stg_frac/n1021 ), .IN2(n1327), .QN(n6279) );
  NAND2X0 U8949 ( .IN1(n8793), .IN2(n8794), .QN(n8776) );
  MUX21X1 U8950 ( .IN1(n6336), .IN2(n6337), .S(\i_m4stg_frac/n1474 ), .Q(n8794) );
  NOR2X0 U8951 ( .IN1(n1135), .IN2(n6466), .QN(n7109) );
  MUX21X1 U8952 ( .IN1(n6338), .IN2(n6339), .S(\i_m4stg_frac/n1473 ), .Q(n8793) );
  NOR2X0 U8953 ( .IN1(n6466), .IN2(\i_m4stg_frac/n1018 ), .QN(n7100) );
  OR2X1 U8954 ( .IN1(\i_m4stg_frac/n1017 ), .IN2(\i_m4stg_frac/n1016 ), .Q(
        n6466) );
  XNOR3X1 U8955 ( .IN1(n6621), .IN2(n8736), .IN3(n8738), .Q(n6278) );
  XNOR3X1 U8956 ( .IN1(n8761), .IN2(n8760), .IN3(n8762), .Q(n8738) );
  AND2X1 U8957 ( .IN1(n8795), .IN2(n8796), .Q(n8762) );
  MUX21X1 U8958 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1468 ), .Q(n8796) );
  MUX21X1 U8959 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1469 ), .Q(n8795) );
  AND2X1 U8960 ( .IN1(n8797), .IN2(n8798), .Q(n8760) );
  MUX21X1 U8961 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1471 ), .Q(n8798) );
  MUX21X1 U8962 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1470 ), .Q(n8797) );
  MUX21X1 U8963 ( .IN1(n6621), .IN2(n6622), .S(\i_m4stg_frac/n1467 ), .Q(n8761) );
  AO22X1 U8964 ( .IN1(n8788), .IN2(n8787), .IN3(n8799), .IN4(n8800), .Q(n8736)
         );
  OR2X1 U8965 ( .IN1(n8788), .IN2(n8787), .Q(n8800) );
  INVX0 U8966 ( .INP(n6643), .ZN(n8799) );
  NAND2X0 U8967 ( .IN1(n8801), .IN2(n8802), .QN(n8787) );
  MUX21X1 U8968 ( .IN1(n6643), .IN2(n6644), .S(\i_m4stg_frac/n1467 ), .Q(n8802) );
  MUX21X1 U8969 ( .IN1(n6395), .IN2(n6294), .S(\i_m4stg_frac/n1468 ), .Q(n8801) );
  NOR2X0 U8970 ( .IN1(\i_m4stg_frac/n1007 ), .IN2(\i_m4stg_frac/n1008 ), .QN(
        n6377) );
  NAND2X0 U8971 ( .IN1(n8803), .IN2(n8804), .QN(n8788) );
  MUX21X1 U8972 ( .IN1(n6314), .IN2(n6315), .S(\i_m4stg_frac/n1470 ), .Q(n8804) );
  AND2X1 U8973 ( .IN1(\i_m4stg_frac/n1012 ), .IN2(n1169), .Q(n6351) );
  INVX0 U8974 ( .INP(n6399), .ZN(n6347) );
  NAND2X0 U8975 ( .IN1(n1169), .IN2(n913), .QN(n6399) );
  MUX21X1 U8976 ( .IN1(n6312), .IN2(n6313), .S(\i_m4stg_frac/n1469 ), .Q(n8803) );
  NOR2X0 U8977 ( .IN1(\i_m4stg_frac/n1011 ), .IN2(\i_m4stg_frac/n1012 ), .QN(
        n6418) );
  NOR2X0 U8978 ( .IN1(n951), .IN2(n6356), .QN(n8737) );
  NAND2X0 U8979 ( .IN1(n1145), .IN2(n936), .QN(n6356) );
  AO22X1 U8980 ( .IN1(inq_in2[43]), .IN2(n1603), .IN3(n1391), .IN4(n917), .Q(
        \fpu_mul_frac_dp/n999 ) );
  AO22X1 U8981 ( .IN1(inq_in2[44]), .IN2(n1603), .IN3(n1391), .IN4(n880), .Q(
        \fpu_mul_frac_dp/n998 ) );
  AO22X1 U8982 ( .IN1(inq_in2[45]), .IN2(n1603), .IN3(n1391), .IN4(n1044), .Q(
        \fpu_mul_frac_dp/n997 ) );
  AO22X1 U8983 ( .IN1(inq_in2[46]), .IN2(n1603), .IN3(n1391), .IN4(n918), .Q(
        \fpu_mul_frac_dp/n996 ) );
  AO22X1 U8984 ( .IN1(inq_in2[47]), .IN2(n1603), .IN3(n1391), .IN4(n890), .Q(
        \fpu_mul_frac_dp/n995 ) );
  AO22X1 U8985 ( .IN1(inq_in2[48]), .IN2(n1603), .IN3(n1391), .IN4(n1042), .Q(
        \fpu_mul_frac_dp/n994 ) );
  AO22X1 U8986 ( .IN1(inq_in2[49]), .IN2(n1603), .IN3(n1391), .IN4(n891), .Q(
        \fpu_mul_frac_dp/n993 ) );
  AO22X1 U8987 ( .IN1(inq_in2[50]), .IN2(n1603), .IN3(n1391), .IN4(n916), .Q(
        \fpu_mul_frac_dp/n992 ) );
  AO22X1 U8988 ( .IN1(inq_in2[51]), .IN2(n1604), .IN3(n1391), .IN4(n1132), .Q(
        \fpu_mul_frac_dp/n991 ) );
  AO22X1 U8989 ( .IN1(inq_in2[52]), .IN2(n1604), .IN3(n1390), .IN4(n942), .Q(
        \fpu_mul_frac_dp/n990 ) );
  AO22X1 U8990 ( .IN1(inq_in2[53]), .IN2(n1604), .IN3(n1390), .IN4(n1151), .Q(
        \fpu_mul_frac_dp/n989 ) );
  AO21X1 U8991 ( .IN1(n1386), .IN2(n1224), .IN3(n1632), .Q(
        \fpu_mul_frac_dp/n988 ) );
  AO22X1 U8992 ( .IN1(m3bstg_ld0_inv[0]), .IN2(n1604), .IN3(m3stg_ld0_inv[0]), 
        .IN4(n1384), .Q(\fpu_mul_frac_dp/n987 ) );
  AO22X1 U8993 ( .IN1(m3bstg_ld0_inv[1]), .IN2(n1604), .IN3(m3stg_ld0_inv[1]), 
        .IN4(n1384), .Q(\fpu_mul_frac_dp/n986 ) );
  AO22X1 U8994 ( .IN1(m3bstg_ld0_inv[2]), .IN2(n1604), .IN3(m3stg_ld0_inv[2]), 
        .IN4(n1384), .Q(\fpu_mul_frac_dp/n985 ) );
  AO22X1 U8995 ( .IN1(m3bstg_ld0_inv[3]), .IN2(n1604), .IN3(m3stg_ld0_inv[3]), 
        .IN4(n1384), .Q(\fpu_mul_frac_dp/n984 ) );
  AO22X1 U8996 ( .IN1(m3bstg_ld0_inv[4]), .IN2(n1604), .IN3(m3stg_ld0_inv[4]), 
        .IN4(n1384), .Q(\fpu_mul_frac_dp/n983 ) );
  AO22X1 U8997 ( .IN1(m3bstg_ld0_inv[5]), .IN2(n1604), .IN3(m3stg_ld0_inv[5]), 
        .IN4(n1383), .Q(\fpu_mul_frac_dp/n982 ) );
  AO22X1 U8998 ( .IN1(m3bstg_ld0_inv[6]), .IN2(n1604), .IN3(m3stg_ld0_inv[6]), 
        .IN4(n1384), .Q(\fpu_mul_frac_dp/n981 ) );
  AO222X1 U8999 ( .IN1(n8805), .IN2(n1340), .IN3(n1592), .IN4(n8806), .IN5(
        n1383), .IN6(n884), .Q(\fpu_mul_frac_dp/n980 ) );
  OAI21X1 U9000 ( .IN1(n895), .IN2(n8807), .IN3(n8808), .QN(n8806) );
  AO222X1 U9001 ( .IN1(n8805), .IN2(n1051), .IN3(n1592), .IN4(n8809), .IN5(
        n1383), .IN6(n879), .Q(\fpu_mul_frac_dp/n979 ) );
  NAND2X0 U9002 ( .IN1(n8810), .IN2(n8811), .QN(n8809) );
  NAND3X0 U9003 ( .IN1(n1115), .IN2(n895), .IN3(n8812), .QN(n8811) );
  AO222X1 U9004 ( .IN1(n8805), .IN2(n1150), .IN3(n8813), .IN4(n1592), .IN5(
        n1383), .IN6(n906), .Q(\fpu_mul_frac_dp/n978 ) );
  MUX21X1 U9005 ( .IN1(n8814), .IN2(n8815), .S(n106), .Q(n8813) );
  INVX0 U9006 ( .INP(n8810), .ZN(n8815) );
  OA22X1 U9007 ( .IN1(n8816), .IN2(n8817), .IN3(n8818), .IN4(n8819), .Q(n8810)
         );
  OR2X1 U9008 ( .IN1(n452), .IN2(n8820), .Q(n8818) );
  AO22X1 U9009 ( .IN1(n8812), .IN2(n8817), .IN3(n8821), .IN4(n8822), .Q(n8814)
         );
  NOR2X0 U9010 ( .IN1(n1115), .IN2(n8820), .QN(n8821) );
  AO22X1 U9011 ( .IN1(n1595), .IN2(n8823), .IN3(n1387), .IN4(n1033), .Q(
        \fpu_mul_frac_dp/n977 ) );
  NAND4X0 U9012 ( .IN1(n8824), .IN2(n8825), .IN3(n8826), .IN4(n8808), .QN(
        n8823) );
  NAND2X0 U9013 ( .IN1(n8812), .IN2(n8827), .QN(n8826) );
  NAND2X0 U9014 ( .IN1(n8807), .IN2(n1280), .QN(n8825) );
  MUX21X1 U9015 ( .IN1(n8828), .IN2(n8829), .S(n110), .Q(n8824) );
  NAND2X0 U9016 ( .IN1(n8822), .IN2(n8830), .QN(n8829) );
  OA22X1 U9017 ( .IN1(n8831), .IN2(n8816), .IN3(n8830), .IN4(n8819), .Q(n8828)
         );
  NOR2X0 U9018 ( .IN1(n1166), .IN2(n8817), .QN(n8831) );
  NAND2X0 U9019 ( .IN1(n98), .IN2(n452), .QN(n8817) );
  AO222X1 U9020 ( .IN1(n8805), .IN2(n1059), .IN3(n1592), .IN4(n8832), .IN5(
        n1383), .IN6(n908), .Q(\fpu_mul_frac_dp/n976 ) );
  NAND3X0 U9021 ( .IN1(n8808), .IN2(n8833), .IN3(n8834), .QN(n8832) );
  MUX21X1 U9022 ( .IN1(n8835), .IN2(n8836), .S(n888), .Q(n8834) );
  OA22X1 U9023 ( .IN1(n8827), .IN2(n8816), .IN3(n8837), .IN4(n8819), .Q(n8836)
         );
  NAND2X0 U9024 ( .IN1(n8822), .IN2(n8837), .QN(n8835) );
  INVX0 U9025 ( .INP(n8819), .ZN(n8822) );
  NOR2X0 U9026 ( .IN1(n8838), .IN2(n1723), .QN(n8805) );
  AO22X1 U9027 ( .IN1(n1594), .IN2(n8839), .IN3(n1387), .IN4(n1036), .Q(
        \fpu_mul_frac_dp/n975 ) );
  AO22X1 U9028 ( .IN1(n1595), .IN2(n8839), .IN3(n1387), .IN4(n1035), .Q(
        \fpu_mul_frac_dp/n974 ) );
  NAND3X0 U9029 ( .IN1(n8840), .IN2(n8808), .IN3(n8841), .QN(n8839) );
  MUX21X1 U9030 ( .IN1(n8842), .IN2(n8843), .S(n118), .Q(n8841) );
  OA21X1 U9031 ( .IN1(n8844), .IN2(n8819), .IN3(n8833), .Q(n8843) );
  NAND2X0 U9032 ( .IN1(n8812), .IN2(n8845), .QN(n8833) );
  OA22X1 U9033 ( .IN1(n8845), .IN2(n8816), .IN3(n8819), .IN4(n8846), .Q(n8842)
         );
  INVX0 U9034 ( .INP(n8844), .ZN(n8846) );
  NOR2X0 U9035 ( .IN1(n8837), .IN2(n888), .QN(n8844) );
  INVX0 U9036 ( .INP(n8812), .ZN(n8816) );
  NOR2X0 U9037 ( .IN1(n8847), .IN2(n8807), .QN(n8812) );
  NAND3X0 U9038 ( .IN1(n8838), .IN2(n1119), .IN3(n8820), .QN(n8808) );
  NAND4X0 U9039 ( .IN1(n1114), .IN2(n900), .IN3(n8848), .IN4(n8849), .QN(n8820) );
  NOR4X0 U9040 ( .IN1(n142), .IN2(n138), .IN3(n134), .IN4(n130), .QN(n8849) );
  NAND3X0 U9041 ( .IN1(n114), .IN2(n110), .IN3(n118), .QN(n8848) );
  NAND2X0 U9042 ( .IN1(n8807), .IN2(n1279), .QN(n8840) );
  INVX0 U9043 ( .INP(n8838), .ZN(n8807) );
  NAND3X0 U9044 ( .IN1(n8850), .IN2(n8851), .IN3(n8852), .QN(
        \fpu_mul_frac_dp/n973 ) );
  MUX21X1 U9045 ( .IN1(n8853), .IN2(n8854), .S(n8855), .Q(n8852) );
  NAND2X0 U9046 ( .IN1(n8856), .IN2(m5stg_fmulda), .QN(n8854) );
  NAND2X0 U9047 ( .IN1(mul_frac_out[0]), .IN2(n1407), .QN(n8850) );
  NAND3X0 U9048 ( .IN1(n8857), .IN2(n8851), .IN3(n8858), .QN(
        \fpu_mul_frac_dp/n972 ) );
  MUX21X1 U9049 ( .IN1(n8859), .IN2(n8860), .S(n8861), .Q(n8858) );
  NAND2X0 U9050 ( .IN1(mul_frac_out[1]), .IN2(n1407), .QN(n8857) );
  NAND3X0 U9051 ( .IN1(n8862), .IN2(n8851), .IN3(n8863), .QN(
        \fpu_mul_frac_dp/n971 ) );
  MUX21X1 U9052 ( .IN1(n8864), .IN2(n8865), .S(n8866), .Q(n8863) );
  OR2X1 U9053 ( .IN1(n8860), .IN2(n8861), .Q(n8864) );
  NAND3X0 U9054 ( .IN1(m5stg_fmulda), .IN2(n8867), .IN3(n8856), .QN(n8860) );
  NAND2X0 U9055 ( .IN1(mul_frac_out[2]), .IN2(n1408), .QN(n8862) );
  NAND3X0 U9056 ( .IN1(n8868), .IN2(n8851), .IN3(n8869), .QN(
        \fpu_mul_frac_dp/n970 ) );
  MUX21X1 U9057 ( .IN1(n8870), .IN2(n8871), .S(n8872), .Q(n8869) );
  NAND2X0 U9058 ( .IN1(n8856), .IN2(n8873), .QN(n8871) );
  NAND2X0 U9059 ( .IN1(mul_frac_out[3]), .IN2(n1407), .QN(n8868) );
  NAND3X0 U9060 ( .IN1(n8874), .IN2(n8851), .IN3(n8875), .QN(
        \fpu_mul_frac_dp/n969 ) );
  MUX21X1 U9061 ( .IN1(n8876), .IN2(n8877), .S(n8878), .Q(n8875) );
  NAND3X0 U9062 ( .IN1(n8873), .IN2(n8879), .IN3(n8856), .QN(n8877) );
  NAND2X0 U9063 ( .IN1(mul_frac_out[4]), .IN2(n1407), .QN(n8874) );
  NAND3X0 U9064 ( .IN1(n8880), .IN2(n8851), .IN3(n8881), .QN(
        \fpu_mul_frac_dp/n968 ) );
  MUX21X1 U9065 ( .IN1(n8882), .IN2(n8883), .S(n8884), .Q(n8881) );
  NAND2X0 U9066 ( .IN1(n8856), .IN2(n8885), .QN(n8883) );
  NAND2X0 U9067 ( .IN1(mul_frac_out[5]), .IN2(n1407), .QN(n8880) );
  NAND3X0 U9068 ( .IN1(n8886), .IN2(n8851), .IN3(n8887), .QN(
        \fpu_mul_frac_dp/n967 ) );
  MUX21X1 U9069 ( .IN1(n8888), .IN2(n8889), .S(n8890), .Q(n8887) );
  NAND3X0 U9070 ( .IN1(n8885), .IN2(n8891), .IN3(n8856), .QN(n8889) );
  NAND2X0 U9071 ( .IN1(mul_frac_out[6]), .IN2(n1407), .QN(n8886) );
  NAND3X0 U9072 ( .IN1(n8892), .IN2(n8851), .IN3(n8893), .QN(
        \fpu_mul_frac_dp/n966 ) );
  MUX21X1 U9073 ( .IN1(n8894), .IN2(n8895), .S(n8896), .Q(n8893) );
  NAND2X0 U9074 ( .IN1(n8856), .IN2(n8897), .QN(n8895) );
  NAND2X0 U9075 ( .IN1(mul_frac_out[7]), .IN2(n1407), .QN(n8892) );
  NAND3X0 U9076 ( .IN1(n8898), .IN2(n8851), .IN3(n8899), .QN(
        \fpu_mul_frac_dp/n965 ) );
  MUX21X1 U9077 ( .IN1(n8900), .IN2(n8901), .S(n8902), .Q(n8899) );
  NAND3X0 U9078 ( .IN1(n8897), .IN2(n8903), .IN3(n8856), .QN(n8901) );
  NAND2X0 U9079 ( .IN1(mul_frac_out[8]), .IN2(n1407), .QN(n8898) );
  NAND3X0 U9080 ( .IN1(n8904), .IN2(n8851), .IN3(n8905), .QN(
        \fpu_mul_frac_dp/n964 ) );
  MUX21X1 U9081 ( .IN1(n8906), .IN2(n8907), .S(n8908), .Q(n8905) );
  NAND2X0 U9082 ( .IN1(n8856), .IN2(n8909), .QN(n8907) );
  NAND2X0 U9083 ( .IN1(mul_frac_out[9]), .IN2(n1407), .QN(n8904) );
  NAND3X0 U9084 ( .IN1(n8910), .IN2(n8851), .IN3(n8911), .QN(
        \fpu_mul_frac_dp/n963 ) );
  MUX21X1 U9085 ( .IN1(n8912), .IN2(n8913), .S(n8914), .Q(n8911) );
  NAND3X0 U9086 ( .IN1(n8909), .IN2(n8915), .IN3(n8856), .QN(n8913) );
  NAND2X0 U9087 ( .IN1(mul_frac_out[10]), .IN2(n1407), .QN(n8910) );
  NAND3X0 U9088 ( .IN1(n8916), .IN2(n8851), .IN3(n8917), .QN(
        \fpu_mul_frac_dp/n962 ) );
  MUX21X1 U9089 ( .IN1(n8918), .IN2(n8919), .S(n8920), .Q(n8917) );
  NAND2X0 U9090 ( .IN1(n8856), .IN2(n8921), .QN(n8919) );
  NAND2X0 U9091 ( .IN1(mul_frac_out[11]), .IN2(n1407), .QN(n8916) );
  NAND3X0 U9092 ( .IN1(n8922), .IN2(n8851), .IN3(n8923), .QN(
        \fpu_mul_frac_dp/n961 ) );
  MUX21X1 U9093 ( .IN1(n8924), .IN2(n8925), .S(n8926), .Q(n8923) );
  NAND3X0 U9094 ( .IN1(n8921), .IN2(n8927), .IN3(n8856), .QN(n8925) );
  NAND2X0 U9095 ( .IN1(mul_frac_out[12]), .IN2(n1407), .QN(n8922) );
  NAND3X0 U9096 ( .IN1(n8928), .IN2(n8851), .IN3(n8929), .QN(
        \fpu_mul_frac_dp/n960 ) );
  MUX21X1 U9097 ( .IN1(n8930), .IN2(n8931), .S(n8932), .Q(n8929) );
  NAND2X0 U9098 ( .IN1(n8856), .IN2(n8933), .QN(n8931) );
  NAND2X0 U9099 ( .IN1(mul_frac_out[13]), .IN2(n1407), .QN(n8928) );
  NAND3X0 U9100 ( .IN1(n8934), .IN2(n8851), .IN3(n8935), .QN(
        \fpu_mul_frac_dp/n959 ) );
  MUX21X1 U9101 ( .IN1(n8936), .IN2(n8937), .S(n8938), .Q(n8935) );
  NAND3X0 U9102 ( .IN1(n8933), .IN2(n8939), .IN3(n8856), .QN(n8937) );
  NAND2X0 U9103 ( .IN1(mul_frac_out[14]), .IN2(n1408), .QN(n8934) );
  NAND3X0 U9104 ( .IN1(n8940), .IN2(n8851), .IN3(n8941), .QN(
        \fpu_mul_frac_dp/n958 ) );
  MUX21X1 U9105 ( .IN1(n8942), .IN2(n8943), .S(n8944), .Q(n8941) );
  NAND2X0 U9106 ( .IN1(n8856), .IN2(n8945), .QN(n8943) );
  NAND2X0 U9107 ( .IN1(mul_frac_out[15]), .IN2(n1408), .QN(n8940) );
  NAND3X0 U9108 ( .IN1(n8946), .IN2(n8851), .IN3(n8947), .QN(
        \fpu_mul_frac_dp/n957 ) );
  MUX21X1 U9109 ( .IN1(n8948), .IN2(n8949), .S(n8950), .Q(n8947) );
  NAND3X0 U9110 ( .IN1(n8945), .IN2(n8951), .IN3(n8856), .QN(n8949) );
  NAND2X0 U9111 ( .IN1(mul_frac_out[16]), .IN2(n1408), .QN(n8946) );
  NAND3X0 U9112 ( .IN1(n8952), .IN2(n8851), .IN3(n8953), .QN(
        \fpu_mul_frac_dp/n956 ) );
  MUX21X1 U9113 ( .IN1(n8954), .IN2(n8955), .S(n8956), .Q(n8953) );
  NAND2X0 U9114 ( .IN1(n8856), .IN2(n8957), .QN(n8955) );
  NAND2X0 U9115 ( .IN1(mul_frac_out[17]), .IN2(n1408), .QN(n8952) );
  NAND3X0 U9116 ( .IN1(n8958), .IN2(n8851), .IN3(n8959), .QN(
        \fpu_mul_frac_dp/n955 ) );
  MUX21X1 U9117 ( .IN1(n8960), .IN2(n8961), .S(n8962), .Q(n8959) );
  NAND3X0 U9118 ( .IN1(n8957), .IN2(n8963), .IN3(n8856), .QN(n8961) );
  NAND2X0 U9119 ( .IN1(mul_frac_out[18]), .IN2(n1408), .QN(n8958) );
  NAND3X0 U9120 ( .IN1(n8964), .IN2(n8851), .IN3(n8965), .QN(
        \fpu_mul_frac_dp/n954 ) );
  MUX21X1 U9121 ( .IN1(n8966), .IN2(n8967), .S(n8968), .Q(n8965) );
  NAND2X0 U9122 ( .IN1(n8856), .IN2(n8969), .QN(n8967) );
  NAND2X0 U9123 ( .IN1(mul_frac_out[19]), .IN2(n1408), .QN(n8964) );
  NAND3X0 U9124 ( .IN1(n8970), .IN2(n8851), .IN3(n8971), .QN(
        \fpu_mul_frac_dp/n953 ) );
  MUX21X1 U9125 ( .IN1(n8972), .IN2(n8973), .S(n8974), .Q(n8971) );
  NAND3X0 U9126 ( .IN1(n8969), .IN2(n8975), .IN3(n8856), .QN(n8973) );
  NAND2X0 U9127 ( .IN1(mul_frac_out[20]), .IN2(n1408), .QN(n8970) );
  NAND3X0 U9128 ( .IN1(n8976), .IN2(n8851), .IN3(n8977), .QN(
        \fpu_mul_frac_dp/n952 ) );
  MUX21X1 U9129 ( .IN1(n8978), .IN2(n8979), .S(n8980), .Q(n8977) );
  NAND2X0 U9130 ( .IN1(n8856), .IN2(n8981), .QN(n8978) );
  NAND2X0 U9131 ( .IN1(mul_frac_out[21]), .IN2(n1408), .QN(n8976) );
  NAND3X0 U9132 ( .IN1(n8982), .IN2(n8851), .IN3(n8983), .QN(
        \fpu_mul_frac_dp/n951 ) );
  MUX21X1 U9133 ( .IN1(n8984), .IN2(n8985), .S(n8986), .Q(n8983) );
  NAND3X0 U9134 ( .IN1(n8981), .IN2(n8980), .IN3(n8856), .QN(n8984) );
  NAND2X0 U9135 ( .IN1(mul_frac_out[22]), .IN2(n1408), .QN(n8982) );
  NAND3X0 U9136 ( .IN1(n8987), .IN2(n8851), .IN3(n8988), .QN(
        \fpu_mul_frac_dp/n950 ) );
  MUX21X1 U9137 ( .IN1(n8989), .IN2(n8990), .S(n8991), .Q(n8988) );
  NAND2X0 U9138 ( .IN1(n8856), .IN2(n8992), .QN(n8989) );
  NAND2X0 U9139 ( .IN1(mul_frac_out[23]), .IN2(n1408), .QN(n8987) );
  NAND3X0 U9140 ( .IN1(n8993), .IN2(n8851), .IN3(n8994), .QN(
        \fpu_mul_frac_dp/n949 ) );
  MUX21X1 U9141 ( .IN1(n8995), .IN2(n8996), .S(n8997), .Q(n8994) );
  NAND2X0 U9142 ( .IN1(mul_frac_out[24]), .IN2(n1408), .QN(n8993) );
  NAND3X0 U9143 ( .IN1(n8998), .IN2(n8851), .IN3(n8999), .QN(
        \fpu_mul_frac_dp/n948 ) );
  MUX21X1 U9144 ( .IN1(n9000), .IN2(n9001), .S(n9002), .Q(n8999) );
  NAND2X0 U9145 ( .IN1(n9003), .IN2(n8997), .QN(n9000) );
  NAND2X0 U9146 ( .IN1(mul_frac_out[25]), .IN2(n1408), .QN(n8998) );
  NAND3X0 U9147 ( .IN1(n9004), .IN2(n8851), .IN3(n9005), .QN(
        \fpu_mul_frac_dp/n947 ) );
  MUX21X1 U9148 ( .IN1(n9006), .IN2(n9007), .S(n9008), .Q(n9005) );
  NAND3X0 U9149 ( .IN1(n8997), .IN2(n9002), .IN3(n9003), .QN(n9006) );
  INVX0 U9150 ( .INP(n8995), .ZN(n9003) );
  NAND3X0 U9151 ( .IN1(n8992), .IN2(n8991), .IN3(n8856), .QN(n8995) );
  NAND2X0 U9152 ( .IN1(mul_frac_out[26]), .IN2(n1408), .QN(n9004) );
  NAND3X0 U9153 ( .IN1(n9009), .IN2(n8851), .IN3(n9010), .QN(
        \fpu_mul_frac_dp/n946 ) );
  MUX21X1 U9154 ( .IN1(n9011), .IN2(n9012), .S(n9013), .Q(n9010) );
  NAND2X0 U9155 ( .IN1(n8856), .IN2(n9014), .QN(n9011) );
  NAND2X0 U9156 ( .IN1(mul_frac_out[27]), .IN2(n1408), .QN(n9009) );
  NAND3X0 U9157 ( .IN1(n9015), .IN2(n8851), .IN3(n9016), .QN(
        \fpu_mul_frac_dp/n945 ) );
  MUX21X1 U9158 ( .IN1(n9017), .IN2(n9018), .S(n9019), .Q(n9016) );
  OA21X1 U9159 ( .IN1(n9013), .IN2(n1796), .IN3(n9012), .Q(n9018) );
  OA21X1 U9160 ( .IN1(n1796), .IN2(n9008), .IN3(n9007), .Q(n9012) );
  OA21X1 U9161 ( .IN1(n1796), .IN2(n9002), .IN3(n9001), .Q(n9007) );
  OA21X1 U9162 ( .IN1(n1796), .IN2(n8997), .IN3(n8996), .Q(n9001) );
  OA21X1 U9163 ( .IN1(n1796), .IN2(n8991), .IN3(n8990), .Q(n8996) );
  OA21X1 U9164 ( .IN1(n1796), .IN2(n8986), .IN3(n8985), .Q(n8990) );
  OA21X1 U9165 ( .IN1(n1796), .IN2(n8980), .IN3(n8979), .Q(n8985) );
  OA21X1 U9166 ( .IN1(n1796), .IN2(n9020), .IN3(n8972), .Q(n8979) );
  OA21X1 U9167 ( .IN1(n1796), .IN2(n8975), .IN3(n8966), .Q(n8972) );
  OA21X1 U9168 ( .IN1(n1796), .IN2(n9021), .IN3(n8960), .Q(n8966) );
  OA21X1 U9169 ( .IN1(n1796), .IN2(n8963), .IN3(n8954), .Q(n8960) );
  OA21X1 U9170 ( .IN1(n1796), .IN2(n9022), .IN3(n8948), .Q(n8954) );
  OA21X1 U9171 ( .IN1(n1796), .IN2(n8951), .IN3(n8942), .Q(n8948) );
  OA21X1 U9172 ( .IN1(n1796), .IN2(n9023), .IN3(n8936), .Q(n8942) );
  OA21X1 U9173 ( .IN1(n1796), .IN2(n8939), .IN3(n8930), .Q(n8936) );
  OA21X1 U9174 ( .IN1(n1796), .IN2(n9024), .IN3(n8924), .Q(n8930) );
  OA21X1 U9175 ( .IN1(n1796), .IN2(n8927), .IN3(n8918), .Q(n8924) );
  OA21X1 U9176 ( .IN1(n1796), .IN2(n9025), .IN3(n8912), .Q(n8918) );
  OA21X1 U9177 ( .IN1(n1796), .IN2(n8915), .IN3(n8906), .Q(n8912) );
  OA21X1 U9178 ( .IN1(n1796), .IN2(n9026), .IN3(n8900), .Q(n8906) );
  OA21X1 U9179 ( .IN1(n1796), .IN2(n8903), .IN3(n8894), .Q(n8900) );
  OA21X1 U9180 ( .IN1(n1796), .IN2(n9027), .IN3(n8888), .Q(n8894) );
  OA21X1 U9181 ( .IN1(n1796), .IN2(n8891), .IN3(n8882), .Q(n8888) );
  OA21X1 U9182 ( .IN1(n1796), .IN2(n9028), .IN3(n8876), .Q(n8882) );
  OA21X1 U9183 ( .IN1(n1796), .IN2(n8879), .IN3(n8870), .Q(n8876) );
  OA21X1 U9184 ( .IN1(n1796), .IN2(n8866), .IN3(n8865), .Q(n8870) );
  OA21X1 U9185 ( .IN1(n1796), .IN2(n9029), .IN3(n8859), .Q(n8865) );
  OA21X1 U9186 ( .IN1(n1796), .IN2(n8867), .IN3(n8853), .Q(n8859) );
  OA21X1 U9187 ( .IN1(n1796), .IN2(m5stg_fmulda), .IN3(n9030), .Q(n8853) );
  NAND3X0 U9188 ( .IN1(n9014), .IN2(n9013), .IN3(n8856), .QN(n9017) );
  NAND2X0 U9189 ( .IN1(mul_frac_out[28]), .IN2(n1408), .QN(n9015) );
  AO221X1 U9190 ( .IN1(n9031), .IN2(n9032), .IN3(mul_frac_out[29]), .IN4(n1383), .IN5(n9033), .Q(\fpu_mul_frac_dp/n944 ) );
  AO21X1 U9191 ( .IN1(n9034), .IN2(n8856), .IN3(n9035), .Q(n9033) );
  XOR3X1 U9192 ( .IN1(m5stg_fmuls), .IN2(n9036), .IN3(n9037), .Q(n9034) );
  INVX0 U9193 ( .INP(n9030), .ZN(n9031) );
  NAND3X0 U9194 ( .IN1(n9038), .IN2(n8851), .IN3(n9039), .QN(
        \fpu_mul_frac_dp/n943 ) );
  MUX21X1 U9195 ( .IN1(n9040), .IN2(n9041), .S(n9042), .Q(n9039) );
  NAND2X0 U9196 ( .IN1(n8856), .IN2(n9043), .QN(n9041) );
  NAND2X0 U9197 ( .IN1(mul_frac_out[30]), .IN2(n1408), .QN(n9038) );
  NAND3X0 U9198 ( .IN1(n9044), .IN2(n8851), .IN3(n9045), .QN(
        \fpu_mul_frac_dp/n942 ) );
  MUX21X1 U9199 ( .IN1(n9046), .IN2(n9047), .S(n9048), .Q(n9045) );
  NAND3X0 U9200 ( .IN1(n9043), .IN2(n9049), .IN3(n8856), .QN(n9046) );
  NAND2X0 U9201 ( .IN1(mul_frac_out[31]), .IN2(n1407), .QN(n9044) );
  NAND3X0 U9202 ( .IN1(n9050), .IN2(n8851), .IN3(n9051), .QN(
        \fpu_mul_frac_dp/n941 ) );
  MUX21X1 U9203 ( .IN1(n9052), .IN2(n9053), .S(n9054), .Q(n9051) );
  NAND2X0 U9204 ( .IN1(n8856), .IN2(n9055), .QN(n9053) );
  NAND2X0 U9205 ( .IN1(mul_frac_out[32]), .IN2(n1407), .QN(n9050) );
  NAND3X0 U9206 ( .IN1(n9056), .IN2(n8851), .IN3(n9057), .QN(
        \fpu_mul_frac_dp/n940 ) );
  MUX21X1 U9207 ( .IN1(n9058), .IN2(n9059), .S(n9060), .Q(n9057) );
  NAND3X0 U9208 ( .IN1(n9055), .IN2(n9061), .IN3(n8856), .QN(n9058) );
  NAND2X0 U9209 ( .IN1(mul_frac_out[33]), .IN2(n1407), .QN(n9056) );
  NAND3X0 U9210 ( .IN1(n9062), .IN2(n8851), .IN3(n9063), .QN(
        \fpu_mul_frac_dp/n939 ) );
  MUX21X1 U9211 ( .IN1(n9064), .IN2(n9065), .S(n9066), .Q(n9063) );
  NAND2X0 U9212 ( .IN1(n8856), .IN2(n9067), .QN(n9065) );
  NAND2X0 U9213 ( .IN1(mul_frac_out[34]), .IN2(n1406), .QN(n9062) );
  NAND3X0 U9214 ( .IN1(n9068), .IN2(n8851), .IN3(n9069), .QN(
        \fpu_mul_frac_dp/n938 ) );
  MUX21X1 U9215 ( .IN1(n9070), .IN2(n9071), .S(n9072), .Q(n9069) );
  NAND3X0 U9216 ( .IN1(n9067), .IN2(n9073), .IN3(n8856), .QN(n9070) );
  NAND2X0 U9217 ( .IN1(mul_frac_out[35]), .IN2(n1406), .QN(n9068) );
  NAND3X0 U9218 ( .IN1(n9074), .IN2(n8851), .IN3(n9075), .QN(
        \fpu_mul_frac_dp/n937 ) );
  MUX21X1 U9219 ( .IN1(n9076), .IN2(n9077), .S(n9078), .Q(n9075) );
  NAND2X0 U9220 ( .IN1(n8856), .IN2(n9079), .QN(n9077) );
  NAND2X0 U9221 ( .IN1(mul_frac_out[36]), .IN2(n1406), .QN(n9074) );
  NAND3X0 U9222 ( .IN1(n9080), .IN2(n8851), .IN3(n9081), .QN(
        \fpu_mul_frac_dp/n936 ) );
  MUX21X1 U9223 ( .IN1(n9082), .IN2(n9083), .S(n9084), .Q(n9081) );
  NAND3X0 U9224 ( .IN1(n9079), .IN2(n9085), .IN3(n8856), .QN(n9082) );
  NAND2X0 U9225 ( .IN1(mul_frac_out[37]), .IN2(n1406), .QN(n9080) );
  NAND3X0 U9226 ( .IN1(n9086), .IN2(n8851), .IN3(n9087), .QN(
        \fpu_mul_frac_dp/n935 ) );
  MUX21X1 U9227 ( .IN1(n9088), .IN2(n9089), .S(n9090), .Q(n9087) );
  NAND2X0 U9228 ( .IN1(n8856), .IN2(n9091), .QN(n9088) );
  NAND2X0 U9229 ( .IN1(mul_frac_out[38]), .IN2(n1407), .QN(n9086) );
  NAND3X0 U9230 ( .IN1(n9092), .IN2(n8851), .IN3(n9093), .QN(
        \fpu_mul_frac_dp/n934 ) );
  MUX21X1 U9231 ( .IN1(n9094), .IN2(n9095), .S(n9096), .Q(n9093) );
  NAND3X0 U9232 ( .IN1(n9091), .IN2(n9090), .IN3(n8856), .QN(n9094) );
  NAND2X0 U9233 ( .IN1(mul_frac_out[39]), .IN2(n1406), .QN(n9092) );
  NAND3X0 U9234 ( .IN1(n9097), .IN2(n8851), .IN3(n9098), .QN(
        \fpu_mul_frac_dp/n933 ) );
  MUX21X1 U9235 ( .IN1(n9099), .IN2(n9100), .S(n9101), .Q(n9098) );
  NAND2X0 U9236 ( .IN1(n8856), .IN2(n9102), .QN(n9099) );
  NAND2X0 U9237 ( .IN1(mul_frac_out[40]), .IN2(n1406), .QN(n9097) );
  NAND3X0 U9238 ( .IN1(n9103), .IN2(n8851), .IN3(n9104), .QN(
        \fpu_mul_frac_dp/n932 ) );
  MUX21X1 U9239 ( .IN1(n9105), .IN2(n9106), .S(n9107), .Q(n9104) );
  NAND3X0 U9240 ( .IN1(n9102), .IN2(n9101), .IN3(n8856), .QN(n9105) );
  NAND2X0 U9241 ( .IN1(mul_frac_out[41]), .IN2(n1406), .QN(n9103) );
  NAND3X0 U9242 ( .IN1(n9108), .IN2(n8851), .IN3(n9109), .QN(
        \fpu_mul_frac_dp/n931 ) );
  MUX21X1 U9243 ( .IN1(n9110), .IN2(n9111), .S(n9112), .Q(n9109) );
  NAND2X0 U9244 ( .IN1(n8856), .IN2(n9113), .QN(n9110) );
  NAND2X0 U9245 ( .IN1(mul_frac_out[42]), .IN2(n1406), .QN(n9108) );
  NAND3X0 U9246 ( .IN1(n9114), .IN2(n8851), .IN3(n9115), .QN(
        \fpu_mul_frac_dp/n930 ) );
  MUX21X1 U9247 ( .IN1(n9116), .IN2(n9117), .S(n9118), .Q(n9115) );
  NAND2X0 U9248 ( .IN1(mul_frac_out[43]), .IN2(n1406), .QN(n9114) );
  NAND3X0 U9249 ( .IN1(n9119), .IN2(n8851), .IN3(n9120), .QN(
        \fpu_mul_frac_dp/n929 ) );
  MUX21X1 U9250 ( .IN1(n9121), .IN2(n9122), .S(n9123), .Q(n9120) );
  NAND2X0 U9251 ( .IN1(n9124), .IN2(n9118), .QN(n9121) );
  NAND2X0 U9252 ( .IN1(mul_frac_out[44]), .IN2(n1406), .QN(n9119) );
  NAND3X0 U9253 ( .IN1(n9125), .IN2(n8851), .IN3(n9126), .QN(
        \fpu_mul_frac_dp/n928 ) );
  MUX21X1 U9254 ( .IN1(n9127), .IN2(n9128), .S(n9129), .Q(n9126) );
  NAND3X0 U9255 ( .IN1(n9123), .IN2(n9118), .IN3(n9124), .QN(n9127) );
  INVX0 U9256 ( .INP(n9116), .ZN(n9124) );
  NAND3X0 U9257 ( .IN1(n9113), .IN2(n9112), .IN3(n8856), .QN(n9116) );
  NAND2X0 U9258 ( .IN1(mul_frac_out[45]), .IN2(n1406), .QN(n9125) );
  NAND3X0 U9259 ( .IN1(n9130), .IN2(n8851), .IN3(n9131), .QN(
        \fpu_mul_frac_dp/n927 ) );
  MUX21X1 U9260 ( .IN1(n9132), .IN2(n9133), .S(n9134), .Q(n9131) );
  NAND2X0 U9261 ( .IN1(n8856), .IN2(n9135), .QN(n9132) );
  NAND2X0 U9262 ( .IN1(mul_frac_out[46]), .IN2(n1406), .QN(n9130) );
  NAND3X0 U9263 ( .IN1(n9136), .IN2(n8851), .IN3(n9137), .QN(
        \fpu_mul_frac_dp/n926 ) );
  MUX21X1 U9264 ( .IN1(n9138), .IN2(n9139), .S(n9140), .Q(n9137) );
  NAND3X0 U9265 ( .IN1(n9135), .IN2(n9134), .IN3(n8856), .QN(n9138) );
  NAND2X0 U9266 ( .IN1(mul_frac_out[47]), .IN2(n1406), .QN(n9136) );
  NAND3X0 U9267 ( .IN1(n9141), .IN2(n8851), .IN3(n9142), .QN(
        \fpu_mul_frac_dp/n925 ) );
  MUX21X1 U9268 ( .IN1(n9143), .IN2(n9144), .S(n9145), .Q(n9142) );
  NAND2X0 U9269 ( .IN1(n8856), .IN2(n9146), .QN(n9143) );
  NAND2X0 U9270 ( .IN1(mul_frac_out[48]), .IN2(n1406), .QN(n9141) );
  NAND3X0 U9271 ( .IN1(n9147), .IN2(n8851), .IN3(n9148), .QN(
        \fpu_mul_frac_dp/n924 ) );
  MUX21X1 U9272 ( .IN1(n9149), .IN2(n9150), .S(n9151), .Q(n9148) );
  NAND3X0 U9273 ( .IN1(n9146), .IN2(n9145), .IN3(n8856), .QN(n9149) );
  NAND2X0 U9274 ( .IN1(mul_frac_out[49]), .IN2(n1406), .QN(n9147) );
  NAND3X0 U9275 ( .IN1(n9152), .IN2(n8851), .IN3(n9153), .QN(
        \fpu_mul_frac_dp/n923 ) );
  MUX21X1 U9276 ( .IN1(n9154), .IN2(n9155), .S(n9156), .Q(n9153) );
  NAND2X0 U9277 ( .IN1(n8856), .IN2(n9157), .QN(n9154) );
  NAND2X0 U9278 ( .IN1(mul_frac_out[50]), .IN2(n1406), .QN(n9152) );
  NAND3X0 U9279 ( .IN1(n9158), .IN2(n8851), .IN3(n9159), .QN(
        \fpu_mul_frac_dp/n922 ) );
  MUX21X1 U9280 ( .IN1(n9160), .IN2(n9161), .S(n9162), .Q(n9159) );
  NAND3X0 U9281 ( .IN1(n9157), .IN2(n9156), .IN3(n8856), .QN(n9161) );
  INVX0 U9282 ( .INP(n1796), .ZN(n8856) );
  OA21X1 U9283 ( .IN1(n1796), .IN2(n9156), .IN3(n9155), .Q(n9160) );
  OA21X1 U9284 ( .IN1(n9151), .IN2(n1796), .IN3(n9150), .Q(n9155) );
  OA21X1 U9285 ( .IN1(n9145), .IN2(n1796), .IN3(n9144), .Q(n9150) );
  OA21X1 U9286 ( .IN1(n9140), .IN2(n1796), .IN3(n9139), .Q(n9144) );
  OA21X1 U9287 ( .IN1(n9134), .IN2(n1796), .IN3(n9133), .Q(n9139) );
  OA21X1 U9288 ( .IN1(n9129), .IN2(n1796), .IN3(n9128), .Q(n9133) );
  OA21X1 U9289 ( .IN1(n9123), .IN2(n1796), .IN3(n9122), .Q(n9128) );
  OA21X1 U9290 ( .IN1(n9118), .IN2(n1796), .IN3(n9117), .Q(n9122) );
  OA21X1 U9291 ( .IN1(n9112), .IN2(n1796), .IN3(n9111), .Q(n9117) );
  OA21X1 U9292 ( .IN1(n9107), .IN2(n1796), .IN3(n9106), .Q(n9111) );
  OA21X1 U9293 ( .IN1(n9101), .IN2(n1796), .IN3(n9100), .Q(n9106) );
  OA21X1 U9294 ( .IN1(n9096), .IN2(n1796), .IN3(n9095), .Q(n9100) );
  OA21X1 U9295 ( .IN1(n9090), .IN2(n1796), .IN3(n9089), .Q(n9095) );
  OA21X1 U9296 ( .IN1(n9084), .IN2(n1796), .IN3(n9083), .Q(n9089) );
  OA21X1 U9297 ( .IN1(n9085), .IN2(n1796), .IN3(n9076), .Q(n9083) );
  OA21X1 U9298 ( .IN1(n9072), .IN2(n1796), .IN3(n9071), .Q(n9076) );
  OA21X1 U9299 ( .IN1(n9073), .IN2(n1796), .IN3(n9064), .Q(n9071) );
  OA21X1 U9300 ( .IN1(n9060), .IN2(n1796), .IN3(n9059), .Q(n9064) );
  OA21X1 U9301 ( .IN1(n9061), .IN2(n1796), .IN3(n9052), .Q(n9059) );
  OA21X1 U9302 ( .IN1(n9048), .IN2(n1796), .IN3(n9047), .Q(n9052) );
  OA21X1 U9303 ( .IN1(n9049), .IN2(n1796), .IN3(n9040), .Q(n9047) );
  OA21X1 U9304 ( .IN1(n9043), .IN2(n1796), .IN3(n9030), .Q(n9040) );
  NAND2X0 U9305 ( .IN1(n1775), .IN2(n1608), .QN(n9030) );
  NOR2X0 U9306 ( .IN1(n9163), .IN2(n9164), .QN(n1775) );
  NAND3X0 U9307 ( .IN1(n1592), .IN2(n1773), .IN3(n9163), .QN(n1796) );
  NOR2X0 U9308 ( .IN1(n1751), .IN2(n1778), .QN(n9035) );
  NAND2X0 U9309 ( .IN1(mul_frac_out[51]), .IN2(n1406), .QN(n9158) );
  NOR2X0 U9310 ( .IN1(\fpu_mul_frac_dp/n383 ), .IN2(n709), .QN(
        \fpu_mul_frac_dp/n832 ) );
  INVX0 U9311 ( .INP(rclk), .ZN(n709) );
  AO22X1 U9312 ( .IN1(inq_in1[0]), .IN2(n1604), .IN3(n1387), .IN4(n1208), .Q(
        \fpu_mul_frac_dp/n1097 ) );
  AO22X1 U9313 ( .IN1(inq_in1[1]), .IN2(n1604), .IN3(n1387), .IN4(n956), .Q(
        \fpu_mul_frac_dp/n1096 ) );
  AO22X1 U9314 ( .IN1(inq_in1[2]), .IN2(n1604), .IN3(n1387), .IN4(n1311), .Q(
        \fpu_mul_frac_dp/n1095 ) );
  AO22X1 U9315 ( .IN1(inq_in1[3]), .IN2(n1604), .IN3(n1387), .IN4(n1180), .Q(
        \fpu_mul_frac_dp/n1094 ) );
  AO22X1 U9316 ( .IN1(inq_in1[4]), .IN2(n1604), .IN3(n1387), .IN4(n1316), .Q(
        \fpu_mul_frac_dp/n1093 ) );
  AO22X1 U9317 ( .IN1(inq_in1[5]), .IN2(n1604), .IN3(n1387), .IN4(n1312), .Q(
        \fpu_mul_frac_dp/n1092 ) );
  AO22X1 U9318 ( .IN1(inq_in1[6]), .IN2(n1604), .IN3(n1387), .IN4(n943), .Q(
        \fpu_mul_frac_dp/n1091 ) );
  AO22X1 U9319 ( .IN1(inq_in1[7]), .IN2(n1604), .IN3(n1387), .IN4(n1317), .Q(
        \fpu_mul_frac_dp/n1090 ) );
  AO22X1 U9320 ( .IN1(inq_in1[8]), .IN2(n1605), .IN3(n1388), .IN4(n1186), .Q(
        \fpu_mul_frac_dp/n1089 ) );
  AO22X1 U9321 ( .IN1(inq_in1[9]), .IN2(n1605), .IN3(n1388), .IN4(n952), .Q(
        \fpu_mul_frac_dp/n1088 ) );
  AO22X1 U9322 ( .IN1(inq_in1[10]), .IN2(n1605), .IN3(n1388), .IN4(n1171), .Q(
        \fpu_mul_frac_dp/n1087 ) );
  AO22X1 U9323 ( .IN1(inq_in1[11]), .IN2(n1605), .IN3(n1388), .IN4(n1121), .Q(
        \fpu_mul_frac_dp/n1086 ) );
  AO22X1 U9324 ( .IN1(inq_in1[12]), .IN2(n1605), .IN3(\fpu_mul_frac_dp/n836 ), 
        .IN4(n1385), .Q(\fpu_mul_frac_dp/n1085 ) );
  AO22X1 U9325 ( .IN1(inq_in1[13]), .IN2(n1605), .IN3(n1388), .IN4(n1314), .Q(
        \fpu_mul_frac_dp/n1084 ) );
  AO22X1 U9326 ( .IN1(inq_in1[14]), .IN2(n1605), .IN3(n1388), .IN4(n1310), .Q(
        \fpu_mul_frac_dp/n1083 ) );
  AO22X1 U9327 ( .IN1(inq_in1[15]), .IN2(n1605), .IN3(n1388), .IN4(n1202), .Q(
        \fpu_mul_frac_dp/n1082 ) );
  AO22X1 U9328 ( .IN1(inq_in1[16]), .IN2(n1605), .IN3(n1388), .IN4(n1159), .Q(
        \fpu_mul_frac_dp/n1081 ) );
  AO22X1 U9329 ( .IN1(inq_in1[17]), .IN2(n1605), .IN3(n1388), .IN4(n899), .Q(
        \fpu_mul_frac_dp/n1080 ) );
  AO22X1 U9330 ( .IN1(inq_in1[18]), .IN2(n1605), .IN3(n1388), .IN4(n960), .Q(
        \fpu_mul_frac_dp/n1079 ) );
  AO22X1 U9331 ( .IN1(inq_in1[19]), .IN2(n1605), .IN3(n1388), .IN4(n882), .Q(
        \fpu_mul_frac_dp/n1078 ) );
  AO22X1 U9332 ( .IN1(inq_in1[20]), .IN2(n1605), .IN3(n1388), .IN4(n1222), .Q(
        \fpu_mul_frac_dp/n1077 ) );
  AO22X1 U9333 ( .IN1(inq_in1[21]), .IN2(n1605), .IN3(n1388), .IN4(n985), .Q(
        \fpu_mul_frac_dp/n1076 ) );
  AO22X1 U9334 ( .IN1(inq_in1[22]), .IN2(n1605), .IN3(n1388), .IN4(n1221), .Q(
        \fpu_mul_frac_dp/n1075 ) );
  AO22X1 U9335 ( .IN1(inq_in1[23]), .IN2(n1605), .IN3(n1389), .IN4(n987), .Q(
        \fpu_mul_frac_dp/n1074 ) );
  AO22X1 U9336 ( .IN1(inq_in1[24]), .IN2(n1606), .IN3(n1389), .IN4(n1201), .Q(
        \fpu_mul_frac_dp/n1073 ) );
  AO22X1 U9337 ( .IN1(inq_in1[25]), .IN2(n1606), .IN3(n1389), .IN4(n978), .Q(
        \fpu_mul_frac_dp/n1072 ) );
  AO22X1 U9338 ( .IN1(inq_in1[26]), .IN2(n1605), .IN3(n1389), .IN4(n1220), .Q(
        \fpu_mul_frac_dp/n1071 ) );
  AO22X1 U9339 ( .IN1(inq_in1[27]), .IN2(n1606), .IN3(n1389), .IN4(n986), .Q(
        \fpu_mul_frac_dp/n1070 ) );
  AO22X1 U9340 ( .IN1(inq_in1[28]), .IN2(n1606), .IN3(\fpu_mul_frac_dp/n813 ), 
        .IN4(n1384), .Q(\fpu_mul_frac_dp/n1069 ) );
  AO22X1 U9341 ( .IN1(inq_in1[29]), .IN2(n1606), .IN3(n1389), .IN4(n1326), .Q(
        \fpu_mul_frac_dp/n1068 ) );
  AO22X1 U9342 ( .IN1(inq_in1[30]), .IN2(n1606), .IN3(n1389), .IN4(n1320), .Q(
        \fpu_mul_frac_dp/n1067 ) );
  AO22X1 U9343 ( .IN1(inq_in1[31]), .IN2(n1606), .IN3(n1389), .IN4(n1319), .Q(
        \fpu_mul_frac_dp/n1066 ) );
  AO22X1 U9344 ( .IN1(inq_in1[32]), .IN2(n1606), .IN3(n1389), .IN4(n967), .Q(
        \fpu_mul_frac_dp/n1065 ) );
  AO22X1 U9345 ( .IN1(inq_in1[33]), .IN2(n1606), .IN3(n1389), .IN4(n1183), .Q(
        \fpu_mul_frac_dp/n1064 ) );
  AO22X1 U9346 ( .IN1(inq_in1[34]), .IN2(n1606), .IN3(n1389), .IN4(n1302), .Q(
        \fpu_mul_frac_dp/n1063 ) );
  AO22X1 U9347 ( .IN1(inq_in1[35]), .IN2(n1606), .IN3(n1389), .IN4(n1182), .Q(
        \fpu_mul_frac_dp/n1062 ) );
  AO22X1 U9348 ( .IN1(inq_in1[36]), .IN2(n1606), .IN3(n1389), .IN4(n947), .Q(
        \fpu_mul_frac_dp/n1061 ) );
  AO22X1 U9349 ( .IN1(inq_in1[37]), .IN2(n1606), .IN3(n1389), .IN4(n1307), .Q(
        \fpu_mul_frac_dp/n1060 ) );
  AO22X1 U9350 ( .IN1(inq_in1[38]), .IN2(n1606), .IN3(n1390), .IN4(n1303), .Q(
        \fpu_mul_frac_dp/n1059 ) );
  AO22X1 U9351 ( .IN1(inq_in1[39]), .IN2(n1606), .IN3(n1390), .IN4(n1187), .Q(
        \fpu_mul_frac_dp/n1058 ) );
  AO22X1 U9352 ( .IN1(inq_in1[40]), .IN2(n1606), .IN3(n1390), .IN4(n1308), .Q(
        \fpu_mul_frac_dp/n1057 ) );
  AO22X1 U9353 ( .IN1(inq_in1[41]), .IN2(n1607), .IN3(n1390), .IN4(n1309), .Q(
        \fpu_mul_frac_dp/n1056 ) );
  AO22X1 U9354 ( .IN1(inq_in1[42]), .IN2(n1607), .IN3(n1390), .IN4(n1304), .Q(
        \fpu_mul_frac_dp/n1055 ) );
  AO22X1 U9355 ( .IN1(inq_in1[43]), .IN2(n1606), .IN3(n1390), .IN4(n1305), .Q(
        \fpu_mul_frac_dp/n1054 ) );
  AO22X1 U9356 ( .IN1(inq_in1[44]), .IN2(n1607), .IN3(n1390), .IN4(n973), .Q(
        \fpu_mul_frac_dp/n1053 ) );
  AO22X1 U9357 ( .IN1(inq_in1[45]), .IN2(n1607), .IN3(n1390), .IN4(n977), .Q(
        \fpu_mul_frac_dp/n1052 ) );
  AO22X1 U9358 ( .IN1(inq_in1[46]), .IN2(n1606), .IN3(n1390), .IN4(n1300), .Q(
        \fpu_mul_frac_dp/n1051 ) );
  AO22X1 U9359 ( .IN1(inq_in1[47]), .IN2(n1607), .IN3(n1390), .IN4(n1193), .Q(
        \fpu_mul_frac_dp/n1050 ) );
  AO22X1 U9360 ( .IN1(inq_in1[48]), .IN2(n1607), .IN3(n1390), .IN4(n1195), .Q(
        \fpu_mul_frac_dp/n1049 ) );
  AO22X1 U9361 ( .IN1(inq_in1[49]), .IN2(n1607), .IN3(n1387), .IN4(n1306), .Q(
        \fpu_mul_frac_dp/n1048 ) );
  AO22X1 U9362 ( .IN1(inq_in1[50]), .IN2(n1607), .IN3(n1390), .IN4(n1301), .Q(
        \fpu_mul_frac_dp/n1047 ) );
  AO22X1 U9363 ( .IN1(inq_in1[51]), .IN2(n1607), .IN3(n1402), .IN4(n1124), .Q(
        \fpu_mul_frac_dp/n1046 ) );
  AO22X1 U9364 ( .IN1(inq_in1[52]), .IN2(n1607), .IN3(n1400), .IN4(n1318), .Q(
        \fpu_mul_frac_dp/n1045 ) );
  AO22X1 U9365 ( .IN1(inq_in1[53]), .IN2(n1607), .IN3(n1400), .IN4(n1315), .Q(
        \fpu_mul_frac_dp/n1044 ) );
  AO21X1 U9366 ( .IN1(n1386), .IN2(n1200), .IN3(n1633), .Q(
        \fpu_mul_frac_dp/n1043 ) );
  AO22X1 U9367 ( .IN1(inq_in2[0]), .IN2(n1607), .IN3(n1401), .IN4(n1158), .Q(
        \fpu_mul_frac_dp/n1042 ) );
  AO22X1 U9368 ( .IN1(inq_in2[1]), .IN2(n1607), .IN3(n1400), .IN4(n939), .Q(
        \fpu_mul_frac_dp/n1041 ) );
  AO22X1 U9369 ( .IN1(inq_in2[2]), .IN2(n1607), .IN3(n1401), .IN4(n1147), .Q(
        \fpu_mul_frac_dp/n1040 ) );
  AO22X1 U9370 ( .IN1(inq_in2[3]), .IN2(n1607), .IN3(n1400), .IN4(n896), .Q(
        \fpu_mul_frac_dp/n1039 ) );
  AO22X1 U9371 ( .IN1(inq_in2[4]), .IN2(n1607), .IN3(n1401), .IN4(n1155), .Q(
        \fpu_mul_frac_dp/n1038 ) );
  AO22X1 U9372 ( .IN1(inq_in2[5]), .IN2(n1608), .IN3(n1401), .IN4(n941), .Q(
        \fpu_mul_frac_dp/n1037 ) );
  AO22X1 U9373 ( .IN1(inq_in2[6]), .IN2(n1607), .IN3(n1401), .IN4(n1149), .Q(
        \fpu_mul_frac_dp/n1036 ) );
  AO22X1 U9374 ( .IN1(inq_in2[7]), .IN2(n1608), .IN3(n1401), .IN4(n953), .Q(
        \fpu_mul_frac_dp/n1035 ) );
  AO22X1 U9375 ( .IN1(inq_in2[8]), .IN2(n1608), .IN3(n1401), .IN4(n898), .Q(
        \fpu_mul_frac_dp/n1034 ) );
  AO22X1 U9376 ( .IN1(inq_in2[9]), .IN2(n1608), .IN3(n1401), .IN4(n1137), .Q(
        \fpu_mul_frac_dp/n1033 ) );
  AO22X1 U9377 ( .IN1(inq_in2[10]), .IN2(n1608), .IN3(n1401), .IN4(n881), .Q(
        \fpu_mul_frac_dp/n1032 ) );
  AO22X1 U9378 ( .IN1(inq_in2[11]), .IN2(n1607), .IN3(n1401), .IN4(n925), .Q(
        \fpu_mul_frac_dp/n1031 ) );
  AO22X1 U9379 ( .IN1(inq_in2[12]), .IN2(n1608), .IN3(n1402), .IN4(n1113), .Q(
        \fpu_mul_frac_dp/n1030 ) );
  AO22X1 U9380 ( .IN1(inq_in2[13]), .IN2(n1608), .IN3(n1401), .IN4(n927), .Q(
        \fpu_mul_frac_dp/n1029 ) );
  AO22X1 U9381 ( .IN1(inq_in2[14]), .IN2(n1608), .IN3(n1400), .IN4(n1054), .Q(
        \fpu_mul_frac_dp/n1028 ) );
  AO22X1 U9382 ( .IN1(inq_in2[15]), .IN2(n1601), .IN3(n1402), .IN4(n892), .Q(
        \fpu_mul_frac_dp/n1027 ) );
  AO22X1 U9383 ( .IN1(inq_in2[16]), .IN2(n1599), .IN3(n1401), .IN4(n1141), .Q(
        \fpu_mul_frac_dp/n1026 ) );
  AO22X1 U9384 ( .IN1(inq_in2[17]), .IN2(n1600), .IN3(n1402), .IN4(n930), .Q(
        \fpu_mul_frac_dp/n1025 ) );
  AO22X1 U9385 ( .IN1(inq_in2[18]), .IN2(n1599), .IN3(n1402), .IN4(n1136), .Q(
        \fpu_mul_frac_dp/n1024 ) );
  AO22X1 U9386 ( .IN1(inq_in2[19]), .IN2(n1599), .IN3(n1402), .IN4(n932), .Q(
        \fpu_mul_frac_dp/n1023 ) );
  AO22X1 U9387 ( .IN1(inq_in2[20]), .IN2(n1600), .IN3(n1401), .IN4(n1156), .Q(
        \fpu_mul_frac_dp/n1022 ) );
  AO22X1 U9388 ( .IN1(inq_in2[21]), .IN2(n1599), .IN3(n1402), .IN4(n940), .Q(
        \fpu_mul_frac_dp/n1021 ) );
  AO22X1 U9389 ( .IN1(inq_in2[22]), .IN2(n1600), .IN3(n1402), .IN4(n1146), .Q(
        \fpu_mul_frac_dp/n1020 ) );
  AO22X1 U9390 ( .IN1(inq_in2[23]), .IN2(n1600), .IN3(n1403), .IN4(n955), .Q(
        \fpu_mul_frac_dp/n1019 ) );
  AO22X1 U9391 ( .IN1(inq_in2[24]), .IN2(n1600), .IN3(n1402), .IN4(n1157), .Q(
        \fpu_mul_frac_dp/n1018 ) );
  AO22X1 U9392 ( .IN1(inq_in2[25]), .IN2(n1600), .IN3(n1403), .IN4(n957), .Q(
        \fpu_mul_frac_dp/n1017 ) );
  AO22X1 U9393 ( .IN1(inq_in2[26]), .IN2(n1600), .IN3(n1402), .IN4(n897), .Q(
        \fpu_mul_frac_dp/n1016 ) );
  AO22X1 U9394 ( .IN1(inq_in2[27]), .IN2(n1600), .IN3(n1403), .IN4(n1148), .Q(
        \fpu_mul_frac_dp/n1015 ) );
  AO22X1 U9395 ( .IN1(inq_in2[28]), .IN2(n1600), .IN3(\fpu_mul_frac_dp/n837 ), 
        .IN4(n1385), .Q(\fpu_mul_frac_dp/n1014 ) );
  AO22X1 U9396 ( .IN1(inq_in2[29]), .IN2(n1600), .IN3(n1402), .IN4(n959), .Q(
        \fpu_mul_frac_dp/n1013 ) );
  AO22X1 U9397 ( .IN1(inq_in2[30]), .IN2(n1600), .IN3(n1403), .IN4(n1160), .Q(
        \fpu_mul_frac_dp/n1012 ) );
  AO22X1 U9398 ( .IN1(inq_in2[31]), .IN2(n1600), .IN3(n1402), .IN4(n958), .Q(
        \fpu_mul_frac_dp/n1011 ) );
  AO22X1 U9399 ( .IN1(inq_in2[32]), .IN2(n1600), .IN3(n1403), .IN4(n887), .Q(
        \fpu_mul_frac_dp/n1010 ) );
  AO22X1 U9400 ( .IN1(inq_in2[33]), .IN2(n1600), .IN3(n1401), .IN4(n1045), .Q(
        \fpu_mul_frac_dp/n1009 ) );
  AO22X1 U9401 ( .IN1(inq_in2[34]), .IN2(n1600), .IN3(n1403), .IN4(n919), .Q(
        \fpu_mul_frac_dp/n1008 ) );
  AO22X1 U9402 ( .IN1(inq_in2[35]), .IN2(n1600), .IN3(n1402), .IN4(n1046), .Q(
        \fpu_mul_frac_dp/n1007 ) );
  AO22X1 U9403 ( .IN1(inq_in2[36]), .IN2(n1600), .IN3(n1403), .IN4(n909), .Q(
        \fpu_mul_frac_dp/n1006 ) );
  AO22X1 U9404 ( .IN1(inq_in2[37]), .IN2(n1600), .IN3(n1403), .IN4(n1048), .Q(
        \fpu_mul_frac_dp/n1005 ) );
  AO22X1 U9405 ( .IN1(inq_in2[38]), .IN2(n1601), .IN3(n1403), .IN4(n920), .Q(
        \fpu_mul_frac_dp/n1004 ) );
  AO22X1 U9406 ( .IN1(inq_in2[39]), .IN2(n1601), .IN3(n1403), .IN4(n889), .Q(
        \fpu_mul_frac_dp/n1003 ) );
  AO22X1 U9407 ( .IN1(inq_in2[40]), .IN2(n1601), .IN3(n1403), .IN4(n1043), .Q(
        \fpu_mul_frac_dp/n1002 ) );
  AO22X1 U9408 ( .IN1(inq_in2[41]), .IN2(n1601), .IN3(n1402), .IN4(n921), .Q(
        \fpu_mul_frac_dp/n1001 ) );
  AO22X1 U9409 ( .IN1(inq_in2[42]), .IN2(n1601), .IN3(n1403), .IN4(n1047), .Q(
        \fpu_mul_frac_dp/n1000 ) );
  NAND2X0 U9410 ( .IN1(n9165), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N9 ) );
  NAND2X0 U9411 ( .IN1(n9167), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N8 ) );
  NAND2X0 U9412 ( .IN1(n9168), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N7 ) );
  NAND2X0 U9413 ( .IN1(n9169), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N6 ) );
  NAND2X0 U9414 ( .IN1(n9170), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N57 ) );
  NAND2X0 U9415 ( .IN1(n9171), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N56 ) );
  AO21X1 U9416 ( .IN1(n9172), .IN2(n1359), .IN3(n9173), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N55 ) );
  AO21X1 U9417 ( .IN1(n9174), .IN2(n1360), .IN3(n9173), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N54 ) );
  AO21X1 U9418 ( .IN1(n9175), .IN2(n1357), .IN3(n9173), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N53 ) );
  AO21X1 U9419 ( .IN1(n9176), .IN2(n1359), .IN3(n9173), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N52 ) );
  AO21X1 U9420 ( .IN1(n1033), .IN2(n1360), .IN3(n9177), .Q(n9173) );
  AO21X1 U9421 ( .IN1(n9178), .IN2(n1357), .IN3(n9177), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N51 ) );
  AO21X1 U9422 ( .IN1(n9179), .IN2(n1358), .IN3(n9177), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N50 ) );
  NAND2X0 U9423 ( .IN1(n9180), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N5 ) );
  AO21X1 U9424 ( .IN1(n9181), .IN2(n1359), .IN3(n9177), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N49 ) );
  AO21X1 U9425 ( .IN1(n9182), .IN2(n1360), .IN3(n9177), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N48 ) );
  AO21X1 U9426 ( .IN1(n9183), .IN2(n1357), .IN3(n9177), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N47 ) );
  AO21X1 U9427 ( .IN1(n9184), .IN2(n1358), .IN3(n9177), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N46 ) );
  AO21X1 U9428 ( .IN1(n9185), .IN2(n1359), .IN3(n9177), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N45 ) );
  AO21X1 U9429 ( .IN1(n9186), .IN2(n1360), .IN3(n9177), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N44 ) );
  AO21X1 U9430 ( .IN1(n9187), .IN2(n1357), .IN3(n9188), .Q(n9177) );
  NAND2X0 U9431 ( .IN1(n9189), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N43 ) );
  AO21X1 U9432 ( .IN1(n9190), .IN2(n1358), .IN3(n9191), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N42 ) );
  NAND2X0 U9433 ( .IN1(n9192), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N41 ) );
  NAND2X0 U9434 ( .IN1(n9193), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N40 ) );
  NAND2X0 U9435 ( .IN1(n9194), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N4 ) );
  AO21X1 U9436 ( .IN1(n9195), .IN2(n1359), .IN3(n9191), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N39 ) );
  AO21X1 U9437 ( .IN1(n9196), .IN2(n1360), .IN3(n9191), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N38 ) );
  AO21X1 U9438 ( .IN1(n9197), .IN2(n1357), .IN3(n9191), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N37 ) );
  AO21X1 U9439 ( .IN1(n1036), .IN2(n1358), .IN3(n9188), .Q(n9191) );
  INVX0 U9440 ( .INP(n9166), .ZN(n9188) );
  NAND2X0 U9441 ( .IN1(n9198), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N36 ) );
  NAND2X0 U9442 ( .IN1(n9199), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N35 ) );
  NAND2X0 U9443 ( .IN1(n9200), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N34 ) );
  NAND2X0 U9444 ( .IN1(n9201), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N33 ) );
  NAND2X0 U9445 ( .IN1(n9202), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N32 ) );
  NAND2X0 U9446 ( .IN1(n9203), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N31 ) );
  NAND2X0 U9447 ( .IN1(n9204), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N30 ) );
  NAND2X0 U9448 ( .IN1(n9205), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N29 ) );
  NAND2X0 U9449 ( .IN1(n9206), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N28 ) );
  NAND2X0 U9450 ( .IN1(n9207), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N27 ) );
  NAND2X0 U9451 ( .IN1(n9208), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N26 ) );
  NAND2X0 U9452 ( .IN1(n9209), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N25 ) );
  NAND2X0 U9453 ( .IN1(n9210), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N24 ) );
  NAND2X0 U9454 ( .IN1(n9211), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N23 ) );
  NAND2X0 U9455 ( .IN1(n9212), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N22 ) );
  NAND2X0 U9456 ( .IN1(n9213), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N21 ) );
  NAND2X0 U9457 ( .IN1(n9214), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N20 ) );
  NAND2X0 U9458 ( .IN1(n9215), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N19 ) );
  NAND2X0 U9459 ( .IN1(n9216), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N18 ) );
  NAND2X0 U9460 ( .IN1(n9217), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N17 ) );
  NAND2X0 U9461 ( .IN1(n9218), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N16 ) );
  NAND2X0 U9462 ( .IN1(n9219), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N15 ) );
  NAND2X0 U9463 ( .IN1(n9220), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N14 ) );
  NAND2X0 U9464 ( .IN1(n9221), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N13 ) );
  NAND2X0 U9465 ( .IN1(n9222), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N12 ) );
  NAND2X0 U9466 ( .IN1(n9223), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N11 ) );
  NAND2X0 U9467 ( .IN1(n9224), .IN2(n9166), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre4/N10 ) );
  AO21X1 U9468 ( .IN1(n9225), .IN2(n9226), .IN3(se_mul), .Q(n9166) );
  NAND2X0 U9469 ( .IN1(n9227), .IN2(n9228), .QN(n9226) );
  NAND2X0 U9470 ( .IN1(n9229), .IN2(n9224), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N9 ) );
  AO221X1 U9471 ( .IN1(n9227), .IN2(n9230), .IN3(n9231), .IN4(n9232), .IN5(
        n9233), .Q(n9224) );
  OAI21X1 U9472 ( .IN1(n9190), .IN2(\fpu_mul_frac_dp/n767 ), .IN3(n1359), .QN(
        n9233) );
  NAND2X0 U9473 ( .IN1(n9229), .IN2(n9165), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N8 ) );
  AO221X1 U9474 ( .IN1(n9234), .IN2(n9235), .IN3(n9231), .IN4(n9236), .IN5(
        n9237), .Q(n9165) );
  AO221X1 U9475 ( .IN1(n9238), .IN2(n9239), .IN3(n9227), .IN4(n9240), .IN5(
        se_mul), .Q(n9237) );
  NAND2X0 U9476 ( .IN1(n9229), .IN2(n9167), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N7 ) );
  AO221X1 U9477 ( .IN1(n9231), .IN2(n9241), .IN3(n9234), .IN4(n9242), .IN5(
        n9243), .Q(n9167) );
  AO221X1 U9478 ( .IN1(n9244), .IN2(n9239), .IN3(n9227), .IN4(n9245), .IN5(
        se_mul), .Q(n9243) );
  INVX0 U9479 ( .INP(n9246), .ZN(n9239) );
  NAND2X0 U9480 ( .IN1(n9229), .IN2(n9168), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N6 ) );
  AO221X1 U9481 ( .IN1(n9227), .IN2(n9247), .IN3(n9231), .IN4(n9248), .IN5(
        n9249), .Q(n9168) );
  AO21X1 U9482 ( .IN1(n9250), .IN2(n1036), .IN3(se_mul), .Q(n9249) );
  AO21X1 U9483 ( .IN1(n9251), .IN2(n1359), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N57 ) );
  NAND2X0 U9484 ( .IN1(n9229), .IN2(n9170), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N56 ) );
  AO21X1 U9485 ( .IN1(n9238), .IN2(n9227), .IN3(se_mul), .Q(n9170) );
  NAND2X0 U9486 ( .IN1(n9229), .IN2(n9171), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N55 ) );
  AO21X1 U9487 ( .IN1(n9244), .IN2(n9227), .IN3(se_mul), .Q(n9171) );
  AO21X1 U9488 ( .IN1(n9172), .IN2(n1360), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N54 ) );
  AO21X1 U9489 ( .IN1(n9174), .IN2(n1357), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N53 ) );
  INVX0 U9490 ( .INP(n9253), .ZN(n9174) );
  AO21X1 U9491 ( .IN1(n9175), .IN2(n1358), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N52 ) );
  INVX0 U9492 ( .INP(n9254), .ZN(n9175) );
  AO21X1 U9493 ( .IN1(n9176), .IN2(n1359), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N51 ) );
  AO21X1 U9494 ( .IN1(n9178), .IN2(n1360), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N50 ) );
  NAND2X0 U9495 ( .IN1(n9229), .IN2(n9169), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N5 ) );
  AO221X1 U9496 ( .IN1(n9227), .IN2(n9255), .IN3(n9231), .IN4(n9256), .IN5(
        n9257), .Q(n9169) );
  AO21X1 U9497 ( .IN1(n9258), .IN2(n1036), .IN3(se_mul), .Q(n9257) );
  AO21X1 U9498 ( .IN1(n9179), .IN2(n1357), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N49 ) );
  AO21X1 U9499 ( .IN1(n9181), .IN2(n1358), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N48 ) );
  AO21X1 U9500 ( .IN1(n9182), .IN2(n1359), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N47 ) );
  AO21X1 U9501 ( .IN1(n9183), .IN2(n1360), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N46 ) );
  AO21X1 U9502 ( .IN1(n9184), .IN2(n1357), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N45 ) );
  AO21X1 U9503 ( .IN1(n9185), .IN2(n1358), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N44 ) );
  AO21X1 U9504 ( .IN1(n9186), .IN2(n1359), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N43 ) );
  INVX0 U9505 ( .INP(n9259), .ZN(n9186) );
  NAND2X0 U9506 ( .IN1(n9229), .IN2(n9189), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N42 ) );
  AO221X1 U9507 ( .IN1(n9231), .IN2(n9228), .IN3(n9227), .IN4(n9260), .IN5(
        se_mul), .Q(n9189) );
  AO21X1 U9508 ( .IN1(n9190), .IN2(n1360), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N41 ) );
  MUX21X1 U9509 ( .IN1(n9261), .IN2(n9262), .S(\fpu_mul_frac_dp/n838 ), .Q(
        n9190) );
  NAND2X0 U9510 ( .IN1(n9263), .IN2(n1380), .QN(n9261) );
  NAND2X0 U9511 ( .IN1(n9229), .IN2(n9192), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N40 ) );
  AO221X1 U9512 ( .IN1(n9231), .IN2(n9238), .IN3(n9227), .IN4(n9235), .IN5(
        se_mul), .Q(n9192) );
  NAND2X0 U9513 ( .IN1(n9229), .IN2(n9180), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N4 ) );
  AO221X1 U9514 ( .IN1(n9227), .IN2(n9264), .IN3(n9231), .IN4(n9265), .IN5(
        n9266), .Q(n9180) );
  AO21X1 U9515 ( .IN1(n9267), .IN2(n1036), .IN3(se_mul), .Q(n9266) );
  NAND2X0 U9516 ( .IN1(n9229), .IN2(n9193), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N39 ) );
  AO221X1 U9517 ( .IN1(n9244), .IN2(n9231), .IN3(n9227), .IN4(n9242), .IN5(
        se_mul), .Q(n9193) );
  AO21X1 U9518 ( .IN1(n9195), .IN2(n1357), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N38 ) );
  INVX0 U9519 ( .INP(n9250), .ZN(n9195) );
  AO22X1 U9520 ( .IN1(n9268), .IN2(n9269), .IN3(\fpu_mul_frac_dp/n838 ), .IN4(
        n9270), .Q(n9250) );
  AO21X1 U9521 ( .IN1(n9196), .IN2(n1358), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N37 ) );
  INVX0 U9522 ( .INP(n9258), .ZN(n9196) );
  AO22X1 U9523 ( .IN1(n9268), .IN2(n9253), .IN3(\fpu_mul_frac_dp/n838 ), .IN4(
        n9271), .Q(n9258) );
  AO21X1 U9524 ( .IN1(n9197), .IN2(n1359), .IN3(n9252), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N36 ) );
  INVX0 U9525 ( .INP(n9229), .ZN(n9252) );
  INVX0 U9526 ( .INP(n9267), .ZN(n9197) );
  AO22X1 U9527 ( .IN1(n9268), .IN2(n9254), .IN3(\fpu_mul_frac_dp/n838 ), .IN4(
        n9272), .Q(n9267) );
  NAND2X0 U9528 ( .IN1(n9229), .IN2(n9198), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N35 ) );
  AO221X1 U9529 ( .IN1(n9273), .IN2(n9231), .IN3(n9227), .IN4(n9274), .IN5(
        se_mul), .Q(n9198) );
  NOR2X0 U9530 ( .IN1(n9176), .IN2(n1033), .QN(n9273) );
  INVX0 U9531 ( .INP(n9275), .ZN(n9176) );
  NAND2X0 U9532 ( .IN1(n9229), .IN2(n9199), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N34 ) );
  AO221X1 U9533 ( .IN1(n9227), .IN2(n9276), .IN3(n9231), .IN4(n9277), .IN5(
        se_mul), .Q(n9199) );
  NAND2X0 U9534 ( .IN1(n9229), .IN2(n9200), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N33 ) );
  AO221X1 U9535 ( .IN1(n9227), .IN2(n9278), .IN3(n9231), .IN4(n9279), .IN5(
        se_mul), .Q(n9200) );
  NAND2X0 U9536 ( .IN1(n9229), .IN2(n9201), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N32 ) );
  AO221X1 U9537 ( .IN1(n9227), .IN2(n9280), .IN3(n9231), .IN4(n9281), .IN5(
        se_mul), .Q(n9201) );
  NAND2X0 U9538 ( .IN1(n9229), .IN2(n9202), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N31 ) );
  AO221X1 U9539 ( .IN1(n9227), .IN2(n9282), .IN3(n9231), .IN4(n9283), .IN5(
        se_mul), .Q(n9202) );
  NAND2X0 U9540 ( .IN1(n9229), .IN2(n9203), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N30 ) );
  AO221X1 U9541 ( .IN1(n9227), .IN2(n9284), .IN3(n9231), .IN4(n9285), .IN5(
        se_mul), .Q(n9203) );
  NAND2X0 U9542 ( .IN1(n9229), .IN2(n9194), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N3 ) );
  NAND4X0 U9543 ( .IN1(n9286), .IN2(n9287), .IN3(n9288), .IN4(n9289), .QN(
        n9194) );
  NOR4X0 U9544 ( .IN1(n9290), .IN2(n9291), .IN3(n9292), .IN4(n9293), .QN(n9289) );
  OR4X1 U9545 ( .IN1(m4stg_frac[40]), .IN2(m4stg_frac[41]), .IN3(
        m4stg_frac[42]), .IN4(m4stg_frac[43]), .Q(n9293) );
  OR4X1 U9546 ( .IN1(m4stg_frac[44]), .IN2(m4stg_frac[45]), .IN3(
        m4stg_frac[46]), .IN4(m4stg_frac[48]), .Q(n9292) );
  OR4X1 U9547 ( .IN1(m4stg_frac[49]), .IN2(m4stg_frac[4]), .IN3(m4stg_frac[50]), .IN4(m4stg_frac[5]), .Q(n9291) );
  OR4X1 U9548 ( .IN1(m4stg_frac[6]), .IN2(m4stg_frac[7]), .IN3(n9294), .IN4(
        m4stg_frac[8]), .Q(n9290) );
  OR2X1 U9549 ( .IN1(se_mul), .IN2(m4stg_frac[9]), .Q(n9294) );
  NOR4X0 U9550 ( .IN1(n9295), .IN2(n9296), .IN3(n9297), .IN4(n9298), .QN(n9288) );
  OR4X1 U9551 ( .IN1(m4stg_frac[21]), .IN2(m4stg_frac[23]), .IN3(
        m4stg_frac[24]), .IN4(m4stg_frac[28]), .Q(n9298) );
  OR4X1 U9552 ( .IN1(m4stg_frac[29]), .IN2(m4stg_frac[2]), .IN3(m4stg_frac[31]), .IN4(m4stg_frac[32]), .Q(n9297) );
  OR4X1 U9553 ( .IN1(m4stg_frac[33]), .IN2(m4stg_frac[34]), .IN3(
        m4stg_frac[35]), .IN4(m4stg_frac[36]), .Q(n9296) );
  OR4X1 U9554 ( .IN1(m4stg_frac[37]), .IN2(m4stg_frac[38]), .IN3(
        m4stg_frac[39]), .IN4(m4stg_frac[3]), .Q(n9295) );
  NOR4X0 U9555 ( .IN1(n9299), .IN2(n9300), .IN3(n9301), .IN4(n9302), .QN(n9287) );
  AO221X1 U9556 ( .IN1(n9187), .IN2(n9303), .IN3(n9304), .IN4(n9305), .IN5(
        n9306), .Q(n9302) );
  AO22X1 U9557 ( .IN1(m4stg_frac[51]), .IN2(n9307), .IN3(m4stg_frac[53]), 
        .IN4(n1411), .Q(n9306) );
  OR4X1 U9558 ( .IN1(n9308), .IN2(n9309), .IN3(n9310), .IN4(n9311), .Q(n9305)
         );
  OR4X1 U9559 ( .IN1(n9312), .IN2(n9313), .IN3(n9314), .IN4(n9315), .Q(n9303)
         );
  OR4X1 U9560 ( .IN1(n9316), .IN2(n9317), .IN3(n9318), .IN4(n9319), .Q(n9315)
         );
  OR4X1 U9561 ( .IN1(n9320), .IN2(n9321), .IN3(n9322), .IN4(n9230), .Q(n9314)
         );
  AO221X1 U9562 ( .IN1(n1378), .IN2(n9323), .IN3(n1364), .IN4(n9324), .IN5(
        n9325), .Q(n9230) );
  AO22X1 U9563 ( .IN1(n1365), .IN2(n9326), .IN3(n1371), .IN4(n9327), .Q(n9325)
         );
  OAI22X1 U9564 ( .IN1(n9328), .IN2(n9246), .IN3(\fpu_mul_frac_dp/n767 ), 
        .IN4(n9329), .QN(n9322) );
  NOR4X0 U9565 ( .IN1(n9330), .IN2(n9331), .IN3(n9332), .IN4(n9333), .QN(n9329) );
  OR4X1 U9566 ( .IN1(n9236), .IN2(n9241), .IN3(n9248), .IN4(n9256), .Q(n9333)
         );
  OR4X1 U9567 ( .IN1(n9265), .IN2(n9334), .IN3(n9335), .IN4(n9336), .Q(n9332)
         );
  OR4X1 U9568 ( .IN1(n9337), .IN2(n9284), .IN3(n9282), .IN4(n9280), .Q(n9331)
         );
  OR4X1 U9569 ( .IN1(n9278), .IN2(n9276), .IN3(n9274), .IN4(n9232), .Q(n9330)
         );
  NAND2X0 U9570 ( .IN1(n1036), .IN2(n908), .QN(n9246) );
  NOR4X0 U9571 ( .IN1(n9338), .IN2(n9339), .IN3(n9340), .IN4(n9341), .QN(n9328) );
  OR3X1 U9572 ( .IN1(n9242), .IN2(n9270), .IN3(n9235), .Q(n9341) );
  OR4X1 U9573 ( .IN1(n9271), .IN2(n9272), .IN3(n9342), .IN4(n9260), .Q(n9340)
         );
  NAND4X0 U9574 ( .IN1(n9262), .IN2(n9185), .IN3(n9184), .IN4(n9183), .QN(
        n9339) );
  INVX0 U9575 ( .INP(n9285), .ZN(n9183) );
  INVX0 U9576 ( .INP(n9343), .ZN(n9184) );
  INVX0 U9577 ( .INP(n9344), .ZN(n9185) );
  INVX0 U9578 ( .INP(n9345), .ZN(n9262) );
  NAND4X0 U9579 ( .IN1(n9182), .IN2(n9181), .IN3(n9179), .IN4(n9178), .QN(
        n9338) );
  INVX0 U9580 ( .INP(n9277), .ZN(n9178) );
  INVX0 U9581 ( .INP(n9279), .ZN(n9179) );
  INVX0 U9582 ( .INP(n9281), .ZN(n9181) );
  INVX0 U9583 ( .INP(n9283), .ZN(n9182) );
  OR4X1 U9584 ( .IN1(n9240), .IN2(n9245), .IN3(n9247), .IN4(n9255), .Q(n9313)
         );
  AO221X1 U9585 ( .IN1(n1366), .IN2(n9327), .IN3(n1363), .IN4(n9326), .IN5(
        n9346), .Q(n9255) );
  AO22X1 U9586 ( .IN1(n1380), .IN2(n9310), .IN3(n1369), .IN4(n9323), .Q(n9346)
         );
  AO221X1 U9587 ( .IN1(m4stg_frac[55]), .IN2(n1411), .IN3(m4stg_frac[54]), 
        .IN4(n1426), .IN5(n9348), .Q(n9310) );
  AO22X1 U9588 ( .IN1(m4stg_frac[53]), .IN2(n1436), .IN3(m4stg_frac[52]), 
        .IN4(n1443), .Q(n9348) );
  AO221X1 U9589 ( .IN1(n1377), .IN2(n9309), .IN3(n1366), .IN4(n9350), .IN5(
        n9351), .Q(n9247) );
  AO22X1 U9590 ( .IN1(n1361), .IN2(n9352), .IN3(n1370), .IN4(n9353), .Q(n9351)
         );
  AO221X1 U9591 ( .IN1(m4stg_frac[56]), .IN2(n1411), .IN3(m4stg_frac[55]), 
        .IN4(n1421), .IN5(n9354), .Q(n9309) );
  AO22X1 U9592 ( .IN1(m4stg_frac[54]), .IN2(n1433), .IN3(m4stg_frac[53]), 
        .IN4(n1439), .Q(n9354) );
  AO221X1 U9593 ( .IN1(n1380), .IN2(n9308), .IN3(n1367), .IN4(n9355), .IN5(
        n9356), .Q(n9245) );
  AO22X1 U9594 ( .IN1(n1364), .IN2(n9357), .IN3(n1372), .IN4(n9358), .Q(n9356)
         );
  AO221X1 U9595 ( .IN1(m4stg_frac[57]), .IN2(n1411), .IN3(m4stg_frac[56]), 
        .IN4(n1421), .IN5(n9359), .Q(n9308) );
  AO22X1 U9596 ( .IN1(m4stg_frac[55]), .IN2(n1432), .IN3(m4stg_frac[54]), 
        .IN4(n1439), .Q(n9359) );
  AO221X1 U9597 ( .IN1(n1379), .IN2(n9360), .IN3(n1361), .IN4(n9361), .IN5(
        n9362), .Q(n9240) );
  AO22X1 U9598 ( .IN1(n1366), .IN2(n9363), .IN3(n1371), .IN4(n9364), .Q(n9362)
         );
  OR4X1 U9599 ( .IN1(n9264), .IN2(n9365), .IN3(n9366), .IN4(n9367), .Q(n9312)
         );
  OR2X1 U9600 ( .IN1(n9368), .IN2(n9369), .Q(n9366) );
  AO221X1 U9601 ( .IN1(n1365), .IN2(n9364), .IN3(n1362), .IN4(n9363), .IN5(
        n9370), .Q(n9264) );
  AO22X1 U9602 ( .IN1(n1378), .IN2(n9311), .IN3(n1369), .IN4(n9360), .Q(n9370)
         );
  AO221X1 U9603 ( .IN1(m4stg_frac[54]), .IN2(n1411), .IN3(m4stg_frac[53]), 
        .IN4(n1421), .IN5(n9371), .Q(n9311) );
  AO22X1 U9604 ( .IN1(m4stg_frac[52]), .IN2(n1432), .IN3(m4stg_frac[51]), 
        .IN4(n1439), .Q(n9371) );
  AO221X1 U9605 ( .IN1(n1362), .IN2(n9372), .IN3(n9373), .IN4(n1033), .IN5(
        n9374), .Q(n9301) );
  OR2X1 U9606 ( .IN1(m4stg_frac[0]), .IN2(m4stg_frac[10]), .Q(n9374) );
  OR4X1 U9607 ( .IN1(n9360), .IN2(n9358), .IN3(n9353), .IN4(n9323), .Q(n9373)
         );
  AO221X1 U9608 ( .IN1(m4stg_frac[59]), .IN2(n1411), .IN3(m4stg_frac[58]), 
        .IN4(n1421), .IN5(n9375), .Q(n9323) );
  AO22X1 U9609 ( .IN1(m4stg_frac[57]), .IN2(n1432), .IN3(m4stg_frac[56]), 
        .IN4(n1439), .Q(n9375) );
  AO221X1 U9610 ( .IN1(m4stg_frac[58]), .IN2(n1411), .IN3(m4stg_frac[57]), 
        .IN4(n1421), .IN5(n9376), .Q(n9360) );
  AO22X1 U9611 ( .IN1(m4stg_frac[56]), .IN2(n1432), .IN3(m4stg_frac[55]), 
        .IN4(n1439), .Q(n9376) );
  OR4X1 U9612 ( .IN1(n9364), .IN2(n9355), .IN3(n9350), .IN4(n9327), .Q(n9372)
         );
  OR4X1 U9613 ( .IN1(m4stg_frac[11]), .IN2(m4stg_frac[12]), .IN3(
        m4stg_frac[15]), .IN4(m4stg_frac[16]), .Q(n9300) );
  OR4X1 U9614 ( .IN1(m4stg_frac[17]), .IN2(m4stg_frac[19]), .IN3(m4stg_frac[1]), .IN4(m4stg_frac[20]), .Q(n9299) );
  NOR4X0 U9615 ( .IN1(n9377), .IN2(n9378), .IN3(n9379), .IN4(n9380), .QN(n9286) );
  OR4X1 U9616 ( .IN1(n9381), .IN2(n9382), .IN3(n9383), .IN4(n9384), .Q(n9380)
         );
  OR4X1 U9617 ( .IN1(n9385), .IN2(n9386), .IN3(n9387), .IN4(n9388), .Q(n9379)
         );
  OR4X1 U9618 ( .IN1(n9389), .IN2(n9390), .IN3(n9391), .IN4(n9392), .Q(n9378)
         );
  OR4X1 U9619 ( .IN1(n9393), .IN2(n9394), .IN3(n9395), .IN4(n9396), .Q(n9377)
         );
  AND2X1 U9620 ( .IN1(m4stg_frac[52]), .IN2(n879), .Q(n9396) );
  NAND2X0 U9621 ( .IN1(n9229), .IN2(n9204), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N29 ) );
  AO221X1 U9622 ( .IN1(n9227), .IN2(n9337), .IN3(n9231), .IN4(n9343), .IN5(
        se_mul), .Q(n9204) );
  NAND2X0 U9623 ( .IN1(n9229), .IN2(n9205), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N28 ) );
  AO221X1 U9624 ( .IN1(n9227), .IN2(n9336), .IN3(n9231), .IN4(n9344), .IN5(
        se_mul), .Q(n9205) );
  NAND2X0 U9625 ( .IN1(n9229), .IN2(n9206), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N27 ) );
  AO221X1 U9626 ( .IN1(n9259), .IN2(n9231), .IN3(n9227), .IN4(n9335), .IN5(
        se_mul), .Q(n9206) );
  NAND2X0 U9627 ( .IN1(n9229), .IN2(n9207), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N26 ) );
  AO221X1 U9628 ( .IN1(n9231), .IN2(n9260), .IN3(n9227), .IN4(n9334), .IN5(
        n9397), .Q(n9207) );
  AO21X1 U9629 ( .IN1(n9398), .IN2(n9399), .IN3(se_mul), .Q(n9397) );
  NAND2X0 U9630 ( .IN1(n9229), .IN2(n9208), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N25 ) );
  AO221X1 U9631 ( .IN1(n9231), .IN2(n9345), .IN3(n9227), .IN4(n9232), .IN5(
        n9400), .Q(n9208) );
  NAND2X0 U9632 ( .IN1(n9401), .IN2(n1358), .QN(n9400) );
  NAND3X0 U9633 ( .IN1(n9234), .IN2(n1377), .IN3(n9263), .QN(n9401) );
  AO221X1 U9634 ( .IN1(n1378), .IN2(n9402), .IN3(n1368), .IN4(n9403), .IN5(
        n9404), .Q(n9232) );
  AO22X1 U9635 ( .IN1(n1362), .IN2(n9405), .IN3(n1370), .IN4(n9406), .Q(n9404)
         );
  AO221X1 U9636 ( .IN1(n1377), .IN2(n9407), .IN3(n1370), .IN4(n9408), .IN5(
        n9409), .Q(n9345) );
  AO22X1 U9637 ( .IN1(n1363), .IN2(n9410), .IN3(n1366), .IN4(n9411), .Q(n9409)
         );
  NAND2X0 U9638 ( .IN1(n9229), .IN2(n9209), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N24 ) );
  AO221X1 U9639 ( .IN1(n9231), .IN2(n9235), .IN3(n9227), .IN4(n9236), .IN5(
        n9412), .Q(n9209) );
  AO21X1 U9640 ( .IN1(n9234), .IN2(n9238), .IN3(se_mul), .Q(n9412) );
  AND2X1 U9641 ( .IN1(n1380), .IN2(n9413), .Q(n9238) );
  AO221X1 U9642 ( .IN1(n1380), .IN2(n9414), .IN3(n1364), .IN4(n9415), .IN5(
        n9416), .Q(n9236) );
  AO22X1 U9643 ( .IN1(n1367), .IN2(n9417), .IN3(n1372), .IN4(n9418), .Q(n9416)
         );
  AO221X1 U9644 ( .IN1(n1368), .IN2(n9419), .IN3(n1363), .IN4(n9420), .IN5(
        n9421), .Q(n9235) );
  AO22X1 U9645 ( .IN1(n1369), .IN2(n9422), .IN3(n1377), .IN4(n9423), .Q(n9421)
         );
  NAND2X0 U9646 ( .IN1(n9229), .IN2(n9210), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N23 ) );
  AO221X1 U9647 ( .IN1(n9227), .IN2(n9241), .IN3(n9231), .IN4(n9242), .IN5(
        n9424), .Q(n9210) );
  AO21X1 U9648 ( .IN1(n9244), .IN2(n9234), .IN3(se_mul), .Q(n9424) );
  NOR2X0 U9649 ( .IN1(n9425), .IN2(n9304), .QN(n9244) );
  AO221X1 U9650 ( .IN1(n1369), .IN2(n9426), .IN3(n1379), .IN4(n9427), .IN5(
        n9428), .Q(n9242) );
  AO22X1 U9651 ( .IN1(n1368), .IN2(n9429), .IN3(n1362), .IN4(n9430), .Q(n9428)
         );
  AO221X1 U9652 ( .IN1(n1379), .IN2(n9431), .IN3(n1361), .IN4(n9432), .IN5(
        n9433), .Q(n9241) );
  AO22X1 U9653 ( .IN1(n1365), .IN2(n9434), .IN3(n1371), .IN4(n9435), .Q(n9433)
         );
  NAND2X0 U9654 ( .IN1(n9229), .IN2(n9211), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N22 ) );
  AO221X1 U9655 ( .IN1(n9231), .IN2(n9270), .IN3(n9398), .IN4(n9269), .IN5(
        n9436), .Q(n9211) );
  AO21X1 U9656 ( .IN1(n9227), .IN2(n9248), .IN3(se_mul), .Q(n9436) );
  AO221X1 U9657 ( .IN1(n1378), .IN2(n9437), .IN3(n1362), .IN4(n9438), .IN5(
        n9439), .Q(n9248) );
  AO22X1 U9658 ( .IN1(n1366), .IN2(n9440), .IN3(n1369), .IN4(n9441), .Q(n9439)
         );
  AO221X1 U9659 ( .IN1(n1367), .IN2(n9442), .IN3(n1377), .IN4(n9443), .IN5(
        n9444), .Q(n9270) );
  AO22X1 U9660 ( .IN1(n1370), .IN2(n9445), .IN3(n1364), .IN4(n9446), .Q(n9444)
         );
  NAND2X0 U9661 ( .IN1(n9229), .IN2(n9212), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N21 ) );
  AO221X1 U9662 ( .IN1(n9231), .IN2(n9271), .IN3(n9398), .IN4(n9253), .IN5(
        n9447), .Q(n9212) );
  AO21X1 U9663 ( .IN1(n9227), .IN2(n9256), .IN3(se_mul), .Q(n9447) );
  AO221X1 U9664 ( .IN1(n1372), .IN2(n9402), .IN3(n1378), .IN4(n9324), .IN5(
        n9448), .Q(n9256) );
  AO22X1 U9665 ( .IN1(n1367), .IN2(n9406), .IN3(n1363), .IN4(n9403), .Q(n9448)
         );
  AO221X1 U9666 ( .IN1(n1366), .IN2(n9408), .IN3(n1364), .IN4(n9411), .IN5(
        n9449), .Q(n9271) );
  AO22X1 U9667 ( .IN1(n1371), .IN2(n9407), .IN3(n1378), .IN4(n9405), .Q(n9449)
         );
  NAND2X0 U9668 ( .IN1(n9229), .IN2(n9213), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N20 ) );
  AO221X1 U9669 ( .IN1(n9231), .IN2(n9272), .IN3(n9398), .IN4(n9254), .IN5(
        n9450), .Q(n9213) );
  AO21X1 U9670 ( .IN1(n9227), .IN2(n9265), .IN3(se_mul), .Q(n9450) );
  AO221X1 U9671 ( .IN1(n1371), .IN2(n9414), .IN3(n1380), .IN4(n9361), .IN5(
        n9451), .Q(n9265) );
  AO22X1 U9672 ( .IN1(n1361), .IN2(n9417), .IN3(n1367), .IN4(n9418), .Q(n9451)
         );
  AO221X1 U9673 ( .IN1(n1365), .IN2(n9422), .IN3(n1363), .IN4(n9419), .IN5(
        n9452), .Q(n9272) );
  AO22X1 U9674 ( .IN1(n1377), .IN2(n9415), .IN3(n1370), .IN4(n9423), .Q(n9452)
         );
  NAND2X0 U9675 ( .IN1(n9229), .IN2(n9214), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N19 ) );
  AO221X1 U9676 ( .IN1(n9227), .IN2(n9321), .IN3(n9231), .IN4(n9274), .IN5(
        n9453), .Q(n9214) );
  AO21X1 U9677 ( .IN1(n9398), .IN2(n9275), .IN3(se_mul), .Q(n9453) );
  AND2X1 U9678 ( .IN1(n9234), .IN2(\fpu_mul_frac_dp/n765 ), .Q(n9398) );
  AO222X1 U9679 ( .IN1(n1369), .IN2(n9427), .IN3(n9454), .IN4(n1033), .IN5(
        n1380), .IN6(n9432), .Q(n9274) );
  AO221X1 U9680 ( .IN1(n1377), .IN2(n9357), .IN3(n1372), .IN4(n9431), .IN5(
        n9455), .Q(n9321) );
  AO22X1 U9681 ( .IN1(n1364), .IN2(n9434), .IN3(n1368), .IN4(n9435), .Q(n9455)
         );
  NAND2X0 U9682 ( .IN1(n9229), .IN2(n9215), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N18 ) );
  AO221X1 U9683 ( .IN1(n9231), .IN2(n9276), .IN3(n9234), .IN4(n9277), .IN5(
        n9456), .Q(n9215) );
  AO21X1 U9684 ( .IN1(n9227), .IN2(n9320), .IN3(se_mul), .Q(n9456) );
  AO221X1 U9685 ( .IN1(n1380), .IN2(n9352), .IN3(n1371), .IN4(n9437), .IN5(
        n9457), .Q(n9320) );
  AO22X1 U9686 ( .IN1(n1362), .IN2(n9440), .IN3(n1365), .IN4(n9441), .Q(n9457)
         );
  AO222X1 U9687 ( .IN1(n1379), .IN2(n9446), .IN3(n1370), .IN4(n9458), .IN5(
        n9399), .IN6(n1033), .Q(n9277) );
  INVX0 U9688 ( .INP(n9459), .ZN(n9399) );
  AO221X1 U9689 ( .IN1(n1370), .IN2(n9443), .IN3(n1379), .IN4(n9438), .IN5(
        n9460), .Q(n9276) );
  AO22X1 U9690 ( .IN1(n1363), .IN2(n9442), .IN3(n1366), .IN4(n9445), .Q(n9460)
         );
  NAND2X0 U9691 ( .IN1(n9229), .IN2(n9216), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N17 ) );
  AO221X1 U9692 ( .IN1(n9231), .IN2(n9278), .IN3(n9234), .IN4(n9279), .IN5(
        n9461), .Q(n9216) );
  AO21X1 U9693 ( .IN1(n9227), .IN2(n9319), .IN3(se_mul), .Q(n9461) );
  AO221X1 U9694 ( .IN1(n1379), .IN2(n9326), .IN3(n1361), .IN4(n9406), .IN5(
        n9462), .Q(n9319) );
  AO22X1 U9695 ( .IN1(n1372), .IN2(n9324), .IN3(n1367), .IN4(n9402), .Q(n9462)
         );
  AO222X1 U9696 ( .IN1(n1377), .IN2(n9411), .IN3(n9263), .IN4(n1367), .IN5(
        n1372), .IN6(n9410), .Q(n9279) );
  AO221X1 U9697 ( .IN1(n1378), .IN2(n9403), .IN3(n1369), .IN4(n9405), .IN5(
        n9463), .Q(n9278) );
  AO22X1 U9698 ( .IN1(n1361), .IN2(n9408), .IN3(n1368), .IN4(n9407), .Q(n9463)
         );
  NAND2X0 U9699 ( .IN1(n9229), .IN2(n9217), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N16 ) );
  AO221X1 U9700 ( .IN1(n9231), .IN2(n9280), .IN3(n9234), .IN4(n9281), .IN5(
        n9464), .Q(n9217) );
  AO21X1 U9701 ( .IN1(n9227), .IN2(n9318), .IN3(se_mul), .Q(n9464) );
  AO221X1 U9702 ( .IN1(n1377), .IN2(n9363), .IN3(n1362), .IN4(n9418), .IN5(
        n9465), .Q(n9318) );
  AO22X1 U9703 ( .IN1(n1369), .IN2(n9361), .IN3(n1365), .IN4(n9414), .Q(n9465)
         );
  AO222X1 U9704 ( .IN1(n1366), .IN2(n9413), .IN3(n1379), .IN4(n9419), .IN5(
        n1371), .IN6(n9420), .Q(n9281) );
  AO221X1 U9705 ( .IN1(n1380), .IN2(n9417), .IN3(n1364), .IN4(n9422), .IN5(
        n9466), .Q(n9280) );
  AO22X1 U9706 ( .IN1(n1370), .IN2(n9415), .IN3(n1366), .IN4(n9423), .Q(n9466)
         );
  NAND2X0 U9707 ( .IN1(n9229), .IN2(n9218), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N15 ) );
  AO221X1 U9708 ( .IN1(n9231), .IN2(n9282), .IN3(n9234), .IN4(n9283), .IN5(
        n9467), .Q(n9218) );
  AO21X1 U9709 ( .IN1(n9227), .IN2(n9317), .IN3(se_mul), .Q(n9467) );
  AO221X1 U9710 ( .IN1(n1379), .IN2(n9355), .IN3(n1370), .IN4(n9357), .IN5(
        n9468), .Q(n9317) );
  AO22X1 U9711 ( .IN1(n1364), .IN2(n9435), .IN3(n1367), .IN4(n9431), .Q(n9468)
         );
  AO222X1 U9712 ( .IN1(n1370), .IN2(n9430), .IN3(n9469), .IN4(n1366), .IN5(
        n1377), .IN6(n9429), .Q(n9283) );
  AO221X1 U9713 ( .IN1(n1361), .IN2(n9426), .IN3(n1365), .IN4(n9427), .IN5(
        n9470), .Q(n9282) );
  AO22X1 U9714 ( .IN1(n1379), .IN2(n9434), .IN3(n1372), .IN4(n9432), .Q(n9470)
         );
  NAND2X0 U9715 ( .IN1(n9229), .IN2(n9219), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N14 ) );
  AO221X1 U9716 ( .IN1(n9231), .IN2(n9284), .IN3(n9234), .IN4(n9285), .IN5(
        n9471), .Q(n9219) );
  AO21X1 U9717 ( .IN1(n9227), .IN2(n9316), .IN3(se_mul), .Q(n9471) );
  AO221X1 U9718 ( .IN1(n1378), .IN2(n9350), .IN3(n1372), .IN4(n9352), .IN5(
        n9472), .Q(n9316) );
  AO22X1 U9719 ( .IN1(n1362), .IN2(n9441), .IN3(n1368), .IN4(n9437), .Q(n9472)
         );
  AO222X1 U9720 ( .IN1(n1371), .IN2(n9446), .IN3(n9269), .IN4(n1033), .IN5(
        n1379), .IN6(n9442), .Q(n9285) );
  INVX0 U9721 ( .INP(n9172), .ZN(n9269) );
  MUX21X1 U9722 ( .IN1(n9473), .IN2(n9474), .S(\fpu_mul_frac_dp/n833 ), .Q(
        n9172) );
  INVX0 U9723 ( .INP(n9458), .ZN(n9474) );
  NAND2X0 U9724 ( .IN1(m4stg_frac_105), .IN2(n1447), .QN(n9473) );
  AO221X1 U9725 ( .IN1(n1369), .IN2(n9438), .IN3(n1377), .IN4(n9440), .IN5(
        n9475), .Q(n9284) );
  AO22X1 U9726 ( .IN1(n1368), .IN2(n9443), .IN3(n1361), .IN4(n9445), .Q(n9475)
         );
  NAND2X0 U9727 ( .IN1(n9229), .IN2(n9220), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N13 ) );
  AO221X1 U9728 ( .IN1(n9231), .IN2(n9337), .IN3(n9234), .IN4(n9343), .IN5(
        n9476), .Q(n9220) );
  AO21X1 U9729 ( .IN1(n9227), .IN2(n9368), .IN3(se_mul), .Q(n9476) );
  AO221X1 U9730 ( .IN1(n1377), .IN2(n9327), .IN3(n1371), .IN4(n9326), .IN5(
        n9477), .Q(n9368) );
  AO22X1 U9731 ( .IN1(n1365), .IN2(n9324), .IN3(n1362), .IN4(n9402), .Q(n9477)
         );
  AO221X1 U9732 ( .IN1(m4stg_frac[75]), .IN2(n1411), .IN3(m4stg_frac[74]), 
        .IN4(n1421), .IN5(n9478), .Q(n9402) );
  AO22X1 U9733 ( .IN1(m4stg_frac[73]), .IN2(n1433), .IN3(m4stg_frac[72]), 
        .IN4(n1439), .Q(n9478) );
  AO221X1 U9734 ( .IN1(m4stg_frac[71]), .IN2(n1411), .IN3(m4stg_frac[70]), 
        .IN4(n1421), .IN5(n9479), .Q(n9324) );
  AO22X1 U9735 ( .IN1(m4stg_frac[69]), .IN2(n1432), .IN3(m4stg_frac[68]), 
        .IN4(n1439), .Q(n9479) );
  AO221X1 U9736 ( .IN1(m4stg_frac[67]), .IN2(n1411), .IN3(m4stg_frac[66]), 
        .IN4(n1421), .IN5(n9480), .Q(n9326) );
  AO22X1 U9737 ( .IN1(m4stg_frac[65]), .IN2(n1432), .IN3(m4stg_frac[64]), 
        .IN4(n1439), .Q(n9480) );
  AO221X1 U9738 ( .IN1(m4stg_frac[63]), .IN2(n1412), .IN3(m4stg_frac[62]), 
        .IN4(n1421), .IN5(n9481), .Q(n9327) );
  AO22X1 U9739 ( .IN1(m4stg_frac[61]), .IN2(n1432), .IN3(m4stg_frac[60]), 
        .IN4(n1439), .Q(n9481) );
  AO222X1 U9740 ( .IN1(n1372), .IN2(n9411), .IN3(n1378), .IN4(n9408), .IN5(
        n9253), .IN6(n1033), .Q(n9343) );
  MUX21X1 U9741 ( .IN1(n9263), .IN2(n9410), .S(\fpu_mul_frac_dp/n833 ), .Q(
        n9253) );
  AO221X1 U9742 ( .IN1(m4stg_frac[103]), .IN2(n1411), .IN3(m4stg_frac[102]), 
        .IN4(n1421), .IN5(n9482), .Q(n9410) );
  AO22X1 U9743 ( .IN1(m4stg_frac[101]), .IN2(n1433), .IN3(m4stg_frac[100]), 
        .IN4(n1439), .Q(n9482) );
  NOR2X0 U9744 ( .IN1(n9251), .IN2(n879), .QN(n9263) );
  AO221X1 U9745 ( .IN1(m4stg_frac[95]), .IN2(n1412), .IN3(n1430), .IN4(
        m4stg_frac[94]), .IN5(n9483), .Q(n9408) );
  AO22X1 U9746 ( .IN1(m4stg_frac[93]), .IN2(n1432), .IN3(m4stg_frac[92]), 
        .IN4(n1439), .Q(n9483) );
  AO221X1 U9747 ( .IN1(m4stg_frac[99]), .IN2(n1412), .IN3(m4stg_frac[98]), 
        .IN4(n1421), .IN5(n9484), .Q(n9411) );
  AO22X1 U9748 ( .IN1(m4stg_frac[97]), .IN2(n1433), .IN3(m4stg_frac[96]), 
        .IN4(n1439), .Q(n9484) );
  AO221X1 U9749 ( .IN1(n1372), .IN2(n9403), .IN3(n1378), .IN4(n9406), .IN5(
        n9485), .Q(n9337) );
  AO22X1 U9750 ( .IN1(n1363), .IN2(n9407), .IN3(n1365), .IN4(n9405), .Q(n9485)
         );
  AO221X1 U9751 ( .IN1(m4stg_frac[87]), .IN2(n1412), .IN3(m4stg_frac[86]), 
        .IN4(n1422), .IN5(n9486), .Q(n9405) );
  AO22X1 U9752 ( .IN1(m4stg_frac[85]), .IN2(n1433), .IN3(m4stg_frac[84]), 
        .IN4(n1439), .Q(n9486) );
  AO221X1 U9753 ( .IN1(m4stg_frac[91]), .IN2(n1412), .IN3(m4stg_frac[88]), 
        .IN4(n1439), .IN5(n9487), .Q(n9407) );
  NAND2X0 U9754 ( .IN1(n9488), .IN2(n9489), .QN(n9487) );
  AO221X1 U9755 ( .IN1(m4stg_frac[79]), .IN2(n1412), .IN3(m4stg_frac[78]), 
        .IN4(n1422), .IN5(n9490), .Q(n9406) );
  AO22X1 U9756 ( .IN1(m4stg_frac[77]), .IN2(n1432), .IN3(m4stg_frac[76]), 
        .IN4(n1440), .Q(n9490) );
  AO221X1 U9757 ( .IN1(m4stg_frac[83]), .IN2(n1412), .IN3(m4stg_frac[82]), 
        .IN4(n1422), .IN5(n9491), .Q(n9403) );
  AO22X1 U9758 ( .IN1(m4stg_frac[81]), .IN2(n1433), .IN3(m4stg_frac[80]), 
        .IN4(n1440), .Q(n9491) );
  NAND2X0 U9759 ( .IN1(n9229), .IN2(n9221), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N12 ) );
  AO221X1 U9760 ( .IN1(n9231), .IN2(n9336), .IN3(n9234), .IN4(n9344), .IN5(
        n9492), .Q(n9221) );
  AO21X1 U9761 ( .IN1(n9227), .IN2(n9369), .IN3(se_mul), .Q(n9492) );
  AO221X1 U9762 ( .IN1(n1380), .IN2(n9364), .IN3(n1369), .IN4(n9363), .IN5(
        n9493), .Q(n9369) );
  AO22X1 U9763 ( .IN1(n1366), .IN2(n9361), .IN3(n1364), .IN4(n9414), .Q(n9493)
         );
  AO221X1 U9764 ( .IN1(m4stg_frac[74]), .IN2(n1412), .IN3(m4stg_frac[73]), 
        .IN4(n1422), .IN5(n9494), .Q(n9414) );
  AO22X1 U9765 ( .IN1(m4stg_frac[72]), .IN2(n1432), .IN3(m4stg_frac[71]), 
        .IN4(n1440), .Q(n9494) );
  AO221X1 U9766 ( .IN1(m4stg_frac[70]), .IN2(n1412), .IN3(m4stg_frac[69]), 
        .IN4(n1422), .IN5(n9495), .Q(n9361) );
  AO22X1 U9767 ( .IN1(m4stg_frac[68]), .IN2(n1433), .IN3(m4stg_frac[67]), 
        .IN4(n1440), .Q(n9495) );
  AO221X1 U9768 ( .IN1(m4stg_frac[66]), .IN2(n1412), .IN3(m4stg_frac[65]), 
        .IN4(n1422), .IN5(n9496), .Q(n9363) );
  AO22X1 U9769 ( .IN1(m4stg_frac[64]), .IN2(n1433), .IN3(m4stg_frac[63]), 
        .IN4(n1440), .Q(n9496) );
  AO221X1 U9770 ( .IN1(m4stg_frac[62]), .IN2(n1412), .IN3(m4stg_frac[61]), 
        .IN4(n1422), .IN5(n9497), .Q(n9364) );
  AO22X1 U9771 ( .IN1(m4stg_frac[60]), .IN2(n1433), .IN3(m4stg_frac[59]), 
        .IN4(n1440), .Q(n9497) );
  AO222X1 U9772 ( .IN1(n1369), .IN2(n9419), .IN3(n1380), .IN4(n9422), .IN5(
        n9254), .IN6(n1033), .Q(n9344) );
  MUX21X1 U9773 ( .IN1(n9413), .IN2(n9420), .S(\fpu_mul_frac_dp/n833 ), .Q(
        n9254) );
  AO221X1 U9774 ( .IN1(m4stg_frac[102]), .IN2(n1412), .IN3(m4stg_frac[101]), 
        .IN4(n1422), .IN5(n9498), .Q(n9420) );
  AO22X1 U9775 ( .IN1(m4stg_frac[100]), .IN2(n1433), .IN3(m4stg_frac[99]), 
        .IN4(n1440), .Q(n9498) );
  AO222X1 U9776 ( .IN1(m4stg_frac[103]), .IN2(n1446), .IN3(m4stg_frac_105), 
        .IN4(n1423), .IN5(m4stg_frac[104]), .IN6(n1431), .Q(n9413) );
  AO221X1 U9777 ( .IN1(m4stg_frac[94]), .IN2(n1412), .IN3(m4stg_frac[93]), 
        .IN4(n1422), .IN5(n9499), .Q(n9422) );
  AO22X1 U9778 ( .IN1(m4stg_frac[92]), .IN2(n1433), .IN3(m4stg_frac[91]), 
        .IN4(n1440), .Q(n9499) );
  AO221X1 U9779 ( .IN1(m4stg_frac[98]), .IN2(n1412), .IN3(m4stg_frac[97]), 
        .IN4(n1422), .IN5(n9500), .Q(n9419) );
  AO22X1 U9780 ( .IN1(m4stg_frac[96]), .IN2(n1434), .IN3(n1446), .IN4(
        m4stg_frac[95]), .Q(n9500) );
  AO221X1 U9781 ( .IN1(n1379), .IN2(n9418), .IN3(n1370), .IN4(n9417), .IN5(
        n9501), .Q(n9336) );
  AO22X1 U9782 ( .IN1(n1367), .IN2(n9415), .IN3(n1363), .IN4(n9423), .Q(n9501)
         );
  AO221X1 U9783 ( .IN1(m4stg_frac[90]), .IN2(n1413), .IN3(m4stg_frac[89]), 
        .IN4(n1422), .IN5(n9502), .Q(n9423) );
  AO22X1 U9784 ( .IN1(m4stg_frac[88]), .IN2(n1433), .IN3(m4stg_frac[87]), 
        .IN4(n1440), .Q(n9502) );
  AO221X1 U9785 ( .IN1(m4stg_frac[86]), .IN2(n1413), .IN3(m4stg_frac[85]), 
        .IN4(n1422), .IN5(n9503), .Q(n9415) );
  AO22X1 U9786 ( .IN1(m4stg_frac[84]), .IN2(n1434), .IN3(m4stg_frac[83]), 
        .IN4(n1440), .Q(n9503) );
  AO221X1 U9787 ( .IN1(m4stg_frac[82]), .IN2(n1413), .IN3(m4stg_frac[81]), 
        .IN4(n1423), .IN5(n9504), .Q(n9417) );
  AO22X1 U9788 ( .IN1(m4stg_frac[80]), .IN2(n1433), .IN3(m4stg_frac[79]), 
        .IN4(n1440), .Q(n9504) );
  AO221X1 U9789 ( .IN1(m4stg_frac[78]), .IN2(n1413), .IN3(m4stg_frac[77]), 
        .IN4(n1423), .IN5(n9505), .Q(n9418) );
  AO22X1 U9790 ( .IN1(m4stg_frac[76]), .IN2(n1433), .IN3(m4stg_frac[75]), 
        .IN4(n1440), .Q(n9505) );
  NAND2X0 U9791 ( .IN1(n9229), .IN2(n9222), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N11 ) );
  AO221X1 U9792 ( .IN1(n9259), .IN2(n9234), .IN3(n9231), .IN4(n9335), .IN5(
        n9506), .Q(n9222) );
  AO21X1 U9793 ( .IN1(n9227), .IN2(n9367), .IN3(se_mul), .Q(n9506) );
  AO221X1 U9794 ( .IN1(n1368), .IN2(n9357), .IN3(n1363), .IN4(n9431), .IN5(
        n9507), .Q(n9367) );
  AO22X1 U9795 ( .IN1(n1380), .IN2(n9358), .IN3(n1371), .IN4(n9355), .Q(n9507)
         );
  AO221X1 U9796 ( .IN1(m4stg_frac[65]), .IN2(n1413), .IN3(m4stg_frac[64]), 
        .IN4(n1423), .IN5(n9508), .Q(n9355) );
  AO22X1 U9797 ( .IN1(m4stg_frac[63]), .IN2(n1434), .IN3(m4stg_frac[62]), 
        .IN4(n1440), .Q(n9508) );
  AO221X1 U9798 ( .IN1(m4stg_frac[61]), .IN2(n1413), .IN3(m4stg_frac[60]), 
        .IN4(n1423), .IN5(n9509), .Q(n9358) );
  AO22X1 U9799 ( .IN1(m4stg_frac[59]), .IN2(n1433), .IN3(m4stg_frac[58]), 
        .IN4(n1440), .Q(n9509) );
  AO221X1 U9800 ( .IN1(m4stg_frac[73]), .IN2(n1413), .IN3(m4stg_frac[72]), 
        .IN4(n1423), .IN5(n9510), .Q(n9431) );
  AO22X1 U9801 ( .IN1(m4stg_frac[71]), .IN2(n1434), .IN3(m4stg_frac[70]), 
        .IN4(n1440), .Q(n9510) );
  AO221X1 U9802 ( .IN1(m4stg_frac[69]), .IN2(n1413), .IN3(m4stg_frac[68]), 
        .IN4(n1423), .IN5(n9511), .Q(n9357) );
  AO22X1 U9803 ( .IN1(m4stg_frac[67]), .IN2(n1434), .IN3(m4stg_frac[66]), 
        .IN4(n1440), .Q(n9511) );
  AO221X1 U9804 ( .IN1(n1364), .IN2(n9427), .IN3(n1366), .IN4(n9432), .IN5(
        n9512), .Q(n9335) );
  AO22X1 U9805 ( .IN1(n1371), .IN2(n9434), .IN3(n1380), .IN4(n9435), .Q(n9512)
         );
  AO221X1 U9806 ( .IN1(m4stg_frac[77]), .IN2(n1413), .IN3(m4stg_frac[76]), 
        .IN4(n1423), .IN5(n9513), .Q(n9435) );
  AO22X1 U9807 ( .IN1(m4stg_frac[75]), .IN2(n1434), .IN3(m4stg_frac[74]), 
        .IN4(n1441), .Q(n9513) );
  AO221X1 U9808 ( .IN1(m4stg_frac[81]), .IN2(n1415), .IN3(m4stg_frac[80]), 
        .IN4(n1423), .IN5(n9514), .Q(n9434) );
  AO22X1 U9809 ( .IN1(m4stg_frac[79]), .IN2(n1434), .IN3(m4stg_frac[78]), 
        .IN4(n1441), .Q(n9514) );
  AO221X1 U9810 ( .IN1(m4stg_frac[85]), .IN2(n1413), .IN3(m4stg_frac[84]), 
        .IN4(n1423), .IN5(n9515), .Q(n9432) );
  AO22X1 U9811 ( .IN1(m4stg_frac[83]), .IN2(n1434), .IN3(m4stg_frac[82]), 
        .IN4(n1441), .Q(n9515) );
  AO221X1 U9812 ( .IN1(m4stg_frac[86]), .IN2(n1446), .IN3(m4stg_frac[87]), 
        .IN4(n1431), .IN5(n9516), .Q(n9427) );
  AO21X1 U9813 ( .IN1(m4stg_frac[88]), .IN2(n9347), .IN3(n9517), .Q(n9516) );
  INVX0 U9814 ( .INP(n9518), .ZN(n9517) );
  OA21X1 U9815 ( .IN1(n9454), .IN2(n1033), .IN3(n9342), .Q(n9259) );
  AO21X1 U9816 ( .IN1(\fpu_mul_frac_dp/n765 ), .IN2(n9454), .IN3(n9275), .Q(
        n9342) );
  MUX21X1 U9817 ( .IN1(n9469), .IN2(n9430), .S(\fpu_mul_frac_dp/n833 ), .Q(
        n9275) );
  AO221X1 U9818 ( .IN1(m4stg_frac[101]), .IN2(n1413), .IN3(m4stg_frac[100]), 
        .IN4(n1423), .IN5(n9519), .Q(n9430) );
  AO22X1 U9819 ( .IN1(m4stg_frac[99]), .IN2(n1434), .IN3(m4stg_frac[98]), 
        .IN4(n1441), .Q(n9519) );
  INVX0 U9820 ( .INP(n9425), .ZN(n9469) );
  AO22X1 U9821 ( .IN1(n9520), .IN2(n9521), .IN3(n9251), .IN4(n879), .Q(n9425)
         );
  MUX21X1 U9822 ( .IN1(n1230), .IN2(n979), .S(n884), .Q(n9251) );
  NAND2X0 U9823 ( .IN1(m4stg_frac[102]), .IN2(\fpu_mul_frac_dp/n831 ), .QN(
        n9521) );
  MUX21X1 U9824 ( .IN1(n9429), .IN2(n9426), .S(\fpu_mul_frac_dp/n833 ), .Q(
        n9454) );
  AO221X1 U9825 ( .IN1(m4stg_frac[92]), .IN2(n9347), .IN3(m4stg_frac[91]), 
        .IN4(n1431), .IN5(n9522), .Q(n9426) );
  AO21X1 U9826 ( .IN1(m4stg_frac[93]), .IN2(n1419), .IN3(n9523), .Q(n9522) );
  INVX0 U9827 ( .INP(n9524), .ZN(n9523) );
  AO221X1 U9828 ( .IN1(m4stg_frac[97]), .IN2(n1413), .IN3(m4stg_frac[96]), 
        .IN4(n1423), .IN5(n9525), .Q(n9429) );
  AO22X1 U9829 ( .IN1(m4stg_frac[95]), .IN2(n1434), .IN3(n1446), .IN4(
        m4stg_frac[94]), .Q(n9525) );
  NAND2X0 U9830 ( .IN1(n9229), .IN2(n9223), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre3/N10 ) );
  AO221X1 U9831 ( .IN1(n9227), .IN2(n9365), .IN3(n9231), .IN4(n9334), .IN5(
        n9526), .Q(n9223) );
  AO221X1 U9832 ( .IN1(n9527), .IN2(n9268), .IN3(n9234), .IN4(n9260), .IN5(
        se_mul), .Q(n9526) );
  AO221X1 U9833 ( .IN1(n1378), .IN2(n9445), .IN3(n1372), .IN4(n9442), .IN5(
        n9528), .Q(n9260) );
  AO22X1 U9834 ( .IN1(n1368), .IN2(n9446), .IN3(n1361), .IN4(n9458), .Q(n9528)
         );
  AO221X1 U9835 ( .IN1(n1411), .IN2(m4stg_frac[104]), .IN3(m4stg_frac[103]), 
        .IN4(n1423), .IN5(n9529), .Q(n9458) );
  AO22X1 U9836 ( .IN1(m4stg_frac[102]), .IN2(n1434), .IN3(m4stg_frac[101]), 
        .IN4(n1441), .Q(n9529) );
  AO221X1 U9837 ( .IN1(m4stg_frac[100]), .IN2(n1413), .IN3(m4stg_frac[99]), 
        .IN4(n1424), .IN5(n9530), .Q(n9446) );
  AO22X1 U9838 ( .IN1(m4stg_frac[98]), .IN2(n1434), .IN3(m4stg_frac[97]), 
        .IN4(n1441), .Q(n9530) );
  AO221X1 U9839 ( .IN1(m4stg_frac[96]), .IN2(n1414), .IN3(m4stg_frac[95]), 
        .IN4(n1424), .IN5(n9531), .Q(n9442) );
  AO22X1 U9840 ( .IN1(m4stg_frac[94]), .IN2(n1434), .IN3(m4stg_frac[93]), 
        .IN4(n1441), .Q(n9531) );
  AO221X1 U9841 ( .IN1(m4stg_frac[92]), .IN2(n1413), .IN3(m4stg_frac[91]), 
        .IN4(n1424), .IN5(n9532), .Q(n9445) );
  AO22X1 U9842 ( .IN1(m4stg_frac[90]), .IN2(n1434), .IN3(m4stg_frac[89]), 
        .IN4(n1441), .Q(n9532) );
  NOR2X0 U9843 ( .IN1(n908), .IN2(\fpu_mul_frac_dp/n767 ), .QN(n9234) );
  NOR2X0 U9844 ( .IN1(\fpu_mul_frac_dp/n767 ), .IN2(n9459), .QN(n9527) );
  AO221X1 U9845 ( .IN1(n1377), .IN2(n9441), .IN3(n1371), .IN4(n9440), .IN5(
        n9533), .Q(n9334) );
  AO22X1 U9846 ( .IN1(n1365), .IN2(n9438), .IN3(n1362), .IN4(n9443), .Q(n9533)
         );
  AO221X1 U9847 ( .IN1(m4stg_frac[88]), .IN2(n1414), .IN3(m4stg_frac[87]), 
        .IN4(n1424), .IN5(n9534), .Q(n9443) );
  AO22X1 U9848 ( .IN1(m4stg_frac[86]), .IN2(n1434), .IN3(m4stg_frac[85]), 
        .IN4(n1441), .Q(n9534) );
  AO221X1 U9849 ( .IN1(m4stg_frac[84]), .IN2(n1414), .IN3(m4stg_frac[83]), 
        .IN4(n1424), .IN5(n9535), .Q(n9438) );
  AO22X1 U9850 ( .IN1(m4stg_frac[82]), .IN2(n1435), .IN3(m4stg_frac[81]), 
        .IN4(n1441), .Q(n9535) );
  AO221X1 U9851 ( .IN1(m4stg_frac[80]), .IN2(n1414), .IN3(m4stg_frac[79]), 
        .IN4(n1424), .IN5(n9536), .Q(n9440) );
  AO22X1 U9852 ( .IN1(m4stg_frac[78]), .IN2(n1435), .IN3(m4stg_frac[77]), 
        .IN4(n1441), .Q(n9536) );
  AO221X1 U9853 ( .IN1(m4stg_frac[76]), .IN2(n1414), .IN3(m4stg_frac[75]), 
        .IN4(n1424), .IN5(n9537), .Q(n9441) );
  AO22X1 U9854 ( .IN1(m4stg_frac[74]), .IN2(n1435), .IN3(m4stg_frac[73]), 
        .IN4(n1441), .Q(n9537) );
  NOR2X0 U9855 ( .IN1(n1036), .IN2(\fpu_mul_frac_dp/n838 ), .QN(n9231) );
  AO221X1 U9856 ( .IN1(n1367), .IN2(n9352), .IN3(n1361), .IN4(n9437), .IN5(
        n9538), .Q(n9365) );
  AO22X1 U9857 ( .IN1(n1378), .IN2(n9353), .IN3(n1369), .IN4(n9350), .Q(n9538)
         );
  AO221X1 U9858 ( .IN1(m4stg_frac[64]), .IN2(n1414), .IN3(m4stg_frac[63]), 
        .IN4(n1424), .IN5(n9539), .Q(n9350) );
  AO22X1 U9859 ( .IN1(m4stg_frac[62]), .IN2(n1435), .IN3(m4stg_frac[61]), 
        .IN4(n1441), .Q(n9539) );
  AO221X1 U9860 ( .IN1(m4stg_frac[60]), .IN2(n1414), .IN3(m4stg_frac[59]), 
        .IN4(n1424), .IN5(n9540), .Q(n9353) );
  AO22X1 U9861 ( .IN1(m4stg_frac[58]), .IN2(n1435), .IN3(m4stg_frac[57]), 
        .IN4(n1441), .Q(n9540) );
  AO221X1 U9862 ( .IN1(m4stg_frac[72]), .IN2(n1414), .IN3(m4stg_frac[71]), 
        .IN4(n1424), .IN5(n9541), .Q(n9437) );
  AO22X1 U9863 ( .IN1(m4stg_frac[70]), .IN2(n1435), .IN3(m4stg_frac[69]), 
        .IN4(n1441), .Q(n9541) );
  AO221X1 U9864 ( .IN1(m4stg_frac[68]), .IN2(n1414), .IN3(m4stg_frac[67]), 
        .IN4(n1424), .IN5(n9542), .Q(n9352) );
  AO22X1 U9865 ( .IN1(m4stg_frac[66]), .IN2(n1435), .IN3(m4stg_frac[65]), 
        .IN4(n1441), .Q(n9542) );
  NAND2X0 U9866 ( .IN1(n1357), .IN2(n9543), .QN(n9229) );
  NAND3X0 U9867 ( .IN1(n9227), .IN2(n9228), .IN3(n9225), .QN(n9543) );
  NOR2X0 U9868 ( .IN1(n603), .IN2(m4stg_inc_exp_55), .QN(n9225) );
  NOR2X0 U9869 ( .IN1(n9459), .IN2(n1033), .QN(n9228) );
  INVX0 U9870 ( .INP(n9187), .ZN(n9227) );
  NAND2X0 U9871 ( .IN1(\fpu_mul_frac_dp/n767 ), .IN2(\fpu_mul_frac_dp/n838 ), 
        .QN(n9187) );
  NAND2X0 U9872 ( .IN1(n9544), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N9 ) );
  OAI21X1 U9873 ( .IN1(n9546), .IN2(se_mul), .IN3(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N8 ) );
  NAND2X0 U9874 ( .IN1(n9547), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N7 ) );
  NAND2X0 U9875 ( .IN1(n9548), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N6 ) );
  NAND2X0 U9876 ( .IN1(n9549), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N57 ) );
  NAND2X0 U9877 ( .IN1(n9550), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N56 ) );
  NAND2X0 U9878 ( .IN1(n9551), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N55 ) );
  NAND2X0 U9879 ( .IN1(n9552), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N54 ) );
  NAND2X0 U9880 ( .IN1(n9553), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N53 ) );
  NAND2X0 U9881 ( .IN1(n9554), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N52 ) );
  NAND2X0 U9882 ( .IN1(n9555), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N51 ) );
  NAND2X0 U9883 ( .IN1(n9556), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N50 ) );
  NAND2X0 U9884 ( .IN1(n9557), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N5 ) );
  NAND2X0 U9885 ( .IN1(n9558), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N49 ) );
  NAND2X0 U9886 ( .IN1(n9559), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N48 ) );
  NAND2X0 U9887 ( .IN1(n9560), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N47 ) );
  NAND2X0 U9888 ( .IN1(n9561), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N46 ) );
  NAND2X0 U9889 ( .IN1(n9562), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N45 ) );
  NAND2X0 U9890 ( .IN1(n9563), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N44 ) );
  OAI21X1 U9891 ( .IN1(n9564), .IN2(se_mul), .IN3(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N43 ) );
  NAND2X0 U9892 ( .IN1(n9565), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N42 ) );
  OAI21X1 U9893 ( .IN1(n9566), .IN2(se_mul), .IN3(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N41 ) );
  NAND2X0 U9894 ( .IN1(n9567), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N40 ) );
  OR2X1 U9895 ( .IN1(n9568), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N4 ) );
  OAI21X1 U9896 ( .IN1(n9570), .IN2(se_mul), .IN3(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N39 ) );
  NAND2X0 U9897 ( .IN1(n9571), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N38 ) );
  OAI21X1 U9898 ( .IN1(n9572), .IN2(se_mul), .IN3(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N37 ) );
  NAND2X0 U9899 ( .IN1(n9573), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N36 ) );
  NAND2X0 U9900 ( .IN1(n9574), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N35 ) );
  NAND2X0 U9901 ( .IN1(n9575), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N34 ) );
  NAND2X0 U9902 ( .IN1(n9576), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N33 ) );
  NAND2X0 U9903 ( .IN1(n9577), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N32 ) );
  NAND2X0 U9904 ( .IN1(n9578), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N31 ) );
  NAND2X0 U9905 ( .IN1(n9579), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N30 ) );
  NAND2X0 U9906 ( .IN1(n9580), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N29 ) );
  NAND2X0 U9907 ( .IN1(n9581), .IN2(n9545), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N28 ) );
  INVX0 U9908 ( .INP(n9569), .ZN(n9545) );
  OR2X1 U9909 ( .IN1(n9582), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N27 ) );
  OR2X1 U9910 ( .IN1(n9583), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N26 ) );
  OR2X1 U9911 ( .IN1(n9584), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N25 ) );
  OR2X1 U9912 ( .IN1(n9585), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N24 ) );
  OR2X1 U9913 ( .IN1(n9586), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N23 ) );
  OR2X1 U9914 ( .IN1(n9587), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N22 ) );
  OR2X1 U9915 ( .IN1(n9588), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N21 ) );
  OR2X1 U9916 ( .IN1(n9589), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N20 ) );
  OR2X1 U9917 ( .IN1(n9590), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N19 ) );
  OR2X1 U9918 ( .IN1(n9591), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N18 ) );
  OR2X1 U9919 ( .IN1(n9592), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N17 ) );
  OR2X1 U9920 ( .IN1(n9593), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N16 ) );
  OR2X1 U9921 ( .IN1(n9594), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N15 ) );
  OR2X1 U9922 ( .IN1(n9595), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N14 ) );
  OR2X1 U9923 ( .IN1(n9596), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N13 ) );
  OR2X1 U9924 ( .IN1(n9597), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N12 ) );
  OR2X1 U9925 ( .IN1(n9598), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N11 ) );
  OR2X1 U9926 ( .IN1(n9599), .IN2(n9569), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre2/N10 ) );
  OA21X1 U9927 ( .IN1(n9600), .IN2(m4stg_shl_55), .IN3(n1357), .Q(n9569) );
  OA22X1 U9928 ( .IN1(n9601), .IN2(n9599), .IN3(n8872), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N9 ) );
  AO221X1 U9929 ( .IN1(n9602), .IN2(n9603), .IN3(n9604), .IN4(n9605), .IN5(
        n9606), .Q(n9599) );
  AO22X1 U9930 ( .IN1(n9607), .IN2(n9608), .IN3(n9609), .IN4(n9610), .Q(n9606)
         );
  AOI22X1 U9931 ( .IN1(n9544), .IN2(n9611), .IN3(n8866), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N8 ) );
  AO221X1 U9932 ( .IN1(n9612), .IN2(n9613), .IN3(n9614), .IN4(n9615), .IN5(
        n9616), .Q(n9544) );
  AO221X1 U9933 ( .IN1(n9617), .IN2(n9618), .IN3(n9619), .IN4(n9620), .IN5(
        se_mul), .Q(n9616) );
  MUX21X1 U9934 ( .IN1(n9621), .IN2(n9622), .S(\fpu_mul_frac_dp/n833 ), .Q(
        n9617) );
  OA22X1 U9935 ( .IN1(n8861), .IN2(n2929), .IN3(n9623), .IN4(n9601), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N7 ) );
  NOR2X0 U9936 ( .IN1(se_mul), .IN2(n9546), .QN(n9623) );
  AO221X1 U9937 ( .IN1(n9618), .IN2(n9624), .IN3(n9619), .IN4(n9625), .IN5(
        n9626), .Q(n9546) );
  AO22X1 U9938 ( .IN1(n9614), .IN2(n9627), .IN3(n9612), .IN4(n9628), .Q(n9626)
         );
  INVX0 U9939 ( .INP(n9029), .ZN(n8861) );
  AOI22X1 U9940 ( .IN1(n9547), .IN2(n9611), .IN3(n8867), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N6 ) );
  AO221X1 U9941 ( .IN1(n9612), .IN2(n9629), .IN3(n9619), .IN4(n9630), .IN5(
        n9631), .Q(n9547) );
  AO221X1 U9942 ( .IN1(n9618), .IN2(n9632), .IN3(n9614), .IN4(n9633), .IN5(
        se_mul), .Q(n9631) );
  OA221X1 U9943 ( .IN1(n9162), .IN2(n2929), .IN3(n9600), .IN4(n9634), .IN5(
        n1358), .Q(\fpu_mul_frac_dp/i_m5stg_frac_pre1/N57 ) );
  NAND2X0 U9944 ( .IN1(m4stg_shl_54), .IN2(m4stg_shl_55), .QN(n9634) );
  NAND4X0 U9945 ( .IN1(n9635), .IN2(n9636), .IN3(n9637), .IN4(n9638), .QN(
        m4stg_shl_54) );
  OA22X1 U9946 ( .IN1(n9639), .IN2(n9640), .IN3(n9641), .IN4(n9642), .Q(n9638)
         );
  OA22X1 U9947 ( .IN1(n9643), .IN2(n9520), .IN3(n1230), .IN4(n9307), .Q(n9641)
         );
  INVX0 U9948 ( .INP(n9644), .ZN(n9520) );
  AOI21X1 U9949 ( .IN1(\fpu_mul_frac_dp/n831 ), .IN2(m4stg_frac[102]), .IN3(
        \fpu_mul_frac_dp/n834 ), .QN(n9643) );
  NAND2X0 U9950 ( .IN1(n9644), .IN2(n884), .QN(n9640) );
  OA21X1 U9951 ( .IN1(n879), .IN2(m4stg_frac[103]), .IN3(n9307), .Q(n9644) );
  OA22X1 U9952 ( .IN1(n9645), .IN2(n9646), .IN3(n9647), .IN4(n9648), .Q(n9637)
         );
  INVX0 U9953 ( .INP(n9649), .ZN(n9645) );
  AOI22X1 U9954 ( .IN1(n9650), .IN2(n9651), .IN3(n9652), .IN4(n9614), .QN(
        n9636) );
  OA22X1 U9955 ( .IN1(n9653), .IN2(n9654), .IN3(n9604), .IN4(n9655), .Q(n9635)
         );
  INVX0 U9956 ( .INP(n9656), .ZN(n9162) );
  AOI22X1 U9957 ( .IN1(n9549), .IN2(n9611), .IN3(n9156), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N56 ) );
  NAND4X0 U9958 ( .IN1(n9657), .IN2(n9658), .IN3(n9659), .IN4(n9660), .QN(
        n9549) );
  OA221X1 U9959 ( .IN1(n9661), .IN2(n9639), .IN3(n9662), .IN4(n9642), .IN5(
        n1360), .Q(n9660) );
  AOI22X1 U9960 ( .IN1(n9663), .IN2(\fpu_mul_frac_dp/n834 ), .IN3(n1419), 
        .IN4(m4stg_frac[100]), .QN(n9662) );
  OA22X1 U9961 ( .IN1(n9664), .IN2(n9646), .IN3(n9665), .IN4(n9648), .Q(n9659)
         );
  INVX0 U9962 ( .INP(n9666), .ZN(n9664) );
  AOI22X1 U9963 ( .IN1(n9667), .IN2(n9651), .IN3(n9668), .IN4(n9614), .QN(
        n9658) );
  OA22X1 U9964 ( .IN1(n9669), .IN2(n9655), .IN3(n9670), .IN4(n9654), .Q(n9657)
         );
  AOI22X1 U9965 ( .IN1(n9550), .IN2(n9611), .IN3(n9151), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N55 ) );
  NAND4X0 U9966 ( .IN1(n9671), .IN2(n9672), .IN3(n9673), .IN4(n9674), .QN(
        n9550) );
  OA221X1 U9967 ( .IN1(n9675), .IN2(n9639), .IN3(n9676), .IN4(n9642), .IN5(
        n1359), .Q(n9674) );
  AOI222X1 U9968 ( .IN1(n1447), .IN2(m4stg_frac[102]), .IN3(n1411), .IN4(
        m4stg_frac[99]), .IN5(n1430), .IN6(m4stg_frac[100]), .QN(n9676) );
  NAND2X0 U9969 ( .IN1(n9677), .IN2(m4stg_frac[101]), .QN(n9639) );
  OA22X1 U9970 ( .IN1(n9678), .IN2(n9646), .IN3(n9679), .IN4(n9648), .Q(n9673)
         );
  INVX0 U9971 ( .INP(n9680), .ZN(n9678) );
  AOI22X1 U9972 ( .IN1(n9681), .IN2(n9651), .IN3(n9682), .IN4(n9614), .QN(
        n9672) );
  OA22X1 U9973 ( .IN1(n9683), .IN2(n9655), .IN3(n9684), .IN4(n9654), .Q(n9671)
         );
  AOI22X1 U9974 ( .IN1(n9551), .IN2(n9611), .IN3(n9145), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N54 ) );
  NAND4X0 U9975 ( .IN1(n9685), .IN2(n1358), .IN3(n9686), .IN4(n9687), .QN(
        n9551) );
  OA221X1 U9976 ( .IN1(n9688), .IN2(n9655), .IN3(n9689), .IN4(n9654), .IN5(
        n9690), .Q(n9687) );
  OA22X1 U9977 ( .IN1(n9691), .IN2(n9646), .IN3(n9692), .IN4(n9693), .Q(n9690)
         );
  OA22X1 U9978 ( .IN1(n9694), .IN2(n9648), .IN3(n9695), .IN4(n9696), .Q(n9686)
         );
  INVX0 U9979 ( .INP(n9697), .ZN(n9695) );
  NAND2X0 U9980 ( .IN1(n9677), .IN2(n9698), .QN(n9685) );
  AOI22X1 U9981 ( .IN1(n9552), .IN2(n9611), .IN3(n9140), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N53 ) );
  NAND4X0 U9982 ( .IN1(n9699), .IN2(n1359), .IN3(n9700), .IN4(n9701), .QN(
        n9552) );
  OA221X1 U9983 ( .IN1(n9702), .IN2(n9655), .IN3(n9703), .IN4(n9654), .IN5(
        n9704), .Q(n9701) );
  AOI22X1 U9984 ( .IN1(n9705), .IN2(n9651), .IN3(n9706), .IN4(n9614), .QN(
        n9704) );
  OA22X1 U9985 ( .IN1(n9647), .IN2(n9646), .IN3(n9707), .IN4(n9648), .Q(n9700)
         );
  INVX0 U9986 ( .INP(n9708), .ZN(n9647) );
  NAND2X0 U9987 ( .IN1(n9677), .IN2(n9649), .QN(n9699) );
  AO221X1 U9988 ( .IN1(m4stg_frac[97]), .IN2(n1414), .IN3(m4stg_frac[98]), 
        .IN4(n1424), .IN5(n9709), .Q(n9649) );
  AO22X1 U9989 ( .IN1(m4stg_frac[99]), .IN2(n1435), .IN3(m4stg_frac[100]), 
        .IN4(n1442), .Q(n9709) );
  AOI22X1 U9990 ( .IN1(n9553), .IN2(n9611), .IN3(n9134), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N52 ) );
  NAND4X0 U9991 ( .IN1(n9710), .IN2(n1360), .IN3(n9711), .IN4(n9712), .QN(
        n9553) );
  OA221X1 U9992 ( .IN1(n9713), .IN2(n9654), .IN3(n9714), .IN4(n9655), .IN5(
        n9715), .Q(n9712) );
  AOI22X1 U9993 ( .IN1(n9716), .IN2(n9651), .IN3(n9717), .IN4(n9614), .QN(
        n9715) );
  OA22X1 U9994 ( .IN1(n9665), .IN2(n9646), .IN3(n9718), .IN4(n9648), .Q(n9711)
         );
  INVX0 U9995 ( .INP(n9719), .ZN(n9665) );
  NAND2X0 U9996 ( .IN1(n9677), .IN2(n9666), .QN(n9710) );
  AO221X1 U9997 ( .IN1(m4stg_frac[96]), .IN2(n1414), .IN3(m4stg_frac[97]), 
        .IN4(n1425), .IN5(n9720), .Q(n9666) );
  AO22X1 U9998 ( .IN1(m4stg_frac[98]), .IN2(n1435), .IN3(m4stg_frac[99]), 
        .IN4(n1442), .Q(n9720) );
  AOI22X1 U9999 ( .IN1(n9554), .IN2(n9611), .IN3(n9129), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N51 ) );
  NAND4X0 U10000 ( .IN1(n9721), .IN2(n1357), .IN3(n9722), .IN4(n9723), .QN(
        n9554) );
  OA221X1 U10001 ( .IN1(n9724), .IN2(n9654), .IN3(n9725), .IN4(n9655), .IN5(
        n9726), .Q(n9723) );
  AOI22X1 U10002 ( .IN1(n9727), .IN2(n9651), .IN3(n9728), .IN4(n9614), .QN(
        n9726) );
  OA22X1 U10003 ( .IN1(n9679), .IN2(n9646), .IN3(n9729), .IN4(n9648), .Q(n9722) );
  INVX0 U10004 ( .INP(n9730), .ZN(n9679) );
  NAND2X0 U10005 ( .IN1(n9677), .IN2(n9680), .QN(n9721) );
  AO221X1 U10006 ( .IN1(m4stg_frac[95]), .IN2(n1414), .IN3(m4stg_frac[96]), 
        .IN4(n1425), .IN5(n9731), .Q(n9680) );
  AO22X1 U10007 ( .IN1(m4stg_frac[97]), .IN2(n1435), .IN3(m4stg_frac[98]), 
        .IN4(n1442), .Q(n9731) );
  INVX0 U10008 ( .INP(n9642), .ZN(n9677) );
  NAND2X0 U10009 ( .IN1(n1379), .IN2(n9619), .QN(n9642) );
  AOI22X1 U10010 ( .IN1(n9555), .IN2(n9611), .IN3(n9123), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N50 ) );
  NAND4X0 U10011 ( .IN1(n9732), .IN2(n1358), .IN3(n9733), .IN4(n9734), .QN(
        n9555) );
  OA221X1 U10012 ( .IN1(n9735), .IN2(n9654), .IN3(n9736), .IN4(n9655), .IN5(
        n9737), .Q(n9734) );
  OA22X1 U10013 ( .IN1(n9694), .IN2(n9646), .IN3(n9738), .IN4(n9693), .Q(n9737) );
  INVX0 U10014 ( .INP(n9739), .ZN(n9694) );
  OA22X1 U10015 ( .IN1(n9692), .IN2(n9648), .IN3(n9740), .IN4(n9696), .Q(n9733) );
  INVX0 U10016 ( .INP(n9741), .ZN(n9740) );
  NAND2X0 U10017 ( .IN1(n9742), .IN2(n9743), .QN(n9732) );
  AOI22X1 U10018 ( .IN1(n9548), .IN2(n9611), .IN3(n9744), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N5 ) );
  AO221X1 U10019 ( .IN1(n9612), .IN2(n9745), .IN3(n9619), .IN4(n9746), .IN5(
        n9747), .Q(n9548) );
  AO221X1 U10020 ( .IN1(n9618), .IN2(n9748), .IN3(n9614), .IN4(n9749), .IN5(
        se_mul), .Q(n9747) );
  AND2X1 U10021 ( .IN1(n9268), .IN2(n1035), .Q(n9618) );
  NOR2X0 U10022 ( .IN1(n1033), .IN2(\fpu_mul_frac_dp/n838 ), .QN(n9268) );
  AOI22X1 U10023 ( .IN1(n9556), .IN2(n9611), .IN3(n9118), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N49 ) );
  NAND4X0 U10024 ( .IN1(n9750), .IN2(n1359), .IN3(n9751), .IN4(n9752), .QN(
        n9556) );
  OA221X1 U10025 ( .IN1(n9753), .IN2(n9655), .IN3(n9754), .IN4(n9654), .IN5(
        n9755), .Q(n9752) );
  AOI22X1 U10026 ( .IN1(n9756), .IN2(n9651), .IN3(n9757), .IN4(n9614), .QN(
        n9755) );
  OA22X1 U10027 ( .IN1(n9707), .IN2(n9646), .IN3(n9758), .IN4(n9648), .Q(n9751) );
  INVX0 U10028 ( .INP(n9650), .ZN(n9707) );
  NAND2X0 U10029 ( .IN1(n9742), .IN2(n9708), .QN(n9750) );
  AO221X1 U10030 ( .IN1(m4stg_frac[93]), .IN2(n1414), .IN3(n1430), .IN4(
        m4stg_frac[94]), .IN5(n9759), .Q(n9708) );
  AO22X1 U10031 ( .IN1(m4stg_frac[95]), .IN2(n1435), .IN3(m4stg_frac[96]), 
        .IN4(n1442), .Q(n9759) );
  AOI22X1 U10032 ( .IN1(n9558), .IN2(n9611), .IN3(n9112), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N48 ) );
  NAND4X0 U10033 ( .IN1(n9760), .IN2(n1360), .IN3(n9761), .IN4(n9762), .QN(
        n9558) );
  OA221X1 U10034 ( .IN1(n9763), .IN2(n9654), .IN3(n9764), .IN4(n9655), .IN5(
        n9765), .Q(n9762) );
  AOI22X1 U10035 ( .IN1(n9766), .IN2(n9651), .IN3(n9767), .IN4(n9614), .QN(
        n9765) );
  OA22X1 U10036 ( .IN1(n9718), .IN2(n9646), .IN3(n9768), .IN4(n9648), .Q(n9761) );
  INVX0 U10037 ( .INP(n9667), .ZN(n9718) );
  NAND2X0 U10038 ( .IN1(n9742), .IN2(n9719), .QN(n9760) );
  AO221X1 U10039 ( .IN1(m4stg_frac[92]), .IN2(n1414), .IN3(m4stg_frac[93]), 
        .IN4(n1425), .IN5(n9769), .Q(n9719) );
  AO22X1 U10040 ( .IN1(m4stg_frac[94]), .IN2(n1435), .IN3(n1446), .IN4(
        m4stg_frac[95]), .Q(n9769) );
  AOI22X1 U10041 ( .IN1(n9559), .IN2(n9611), .IN3(n9107), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N47 ) );
  NAND4X0 U10042 ( .IN1(n9770), .IN2(n1357), .IN3(n9771), .IN4(n9772), .QN(
        n9559) );
  OA221X1 U10043 ( .IN1(n9773), .IN2(n9654), .IN3(n9774), .IN4(n9655), .IN5(
        n9775), .Q(n9772) );
  AOI22X1 U10044 ( .IN1(n9776), .IN2(n9651), .IN3(n9777), .IN4(n9614), .QN(
        n9775) );
  OA22X1 U10045 ( .IN1(n9729), .IN2(n9646), .IN3(n9778), .IN4(n9648), .Q(n9771) );
  INVX0 U10046 ( .INP(n9681), .ZN(n9729) );
  NAND2X0 U10047 ( .IN1(n9742), .IN2(n9730), .QN(n9770) );
  AO221X1 U10048 ( .IN1(m4stg_frac[91]), .IN2(n1415), .IN3(m4stg_frac[92]), 
        .IN4(n1425), .IN5(n9779), .Q(n9730) );
  AO22X1 U10049 ( .IN1(m4stg_frac[93]), .IN2(n1435), .IN3(n1446), .IN4(
        m4stg_frac[94]), .Q(n9779) );
  AOI22X1 U10050 ( .IN1(n9560), .IN2(n9611), .IN3(n9101), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N46 ) );
  NAND4X0 U10051 ( .IN1(n9780), .IN2(n1358), .IN3(n9781), .IN4(n9782), .QN(
        n9560) );
  OA221X1 U10052 ( .IN1(n9783), .IN2(n9654), .IN3(n9784), .IN4(n9655), .IN5(
        n9785), .Q(n9782) );
  OA22X1 U10053 ( .IN1(n9692), .IN2(n9646), .IN3(n9786), .IN4(n9693), .Q(n9785) );
  INVX0 U10054 ( .INP(n9787), .ZN(n9786) );
  INVX0 U10055 ( .INP(n9788), .ZN(n9692) );
  OA22X1 U10056 ( .IN1(n9738), .IN2(n9648), .IN3(n9789), .IN4(n9696), .Q(n9781) );
  INVX0 U10057 ( .INP(n9790), .ZN(n9789) );
  INVX0 U10058 ( .INP(n9791), .ZN(n9738) );
  NAND2X0 U10059 ( .IN1(n9742), .IN2(n9739), .QN(n9780) );
  AOI22X1 U10060 ( .IN1(n9561), .IN2(n9611), .IN3(n9096), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N45 ) );
  NAND4X0 U10061 ( .IN1(n9792), .IN2(n1359), .IN3(n9793), .IN4(n9794), .QN(
        n9561) );
  OA221X1 U10062 ( .IN1(n9795), .IN2(n9654), .IN3(n9796), .IN4(n9655), .IN5(
        n9797), .Q(n9794) );
  AOI22X1 U10063 ( .IN1(n9798), .IN2(n9651), .IN3(n9799), .IN4(n9614), .QN(
        n9797) );
  OA22X1 U10064 ( .IN1(n9800), .IN2(n9648), .IN3(n9758), .IN4(n9646), .Q(n9793) );
  INVX0 U10065 ( .INP(n9705), .ZN(n9758) );
  INVX0 U10066 ( .INP(n9756), .ZN(n9800) );
  NAND2X0 U10067 ( .IN1(n9742), .IN2(n9650), .QN(n9792) );
  AO221X1 U10068 ( .IN1(m4stg_frac[92]), .IN2(n1446), .IN3(m4stg_frac[91]), 
        .IN4(n1431), .IN5(n9801), .Q(n9650) );
  NAND2X0 U10069 ( .IN1(n9518), .IN2(n9489), .QN(n9801) );
  NAND2X0 U10070 ( .IN1(m4stg_frac[90]), .IN2(n9347), .QN(n9489) );
  NAND2X0 U10071 ( .IN1(m4stg_frac[89]), .IN2(n1420), .QN(n9518) );
  AOI22X1 U10072 ( .IN1(n9562), .IN2(n9611), .IN3(n9090), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N44 ) );
  NAND4X0 U10073 ( .IN1(n9802), .IN2(n1360), .IN3(n9803), .IN4(n9804), .QN(
        n9562) );
  OA221X1 U10074 ( .IN1(n9805), .IN2(n9654), .IN3(n9806), .IN4(n9655), .IN5(
        n9807), .Q(n9804) );
  AOI22X1 U10075 ( .IN1(n9808), .IN2(n9651), .IN3(n9809), .IN4(n9614), .QN(
        n9807) );
  OA22X1 U10076 ( .IN1(n9810), .IN2(n9648), .IN3(n9768), .IN4(n9646), .Q(n9803) );
  INVX0 U10077 ( .INP(n9716), .ZN(n9768) );
  INVX0 U10078 ( .INP(n9766), .ZN(n9810) );
  NAND2X0 U10079 ( .IN1(n9742), .IN2(n9667), .QN(n9802) );
  AO221X1 U10080 ( .IN1(m4stg_frac[88]), .IN2(n1415), .IN3(m4stg_frac[89]), 
        .IN4(n1425), .IN5(n9811), .Q(n9667) );
  AO22X1 U10081 ( .IN1(m4stg_frac[90]), .IN2(n1435), .IN3(m4stg_frac[91]), 
        .IN4(n1442), .Q(n9811) );
  AOI22X1 U10082 ( .IN1(n9563), .IN2(n9611), .IN3(n9084), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N43 ) );
  NAND4X0 U10083 ( .IN1(n9812), .IN2(n1357), .IN3(n9813), .IN4(n9814), .QN(
        n9563) );
  OA221X1 U10084 ( .IN1(n9815), .IN2(n9654), .IN3(n9816), .IN4(n9655), .IN5(
        n9817), .Q(n9814) );
  AOI22X1 U10085 ( .IN1(n9818), .IN2(n9651), .IN3(n9819), .IN4(n9614), .QN(
        n9817) );
  OA22X1 U10086 ( .IN1(n9820), .IN2(n9648), .IN3(n9778), .IN4(n9646), .Q(n9813) );
  INVX0 U10087 ( .INP(n9727), .ZN(n9778) );
  INVX0 U10088 ( .INP(n9776), .ZN(n9820) );
  NAND2X0 U10089 ( .IN1(n9742), .IN2(n9681), .QN(n9812) );
  AO221X1 U10090 ( .IN1(m4stg_frac[87]), .IN2(n1415), .IN3(m4stg_frac[88]), 
        .IN4(n1425), .IN5(n9821), .Q(n9681) );
  NAND2X0 U10091 ( .IN1(n9488), .IN2(n9524), .QN(n9821) );
  NAND2X0 U10092 ( .IN1(m4stg_frac[90]), .IN2(n1447), .QN(n9524) );
  NAND2X0 U10093 ( .IN1(m4stg_frac[89]), .IN2(n9349), .QN(n9488) );
  OA22X1 U10094 ( .IN1(n9078), .IN2(n2929), .IN3(n9822), .IN4(n9601), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N42 ) );
  NOR2X0 U10095 ( .IN1(se_mul), .IN2(n9564), .QN(n9822) );
  AO222X1 U10096 ( .IN1(n9614), .IN2(n9823), .IN3(n9824), .IN4(n1035), .IN5(
        n9619), .IN6(n9825), .Q(n9564) );
  INVX0 U10097 ( .INP(n9085), .ZN(n9078) );
  AOI22X1 U10098 ( .IN1(n9565), .IN2(n9611), .IN3(n9072), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N41 ) );
  AO221X1 U10099 ( .IN1(n9614), .IN2(n9826), .IN3(n9612), .IN4(n9827), .IN5(
        n9828), .Q(n9565) );
  AO221X1 U10100 ( .IN1(n9619), .IN2(n9652), .IN3(n9829), .IN4(n9830), .IN5(
        se_mul), .Q(n9828) );
  AO221X1 U10101 ( .IN1(n1380), .IN2(n9705), .IN3(n1369), .IN4(n9756), .IN5(
        n9831), .Q(n9652) );
  AO22X1 U10102 ( .IN1(n1361), .IN2(n9832), .IN3(n1366), .IN4(n9798), .Q(n9831) );
  AO221X1 U10103 ( .IN1(m4stg_frac[85]), .IN2(n1415), .IN3(m4stg_frac[86]), 
        .IN4(n1425), .IN5(n9833), .Q(n9705) );
  AO22X1 U10104 ( .IN1(m4stg_frac[87]), .IN2(n1435), .IN3(m4stg_frac[88]), 
        .IN4(n1442), .Q(n9833) );
  OA22X1 U10105 ( .IN1(n9066), .IN2(n2929), .IN3(n9834), .IN4(n9601), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N40 ) );
  NOR2X0 U10106 ( .IN1(se_mul), .IN2(n9566), .QN(n9834) );
  AO221X1 U10107 ( .IN1(n9619), .IN2(n9668), .IN3(n9612), .IN4(n9620), .IN5(
        n9835), .Q(n9566) );
  AO22X1 U10108 ( .IN1(n9829), .IN2(n9615), .IN3(n9614), .IN4(n9836), .Q(n9835) );
  AO221X1 U10109 ( .IN1(n1379), .IN2(n9716), .IN3(n1370), .IN4(n9766), .IN5(
        n9837), .Q(n9668) );
  AO22X1 U10110 ( .IN1(n1364), .IN2(n9838), .IN3(n1367), .IN4(n9808), .Q(n9837) );
  AO221X1 U10111 ( .IN1(m4stg_frac[84]), .IN2(n1415), .IN3(m4stg_frac[85]), 
        .IN4(n1425), .IN5(n9839), .Q(n9716) );
  AO22X1 U10112 ( .IN1(m4stg_frac[86]), .IN2(n1436), .IN3(m4stg_frac[87]), 
        .IN4(n1442), .Q(n9839) );
  INVX0 U10113 ( .INP(n9073), .ZN(n9066) );
  OA22X1 U10114 ( .IN1(n9840), .IN2(n9601), .IN3(n9841), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N4 ) );
  INVX0 U10115 ( .INP(n9557), .ZN(n9840) );
  AO221X1 U10116 ( .IN1(n9612), .IN2(n9842), .IN3(n9614), .IN4(n9843), .IN5(
        n9844), .Q(n9557) );
  AO221X1 U10117 ( .IN1(n9845), .IN2(n9829), .IN3(n9619), .IN4(n9846), .IN5(
        se_mul), .Q(n9844) );
  NOR2X0 U10118 ( .IN1(n9847), .IN2(n9304), .QN(n9845) );
  AOI22X1 U10119 ( .IN1(n9567), .IN2(n9611), .IN3(n9060), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N39 ) );
  AO221X1 U10120 ( .IN1(n9614), .IN2(n9848), .IN3(n9829), .IN4(n9627), .IN5(
        n9849), .Q(n9567) );
  AO221X1 U10121 ( .IN1(n9619), .IN2(n9682), .IN3(n9612), .IN4(n9625), .IN5(
        se_mul), .Q(n9849) );
  AO221X1 U10122 ( .IN1(n1378), .IN2(n9727), .IN3(n1372), .IN4(n9776), .IN5(
        n9850), .Q(n9682) );
  AO22X1 U10123 ( .IN1(n1362), .IN2(n9851), .IN3(n1368), .IN4(n9818), .Q(n9850) );
  AO221X1 U10124 ( .IN1(m4stg_frac[83]), .IN2(n1415), .IN3(m4stg_frac[84]), 
        .IN4(n1425), .IN5(n9852), .Q(n9727) );
  AO22X1 U10125 ( .IN1(m4stg_frac[85]), .IN2(n1436), .IN3(m4stg_frac[86]), 
        .IN4(n1442), .Q(n9852) );
  OA22X1 U10126 ( .IN1(n9054), .IN2(n2929), .IN3(n9853), .IN4(n9601), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N38 ) );
  NOR2X0 U10127 ( .IN1(se_mul), .IN2(n9570), .QN(n9853) );
  AO221X1 U10128 ( .IN1(n9619), .IN2(n9697), .IN3(n9829), .IN4(n9633), .IN5(
        n9854), .Q(n9570) );
  AO22X1 U10129 ( .IN1(n9612), .IN2(n9630), .IN3(n9614), .IN4(n9855), .Q(n9854) );
  AO221X1 U10130 ( .IN1(n1377), .IN2(n9791), .IN3(n1362), .IN4(n9856), .IN5(
        n9857), .Q(n9697) );
  AO22X1 U10131 ( .IN1(n1372), .IN2(n9787), .IN3(n1365), .IN4(n9858), .Q(n9857) );
  INVX0 U10132 ( .INP(n9061), .ZN(n9054) );
  AOI22X1 U10133 ( .IN1(n9571), .IN2(n9611), .IN3(n9048), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N37 ) );
  AO221X1 U10134 ( .IN1(n9614), .IN2(n9859), .IN3(n9612), .IN4(n9746), .IN5(
        n9860), .Q(n9571) );
  AO221X1 U10135 ( .IN1(n9619), .IN2(n9706), .IN3(n9829), .IN4(n9749), .IN5(
        se_mul), .Q(n9860) );
  AO221X1 U10136 ( .IN1(n1380), .IN2(n9756), .IN3(n1371), .IN4(n9798), .IN5(
        n9861), .Q(n9706) );
  AO22X1 U10137 ( .IN1(n1363), .IN2(n9862), .IN3(n1366), .IN4(n9832), .Q(n9861) );
  AO221X1 U10138 ( .IN1(m4stg_frac[81]), .IN2(n1415), .IN3(m4stg_frac[82]), 
        .IN4(n1425), .IN5(n9863), .Q(n9756) );
  AO22X1 U10139 ( .IN1(m4stg_frac[83]), .IN2(n1436), .IN3(m4stg_frac[84]), 
        .IN4(n1442), .Q(n9863) );
  OA22X1 U10140 ( .IN1(n9042), .IN2(n2929), .IN3(n9864), .IN4(n9601), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N36 ) );
  NOR2X0 U10141 ( .IN1(se_mul), .IN2(n9572), .QN(n9864) );
  AO221X1 U10142 ( .IN1(n9619), .IN2(n9717), .IN3(n9612), .IN4(n9846), .IN5(
        n9865), .Q(n9572) );
  AO22X1 U10143 ( .IN1(n9829), .IN2(n9843), .IN3(n9614), .IN4(n9866), .Q(n9865) );
  INVX0 U10144 ( .INP(n9655), .ZN(n9829) );
  INVX0 U10145 ( .INP(n9654), .ZN(n9612) );
  AO221X1 U10146 ( .IN1(n1379), .IN2(n9766), .IN3(n1369), .IN4(n9808), .IN5(
        n9867), .Q(n9717) );
  AO22X1 U10147 ( .IN1(n1361), .IN2(n9868), .IN3(n1367), .IN4(n9838), .Q(n9867) );
  AO221X1 U10148 ( .IN1(m4stg_frac[80]), .IN2(n1415), .IN3(m4stg_frac[81]), 
        .IN4(n1425), .IN5(n9869), .Q(n9766) );
  AO22X1 U10149 ( .IN1(m4stg_frac[82]), .IN2(n1436), .IN3(m4stg_frac[83]), 
        .IN4(n1442), .Q(n9869) );
  INVX0 U10150 ( .INP(n9049), .ZN(n9042) );
  AOI22X1 U10151 ( .IN1(n9573), .IN2(n9611), .IN3(n9032), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N35 ) );
  AO221X1 U10152 ( .IN1(n9619), .IN2(n9728), .IN3(n9614), .IN4(n9870), .IN5(
        n9871), .Q(n9573) );
  OA221X1 U10153 ( .IN1(n9872), .IN2(n9873), .IN3(n9874), .IN4(n9875), .IN5(
        n9876), .Q(n9871) );
  AO221X1 U10154 ( .IN1(n1378), .IN2(n9776), .IN3(n1370), .IN4(n9818), .IN5(
        n9877), .Q(n9728) );
  AO22X1 U10155 ( .IN1(n1364), .IN2(n9878), .IN3(n1368), .IN4(n9851), .Q(n9877) );
  AO221X1 U10156 ( .IN1(m4stg_frac[79]), .IN2(n1415), .IN3(m4stg_frac[80]), 
        .IN4(n1425), .IN5(n9879), .Q(n9776) );
  AO22X1 U10157 ( .IN1(m4stg_frac[81]), .IN2(n1436), .IN3(m4stg_frac[82]), 
        .IN4(n1442), .Q(n9879) );
  AOI22X1 U10158 ( .IN1(n9574), .IN2(n9611), .IN3(n9019), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N34 ) );
  AO221X1 U10159 ( .IN1(n9619), .IN2(n9741), .IN3(n9614), .IN4(n9880), .IN5(
        n9881), .Q(n9574) );
  OA221X1 U10160 ( .IN1(n9882), .IN2(n9873), .IN3(n9883), .IN4(n9875), .IN5(
        n9876), .Q(n9881) );
  AO221X1 U10161 ( .IN1(n1371), .IN2(n9858), .IN3(n1380), .IN4(n9787), .IN5(
        n9884), .Q(n9741) );
  AO22X1 U10162 ( .IN1(n1362), .IN2(n9885), .IN3(n1365), .IN4(n9856), .Q(n9884) );
  AOI22X1 U10163 ( .IN1(n9575), .IN2(n9611), .IN3(n9013), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N33 ) );
  AO221X1 U10164 ( .IN1(n9619), .IN2(n9757), .IN3(n9614), .IN4(n9886), .IN5(
        n9887), .Q(n9575) );
  OA221X1 U10165 ( .IN1(n9888), .IN2(n9873), .IN3(n9889), .IN4(n9875), .IN5(
        n9876), .Q(n9887) );
  AO221X1 U10166 ( .IN1(n1377), .IN2(n9798), .IN3(n1372), .IN4(n9832), .IN5(
        n9890), .Q(n9757) );
  AO22X1 U10167 ( .IN1(n1363), .IN2(n9891), .IN3(n1366), .IN4(n9862), .Q(n9890) );
  AO221X1 U10168 ( .IN1(m4stg_frac[77]), .IN2(n1415), .IN3(m4stg_frac[78]), 
        .IN4(n1426), .IN5(n9892), .Q(n9798) );
  AO22X1 U10169 ( .IN1(m4stg_frac[79]), .IN2(n1436), .IN3(m4stg_frac[80]), 
        .IN4(n1442), .Q(n9892) );
  AOI22X1 U10170 ( .IN1(n9576), .IN2(n9611), .IN3(n9008), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N32 ) );
  AO221X1 U10171 ( .IN1(n9619), .IN2(n9767), .IN3(n9614), .IN4(n9893), .IN5(
        n9894), .Q(n9576) );
  OA221X1 U10172 ( .IN1(n9895), .IN2(n9873), .IN3(n9896), .IN4(n9875), .IN5(
        n9876), .Q(n9894) );
  AO221X1 U10173 ( .IN1(n1380), .IN2(n9808), .IN3(n1371), .IN4(n9838), .IN5(
        n9897), .Q(n9767) );
  AO22X1 U10174 ( .IN1(n1361), .IN2(n9898), .IN3(n1367), .IN4(n9868), .Q(n9897) );
  AO221X1 U10175 ( .IN1(m4stg_frac[76]), .IN2(n1415), .IN3(m4stg_frac[77]), 
        .IN4(n1426), .IN5(n9899), .Q(n9808) );
  AO22X1 U10176 ( .IN1(m4stg_frac[78]), .IN2(n1436), .IN3(m4stg_frac[79]), 
        .IN4(n1442), .Q(n9899) );
  AOI22X1 U10177 ( .IN1(n9577), .IN2(n9611), .IN3(n9002), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N31 ) );
  AO221X1 U10178 ( .IN1(n9619), .IN2(n9777), .IN3(n9614), .IN4(n9900), .IN5(
        n9901), .Q(n9577) );
  OA221X1 U10179 ( .IN1(n9902), .IN2(n9873), .IN3(n9903), .IN4(n9875), .IN5(
        n9876), .Q(n9901) );
  AO221X1 U10180 ( .IN1(n1379), .IN2(n9818), .IN3(n1369), .IN4(n9851), .IN5(
        n9904), .Q(n9777) );
  AO22X1 U10181 ( .IN1(n1364), .IN2(n9905), .IN3(n1368), .IN4(n9878), .Q(n9904) );
  AO221X1 U10182 ( .IN1(m4stg_frac[75]), .IN2(n1415), .IN3(m4stg_frac[76]), 
        .IN4(n1426), .IN5(n9906), .Q(n9818) );
  AO22X1 U10183 ( .IN1(m4stg_frac[77]), .IN2(n1436), .IN3(m4stg_frac[78]), 
        .IN4(n1442), .Q(n9906) );
  AOI22X1 U10184 ( .IN1(n9578), .IN2(n9611), .IN3(n8997), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N30 ) );
  AO221X1 U10185 ( .IN1(n9619), .IN2(n9790), .IN3(n9614), .IN4(n9907), .IN5(
        n9908), .Q(n9578) );
  OA221X1 U10186 ( .IN1(n9909), .IN2(n9873), .IN3(n9910), .IN4(n9875), .IN5(
        n9876), .Q(n9908) );
  AO221X1 U10187 ( .IN1(n1378), .IN2(n9858), .IN3(n1364), .IN4(n9911), .IN5(
        n9912), .Q(n9790) );
  AO22X1 U10188 ( .IN1(n1366), .IN2(n9885), .IN3(n1370), .IN4(n9856), .Q(n9912) );
  OA22X1 U10189 ( .IN1(n9568), .IN2(n9601), .IN3(n9913), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N3 ) );
  OA221X1 U10190 ( .IN1(n9914), .IN2(n9304), .IN3(n9915), .IN4(n1035), .IN5(
        n9916), .Q(n9568) );
  OA21X1 U10191 ( .IN1(n9917), .IN2(n908), .IN3(n1358), .Q(n9916) );
  OA21X1 U10192 ( .IN1(n9918), .IN2(n1035), .IN3(n9919), .Q(n9917) );
  NOR4X0 U10193 ( .IN1(n9920), .IN2(n9921), .IN3(n9922), .IN4(n9923), .QN(
        n9918) );
  NAND4X0 U10194 ( .IN1(n9924), .IN2(n9925), .IN3(n9926), .IN4(n9927), .QN(
        n9923) );
  NAND4X0 U10195 ( .IN1(n9725), .IN2(n9736), .IN3(n9753), .IN4(n9928), .QN(
        n9922) );
  NAND4X0 U10196 ( .IN1(n9764), .IN2(n9774), .IN3(n9784), .IN4(n9796), .QN(
        n9921) );
  NAND4X0 U10197 ( .IN1(n9806), .IN2(n9816), .IN3(n9608), .IN4(n9929), .QN(
        n9920) );
  NOR4X0 U10198 ( .IN1(n9930), .IN2(n9931), .IN3(n9932), .IN4(n9933), .QN(
        n9915) );
  NAND4X0 U10199 ( .IN1(n9934), .IN2(n9603), .IN3(n9935), .IN4(n9936), .QN(
        n9933) );
  NAND4X0 U10200 ( .IN1(n9937), .IN2(n9938), .IN3(n9939), .IN4(n9940), .QN(
        n9932) );
  NAND4X0 U10201 ( .IN1(n9941), .IN2(n9942), .IN3(n9943), .IN4(n9944), .QN(
        n9931) );
  NAND4X0 U10202 ( .IN1(n9945), .IN2(n9919), .IN3(n9946), .IN4(n9947), .QN(
        n9930) );
  NOR2X0 U10203 ( .IN1(n9882), .IN2(n9888), .QN(n9947) );
  NOR4X0 U10204 ( .IN1(n9948), .IN2(n9949), .IN3(n9950), .IN4(n9951), .QN(
        n9919) );
  NAND4X0 U10205 ( .IN1(n9952), .IN2(n9953), .IN3(n9954), .IN4(n9610), .QN(
        n9951) );
  AOI222X1 U10206 ( .IN1(n1377), .IN2(n9955), .IN3(n9956), .IN4(m4stg_frac[0]), 
        .IN5(n1372), .IN6(n9957), .QN(n9610) );
  AND2X1 U10207 ( .IN1(n1447), .IN2(n1365), .Q(n9956) );
  INVX0 U10208 ( .INP(n9624), .ZN(n9954) );
  NAND4X0 U10209 ( .IN1(n9958), .IN2(n9959), .IN3(n9847), .IN4(n9960), .QN(
        n9950) );
  NAND2X0 U10210 ( .IN1(\fpu_mul_frac_dp/n833 ), .IN2(n9622), .QN(n9960) );
  INVX0 U10211 ( .INP(n9621), .ZN(n9847) );
  NAND4X0 U10212 ( .IN1(n9961), .IN2(n9962), .IN3(n9963), .IN4(n9964), .QN(
        n9949) );
  NAND4X0 U10213 ( .IN1(n9965), .IN2(n9966), .IN3(n9967), .IN4(n9968), .QN(
        n9948) );
  NOR2X0 U10214 ( .IN1(n9969), .IN2(n9970), .QN(n9914) );
  OA21X1 U10215 ( .IN1(m4stg_frac[1]), .IN2(m4stg_frac[0]), .IN3(
        \fpu_mul_frac_dp/n834 ), .Q(n9969) );
  AOI22X1 U10216 ( .IN1(n9579), .IN2(n9611), .IN3(n8991), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N29 ) );
  AO221X1 U10217 ( .IN1(n9619), .IN2(n9799), .IN3(n9614), .IN4(n9971), .IN5(
        n9972), .Q(n9579) );
  OA221X1 U10218 ( .IN1(n9973), .IN2(n9873), .IN3(n9974), .IN4(n9875), .IN5(
        n9876), .Q(n9972) );
  AO221X1 U10219 ( .IN1(n1377), .IN2(n9832), .IN3(n1370), .IN4(n9862), .IN5(
        n9975), .Q(n9799) );
  AO22X1 U10220 ( .IN1(n1362), .IN2(n9976), .IN3(n1365), .IN4(n9891), .Q(n9975) );
  AO221X1 U10221 ( .IN1(m4stg_frac[73]), .IN2(n1415), .IN3(m4stg_frac[74]), 
        .IN4(n1426), .IN5(n9977), .Q(n9832) );
  AO22X1 U10222 ( .IN1(m4stg_frac[75]), .IN2(n1436), .IN3(m4stg_frac[76]), 
        .IN4(n1442), .Q(n9977) );
  AOI22X1 U10223 ( .IN1(n9580), .IN2(n9611), .IN3(n8986), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N28 ) );
  AO221X1 U10224 ( .IN1(n9619), .IN2(n9809), .IN3(n9614), .IN4(n9978), .IN5(
        n9979), .Q(n9580) );
  OA221X1 U10225 ( .IN1(n9980), .IN2(n9873), .IN3(n9981), .IN4(n9875), .IN5(
        n9876), .Q(n9979) );
  AO221X1 U10226 ( .IN1(n1380), .IN2(n9838), .IN3(n1372), .IN4(n9868), .IN5(
        n9982), .Q(n9809) );
  AO22X1 U10227 ( .IN1(n1363), .IN2(n9983), .IN3(n1366), .IN4(n9898), .Q(n9982) );
  AO221X1 U10228 ( .IN1(m4stg_frac[72]), .IN2(n1416), .IN3(m4stg_frac[73]), 
        .IN4(n1426), .IN5(n9984), .Q(n9838) );
  AO22X1 U10229 ( .IN1(m4stg_frac[74]), .IN2(n1436), .IN3(m4stg_frac[75]), 
        .IN4(n1442), .Q(n9984) );
  AOI22X1 U10230 ( .IN1(n9581), .IN2(n9611), .IN3(n8980), .IN4(n603), .QN(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N27 ) );
  INVX0 U10231 ( .INP(n9601), .ZN(n9611) );
  AO221X1 U10232 ( .IN1(n9619), .IN2(n9819), .IN3(n9614), .IN4(n9985), .IN5(
        n9986), .Q(n9581) );
  OA221X1 U10233 ( .IN1(n9987), .IN2(n9873), .IN3(n9988), .IN4(n9875), .IN5(
        n9876), .Q(n9986) );
  NAND2X0 U10234 ( .IN1(\fpu_mul_frac_dp/n838 ), .IN2(n1360), .QN(n9875) );
  NAND2X0 U10235 ( .IN1(n908), .IN2(n1357), .QN(n9873) );
  AO221X1 U10236 ( .IN1(n1379), .IN2(n9851), .IN3(n1371), .IN4(n9878), .IN5(
        n9989), .Q(n9819) );
  AO22X1 U10237 ( .IN1(n1361), .IN2(n9990), .IN3(n1367), .IN4(n9905), .Q(n9989) );
  AO221X1 U10238 ( .IN1(m4stg_frac[71]), .IN2(n1416), .IN3(m4stg_frac[72]), 
        .IN4(n1426), .IN5(n9991), .Q(n9851) );
  AO22X1 U10239 ( .IN1(m4stg_frac[73]), .IN2(n1436), .IN3(m4stg_frac[74]), 
        .IN4(n1443), .Q(n9991) );
  OA22X1 U10240 ( .IN1(n9601), .IN2(n9582), .IN3(n8974), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N26 ) );
  INVX0 U10241 ( .INP(n9020), .ZN(n8974) );
  AO221X1 U10242 ( .IN1(n9607), .IN2(n9992), .IN3(n9993), .IN4(n9605), .IN5(
        n9994), .Q(n9582) );
  AO22X1 U10243 ( .IN1(n9602), .IN2(n9929), .IN3(n9609), .IN4(n9934), .Q(n9994) );
  INVX0 U10244 ( .INP(n9995), .ZN(n9929) );
  OA22X1 U10245 ( .IN1(n9601), .IN2(n9583), .IN3(n8968), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N25 ) );
  AO221X1 U10246 ( .IN1(n9653), .IN2(n9605), .IN3(n9604), .IN4(n9607), .IN5(
        n9996), .Q(n9583) );
  AO22X1 U10247 ( .IN1(n9609), .IN2(n9603), .IN3(n9602), .IN4(n9608), .Q(n9996) );
  INVX0 U10248 ( .INP(n9830), .ZN(n9608) );
  AO222X1 U10249 ( .IN1(n1378), .IN2(n9997), .IN3(n9998), .IN4(n1033), .IN5(
        n1372), .IN6(n9999), .Q(n9830) );
  AOI221X1 U10250 ( .IN1(n1378), .IN2(n10000), .IN3(n1371), .IN4(n10001), 
        .IN5(n10002), .QN(n9603) );
  AO22X1 U10251 ( .IN1(n1367), .IN2(n10003), .IN3(n1364), .IN4(n10004), .Q(
        n10002) );
  INVX0 U10252 ( .INP(n9827), .ZN(n9604) );
  AO221X1 U10253 ( .IN1(n1370), .IN2(n10005), .IN3(n1379), .IN4(n10006), .IN5(
        n10007), .Q(n9827) );
  AO22X1 U10254 ( .IN1(n1368), .IN2(n10008), .IN3(n1363), .IN4(n10009), .Q(
        n10007) );
  INVX0 U10255 ( .INP(n9826), .ZN(n9653) );
  AO221X1 U10256 ( .IN1(n1378), .IN2(n9862), .IN3(n1369), .IN4(n9891), .IN5(
        n10010), .Q(n9826) );
  AO22X1 U10257 ( .IN1(n1364), .IN2(n10011), .IN3(n1368), .IN4(n9976), .Q(
        n10010) );
  AO221X1 U10258 ( .IN1(m4stg_frac[69]), .IN2(n1416), .IN3(m4stg_frac[70]), 
        .IN4(n1426), .IN5(n10012), .Q(n9862) );
  AO22X1 U10259 ( .IN1(m4stg_frac[71]), .IN2(n1436), .IN3(m4stg_frac[72]), 
        .IN4(n1443), .Q(n10012) );
  OA22X1 U10260 ( .IN1(n9601), .IN2(n9584), .IN3(n8962), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N24 ) );
  AO221X1 U10261 ( .IN1(n9609), .IN2(n9935), .IN3(n9602), .IN4(n9924), .IN5(
        n10013), .Q(n9584) );
  AO22X1 U10262 ( .IN1(n9670), .IN2(n9605), .IN3(n9669), .IN4(n9607), .Q(
        n10013) );
  INVX0 U10263 ( .INP(n9620), .ZN(n9669) );
  AO221X1 U10264 ( .IN1(n1369), .IN2(n10014), .IN3(n1377), .IN4(n10015), .IN5(
        n10016), .Q(n9620) );
  AO22X1 U10265 ( .IN1(n1365), .IN2(n10017), .IN3(n1361), .IN4(n10018), .Q(
        n10016) );
  INVX0 U10266 ( .INP(n9836), .ZN(n9670) );
  AO221X1 U10267 ( .IN1(n1377), .IN2(n9868), .IN3(n1370), .IN4(n9898), .IN5(
        n10019), .Q(n9836) );
  AO22X1 U10268 ( .IN1(n1362), .IN2(n10020), .IN3(n1365), .IN4(n9983), .Q(
        n10019) );
  AO221X1 U10269 ( .IN1(m4stg_frac[68]), .IN2(n1416), .IN3(m4stg_frac[69]), 
        .IN4(n1426), .IN5(n10021), .Q(n9868) );
  AO22X1 U10270 ( .IN1(m4stg_frac[70]), .IN2(n1436), .IN3(m4stg_frac[71]), 
        .IN4(n1443), .Q(n10021) );
  INVX0 U10271 ( .INP(n9615), .ZN(n9924) );
  AO222X1 U10272 ( .IN1(n1370), .IN2(n10022), .IN3(n10023), .IN4(n1033), .IN5(
        n1378), .IN6(n10024), .Q(n9615) );
  INVX0 U10273 ( .INP(n9613), .ZN(n9935) );
  AO222X1 U10274 ( .IN1(n1371), .IN2(n10025), .IN3(n10026), .IN4(n1033), .IN5(
        n1380), .IN6(n10027), .Q(n9613) );
  OA22X1 U10275 ( .IN1(n9601), .IN2(n9585), .IN3(n8956), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N23 ) );
  AO221X1 U10276 ( .IN1(n9609), .IN2(n9936), .IN3(n9602), .IN4(n9925), .IN5(
        n10028), .Q(n9585) );
  AO22X1 U10277 ( .IN1(n9684), .IN2(n9605), .IN3(n9683), .IN4(n9607), .Q(
        n10028) );
  INVX0 U10278 ( .INP(n9625), .ZN(n9683) );
  AO221X1 U10279 ( .IN1(n1363), .IN2(n10029), .IN3(n1378), .IN4(n10030), .IN5(
        n10031), .Q(n9625) );
  AO22X1 U10280 ( .IN1(n1366), .IN2(n10032), .IN3(n1372), .IN4(n10033), .Q(
        n10031) );
  INVX0 U10281 ( .INP(n9848), .ZN(n9684) );
  AO221X1 U10282 ( .IN1(n1380), .IN2(n9878), .IN3(n1372), .IN4(n9905), .IN5(
        n10034), .Q(n9848) );
  AO22X1 U10283 ( .IN1(n1363), .IN2(n10035), .IN3(n1366), .IN4(n9990), .Q(
        n10034) );
  AO221X1 U10284 ( .IN1(m4stg_frac[67]), .IN2(n1416), .IN3(m4stg_frac[68]), 
        .IN4(n1426), .IN5(n10036), .Q(n9878) );
  AO22X1 U10285 ( .IN1(m4stg_frac[69]), .IN2(n1436), .IN3(m4stg_frac[70]), 
        .IN4(n1443), .Q(n10036) );
  INVX0 U10286 ( .INP(n9627), .ZN(n9925) );
  AO222X1 U10287 ( .IN1(n1372), .IN2(n10037), .IN3(n10038), .IN4(n1033), .IN5(
        n1377), .IN6(n10039), .Q(n9627) );
  INVX0 U10288 ( .INP(n9628), .ZN(n9936) );
  AO221X1 U10289 ( .IN1(n1362), .IN2(n10040), .IN3(n1380), .IN4(n10041), .IN5(
        n10042), .Q(n9628) );
  AO22X1 U10290 ( .IN1(n1367), .IN2(n10043), .IN3(n1371), .IN4(n10044), .Q(
        n10042) );
  OA22X1 U10291 ( .IN1(n9601), .IN2(n9586), .IN3(n8950), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N22 ) );
  AO221X1 U10292 ( .IN1(n9602), .IN2(n9926), .IN3(n9609), .IN4(n9937), .IN5(
        n10045), .Q(n9586) );
  AO22X1 U10293 ( .IN1(n9688), .IN2(n9607), .IN3(n9689), .IN4(n9605), .Q(
        n10045) );
  INVX0 U10294 ( .INP(n9855), .ZN(n9689) );
  AO221X1 U10295 ( .IN1(n1379), .IN2(n9885), .IN3(n1363), .IN4(n10046), .IN5(
        n10047), .Q(n9855) );
  AO22X1 U10296 ( .IN1(n1369), .IN2(n9911), .IN3(n1367), .IN4(n10048), .Q(
        n10047) );
  INVX0 U10297 ( .INP(n9630), .ZN(n9688) );
  AO221X1 U10298 ( .IN1(n1361), .IN2(n10049), .IN3(n1379), .IN4(n10050), .IN5(
        n10051), .Q(n9630) );
  AO22X1 U10299 ( .IN1(n1368), .IN2(n10052), .IN3(n1369), .IN4(n10053), .Q(
        n10051) );
  INVX0 U10300 ( .INP(n9629), .ZN(n9937) );
  AO221X1 U10301 ( .IN1(n1366), .IN2(n10054), .IN3(n1371), .IN4(n10055), .IN5(
        n10056), .Q(n9629) );
  AO22X1 U10302 ( .IN1(n1377), .IN2(n10057), .IN3(n1362), .IN4(n10058), .Q(
        n10056) );
  INVX0 U10303 ( .INP(n9633), .ZN(n9926) );
  AO222X1 U10304 ( .IN1(n1380), .IN2(n10059), .IN3(n10060), .IN4(n1033), .IN5(
        n1371), .IN6(n10061), .Q(n9633) );
  OA22X1 U10305 ( .IN1(n9601), .IN2(n9587), .IN3(n8944), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N21 ) );
  AO221X1 U10306 ( .IN1(n9703), .IN2(n9605), .IN3(n9702), .IN4(n9607), .IN5(
        n10062), .Q(n9587) );
  AO22X1 U10307 ( .IN1(n9609), .IN2(n9938), .IN3(n9602), .IN4(n9927), .Q(
        n10062) );
  INVX0 U10308 ( .INP(n9749), .ZN(n9927) );
  AO222X1 U10309 ( .IN1(n1369), .IN2(n10063), .IN3(n1379), .IN4(n9999), .IN5(
        n10064), .IN6(n1033), .Q(n9749) );
  INVX0 U10310 ( .INP(n9745), .ZN(n9938) );
  AO221X1 U10311 ( .IN1(n1372), .IN2(n10003), .IN3(n1377), .IN4(n10001), .IN5(
        n10065), .Q(n9745) );
  AO22X1 U10312 ( .IN1(n1365), .IN2(n10004), .IN3(n1364), .IN4(n9955), .Q(
        n10065) );
  INVX0 U10313 ( .INP(n9746), .ZN(n9702) );
  AO221X1 U10314 ( .IN1(n1371), .IN2(n10008), .IN3(n1378), .IN4(n10005), .IN5(
        n10066), .Q(n9746) );
  AO22X1 U10315 ( .IN1(n1366), .IN2(n10009), .IN3(n1363), .IN4(n9997), .Q(
        n10066) );
  INVX0 U10316 ( .INP(n9859), .ZN(n9703) );
  AO221X1 U10317 ( .IN1(n1378), .IN2(n9891), .IN3(n1369), .IN4(n9976), .IN5(
        n10067), .Q(n9859) );
  AO22X1 U10318 ( .IN1(n1361), .IN2(n10006), .IN3(n1368), .IN4(n10011), .Q(
        n10067) );
  AO221X1 U10319 ( .IN1(m4stg_frac[65]), .IN2(n1416), .IN3(m4stg_frac[66]), 
        .IN4(n1426), .IN5(n10068), .Q(n9891) );
  AO22X1 U10320 ( .IN1(m4stg_frac[67]), .IN2(n1437), .IN3(m4stg_frac[68]), 
        .IN4(n1443), .Q(n10068) );
  OA22X1 U10321 ( .IN1(n9601), .IN2(n9588), .IN3(n8938), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N20 ) );
  AO221X1 U10322 ( .IN1(n9609), .IN2(n9939), .IN3(n9602), .IN4(n9928), .IN5(
        n10069), .Q(n9588) );
  AO22X1 U10323 ( .IN1(n9713), .IN2(n9605), .IN3(n9714), .IN4(n9607), .Q(
        n10069) );
  INVX0 U10324 ( .INP(n9846), .ZN(n9714) );
  AO221X1 U10325 ( .IN1(n1370), .IN2(n10017), .IN3(n1380), .IN4(n10014), .IN5(
        n10070), .Q(n9846) );
  AO22X1 U10326 ( .IN1(n1364), .IN2(n10024), .IN3(n1365), .IN4(n10018), .Q(
        n10070) );
  INVX0 U10327 ( .INP(n9866), .ZN(n9713) );
  AO221X1 U10328 ( .IN1(n1377), .IN2(n9898), .IN3(n1370), .IN4(n9983), .IN5(
        n10071), .Q(n9866) );
  AO22X1 U10329 ( .IN1(n1362), .IN2(n10015), .IN3(n1366), .IN4(n10020), .Q(
        n10071) );
  AO221X1 U10330 ( .IN1(m4stg_frac[64]), .IN2(n1416), .IN3(m4stg_frac[65]), 
        .IN4(n1426), .IN5(n10072), .Q(n9898) );
  AO22X1 U10331 ( .IN1(m4stg_frac[66]), .IN2(n1437), .IN3(m4stg_frac[67]), 
        .IN4(n1443), .Q(n10072) );
  INVX0 U10332 ( .INP(n9843), .ZN(n9928) );
  AO222X1 U10333 ( .IN1(n1379), .IN2(n10022), .IN3(n1369), .IN4(n10073), .IN5(
        n10074), .IN6(n1033), .Q(n9843) );
  INVX0 U10334 ( .INP(n9842), .ZN(n9939) );
  AO222X1 U10335 ( .IN1(n1362), .IN2(n9622), .IN3(n1365), .IN4(n10075), .IN5(
        \fpu_mul_frac_dp/n765 ), .IN6(n10076), .Q(n9842) );
  OA22X1 U10336 ( .IN1(n9601), .IN2(n9589), .IN3(n8932), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N19 ) );
  AO221X1 U10337 ( .IN1(n9609), .IN2(n9953), .IN3(n9602), .IN4(n9946), .IN5(
        n10077), .Q(n9589) );
  AO22X1 U10338 ( .IN1(n9724), .IN2(n9605), .IN3(n9607), .IN4(n9725), .Q(
        n10077) );
  INVX0 U10339 ( .INP(n9874), .ZN(n9725) );
  AO221X1 U10340 ( .IN1(n1380), .IN2(n10033), .IN3(n1372), .IN4(n10032), .IN5(
        n10078), .Q(n9874) );
  AO22X1 U10341 ( .IN1(n1367), .IN2(n10029), .IN3(n1361), .IN4(n10039), .Q(
        n10078) );
  INVX0 U10342 ( .INP(n9870), .ZN(n9724) );
  AO221X1 U10343 ( .IN1(n1379), .IN2(n9905), .IN3(n1371), .IN4(n9990), .IN5(
        n10079), .Q(n9870) );
  AO22X1 U10344 ( .IN1(n1368), .IN2(n10035), .IN3(n1362), .IN4(n10030), .Q(
        n10079) );
  AO221X1 U10345 ( .IN1(m4stg_frac[63]), .IN2(n1416), .IN3(m4stg_frac[64]), 
        .IN4(n1427), .IN5(n10080), .Q(n9905) );
  AO22X1 U10346 ( .IN1(m4stg_frac[65]), .IN2(n1437), .IN3(m4stg_frac[66]), 
        .IN4(n1443), .Q(n10080) );
  INVX0 U10347 ( .INP(n9872), .ZN(n9946) );
  AO222X1 U10348 ( .IN1(n1364), .IN2(n10041), .IN3(\fpu_mul_frac_dp/n765 ), 
        .IN4(n10081), .IN5(n1368), .IN6(n10082), .Q(n9872) );
  AOI221X1 U10349 ( .IN1(n1363), .IN2(n10083), .IN3(n1367), .IN4(n10040), 
        .IN5(n10084), .QN(n9953) );
  AO22X1 U10350 ( .IN1(n1370), .IN2(n10043), .IN3(n1379), .IN4(n10044), .Q(
        n10084) );
  OA22X1 U10351 ( .IN1(n9601), .IN2(n9590), .IN3(n8926), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N18 ) );
  AO221X1 U10352 ( .IN1(n9735), .IN2(n10085), .IN3(n10086), .IN4(n9736), .IN5(
        n10087), .Q(n9590) );
  AO22X1 U10353 ( .IN1(n9602), .IN2(n10088), .IN3(n9609), .IN4(n9952), .Q(
        n10087) );
  AOI221X1 U10354 ( .IN1(n1368), .IN2(n10058), .IN3(n1362), .IN4(n10089), 
        .IN5(n10090), .QN(n9952) );
  AO22X1 U10355 ( .IN1(n1371), .IN2(n10054), .IN3(n1377), .IN4(n10055), .Q(
        n10090) );
  INVX0 U10356 ( .INP(n9882), .ZN(n10088) );
  AO222X1 U10357 ( .IN1(n1370), .IN2(n10091), .IN3(n1378), .IN4(n10061), .IN5(
        n10092), .IN6(n1033), .Q(n9882) );
  INVX0 U10358 ( .INP(n9883), .ZN(n9736) );
  AO221X1 U10359 ( .IN1(n1369), .IN2(n10052), .IN3(n1379), .IN4(n10053), .IN5(
        n10093), .Q(n9883) );
  AO22X1 U10360 ( .IN1(n1365), .IN2(n10049), .IN3(n1364), .IN4(n10059), .Q(
        n10093) );
  INVX0 U10361 ( .INP(n9880), .ZN(n9735) );
  AO221X1 U10362 ( .IN1(n1378), .IN2(n9911), .IN3(n1369), .IN4(n10048), .IN5(
        n10094), .Q(n9880) );
  AO22X1 U10363 ( .IN1(n1366), .IN2(n10046), .IN3(n1363), .IN4(n10050), .Q(
        n10094) );
  OA22X1 U10364 ( .IN1(n9601), .IN2(n9591), .IN3(n8920), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N17 ) );
  INVX0 U10365 ( .INP(n8927), .ZN(n8920) );
  AO221X1 U10366 ( .IN1(n9754), .IN2(n9605), .IN3(n9607), .IN4(n9753), .IN5(
        n10095), .Q(n9591) );
  AO22X1 U10367 ( .IN1(n9609), .IN2(n9968), .IN3(n9602), .IN4(n10096), .Q(
        n10095) );
  INVX0 U10368 ( .INP(n9888), .ZN(n10096) );
  AO222X1 U10369 ( .IN1(n1367), .IN2(n10000), .IN3(\fpu_mul_frac_dp/n765 ), 
        .IN4(n9998), .IN5(n1364), .IN6(n10001), .Q(n9888) );
  MUX21X1 U10370 ( .IN1(n10063), .IN2(n10097), .S(n906), .Q(n9998) );
  AOI221X1 U10371 ( .IN1(n1377), .IN2(n10003), .IN3(n1372), .IN4(n10004), 
        .IN5(n10098), .QN(n9968) );
  AO22X1 U10372 ( .IN1(n1367), .IN2(n9955), .IN3(n1361), .IN4(n9957), .Q(
        n10098) );
  INVX0 U10373 ( .INP(n9889), .ZN(n9753) );
  AO221X1 U10374 ( .IN1(n1365), .IN2(n9997), .IN3(n1370), .IN4(n10009), .IN5(
        n10099), .Q(n9889) );
  AO22X1 U10375 ( .IN1(n1379), .IN2(n10008), .IN3(n1362), .IN4(n9999), .Q(
        n10099) );
  INVX0 U10376 ( .INP(n9886), .ZN(n9754) );
  AO221X1 U10377 ( .IN1(n1377), .IN2(n9976), .IN3(n1372), .IN4(n10011), .IN5(
        n10100), .Q(n9886) );
  AO22X1 U10378 ( .IN1(n1368), .IN2(n10006), .IN3(n1364), .IN4(n10005), .Q(
        n10100) );
  AO221X1 U10379 ( .IN1(m4stg_frac[61]), .IN2(n1416), .IN3(m4stg_frac[62]), 
        .IN4(n1427), .IN5(n10101), .Q(n9976) );
  AO22X1 U10380 ( .IN1(m4stg_frac[63]), .IN2(n1437), .IN3(m4stg_frac[64]), 
        .IN4(n1443), .Q(n10101) );
  OA22X1 U10381 ( .IN1(n9601), .IN2(n9592), .IN3(n8914), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N16 ) );
  INVX0 U10382 ( .INP(n9025), .ZN(n8914) );
  AO221X1 U10383 ( .IN1(n9609), .IN2(n9967), .IN3(n9602), .IN4(n9944), .IN5(
        n10102), .Q(n9592) );
  AO22X1 U10384 ( .IN1(n10086), .IN2(n9764), .IN3(n9763), .IN4(n10085), .Q(
        n10102) );
  INVX0 U10385 ( .INP(n9893), .ZN(n9763) );
  AO221X1 U10386 ( .IN1(n1380), .IN2(n9983), .IN3(n1371), .IN4(n10020), .IN5(
        n10103), .Q(n9893) );
  AO22X1 U10387 ( .IN1(n1365), .IN2(n10015), .IN3(n1363), .IN4(n10014), .Q(
        n10103) );
  AO221X1 U10388 ( .IN1(m4stg_frac[60]), .IN2(n1416), .IN3(m4stg_frac[61]), 
        .IN4(n1427), .IN5(n10104), .Q(n9983) );
  AO22X1 U10389 ( .IN1(m4stg_frac[62]), .IN2(n1437), .IN3(m4stg_frac[63]), 
        .IN4(n1443), .Q(n10104) );
  INVX0 U10390 ( .INP(n9896), .ZN(n9764) );
  AO221X1 U10391 ( .IN1(n1364), .IN2(n10022), .IN3(n1369), .IN4(n10018), .IN5(
        n10105), .Q(n9896) );
  AO22X1 U10392 ( .IN1(n1380), .IN2(n10017), .IN3(n1367), .IN4(n10024), .Q(
        n10105) );
  INVX0 U10393 ( .INP(n9895), .ZN(n9944) );
  AO222X1 U10394 ( .IN1(n1363), .IN2(n10025), .IN3(\fpu_mul_frac_dp/n765 ), 
        .IN4(n10023), .IN5(n1367), .IN6(n10027), .Q(n9895) );
  MUX21X1 U10395 ( .IN1(n10073), .IN2(n10106), .S(n906), .Q(n10023) );
  AOI222X1 U10396 ( .IN1(n1363), .IN2(n9621), .IN3(\fpu_mul_frac_dp/n765 ), 
        .IN4(n10026), .IN5(n1368), .IN6(n9622), .QN(n9967) );
  MUX21X1 U10397 ( .IN1(n10107), .IN2(n10075), .S(n906), .Q(n10026) );
  OA22X1 U10398 ( .IN1(n9601), .IN2(n9593), .IN3(n8908), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N15 ) );
  AO221X1 U10399 ( .IN1(n9609), .IN2(n9966), .IN3(n9602), .IN4(n9943), .IN5(
        n10108), .Q(n9593) );
  AO22X1 U10400 ( .IN1(n9773), .IN2(n9605), .IN3(n9607), .IN4(n9774), .Q(
        n10108) );
  INVX0 U10401 ( .INP(n9903), .ZN(n9774) );
  AO221X1 U10402 ( .IN1(n1370), .IN2(n10029), .IN3(n1377), .IN4(n10032), .IN5(
        n10109), .Q(n9903) );
  AO22X1 U10403 ( .IN1(n1366), .IN2(n10039), .IN3(n1361), .IN4(n10037), .Q(
        n10109) );
  INVX0 U10404 ( .INP(n9900), .ZN(n9773) );
  AO221X1 U10405 ( .IN1(n1368), .IN2(n10030), .IN3(n1361), .IN4(n10033), .IN5(
        n10110), .Q(n9900) );
  AO22X1 U10406 ( .IN1(n1372), .IN2(n10035), .IN3(n1378), .IN4(n9990), .Q(
        n10110) );
  AO221X1 U10407 ( .IN1(m4stg_frac[59]), .IN2(n1416), .IN3(m4stg_frac[60]), 
        .IN4(n1427), .IN5(n10111), .Q(n9990) );
  AO22X1 U10408 ( .IN1(m4stg_frac[61]), .IN2(n1437), .IN3(m4stg_frac[62]), 
        .IN4(n1443), .Q(n10111) );
  INVX0 U10409 ( .INP(n9902), .ZN(n9943) );
  AO222X1 U10410 ( .IN1(n1368), .IN2(n10041), .IN3(\fpu_mul_frac_dp/n765 ), 
        .IN4(n10038), .IN5(n1363), .IN6(n10044), .Q(n9902) );
  MUX21X1 U10411 ( .IN1(n10112), .IN2(n10082), .S(n906), .Q(n10038) );
  AOI222X1 U10412 ( .IN1(n1379), .IN2(n10043), .IN3(n9624), .IN4(n1033), .IN5(
        n1371), .IN6(n10040), .QN(n9966) );
  MUX21X1 U10413 ( .IN1(n9970), .IN2(n10083), .S(\fpu_mul_frac_dp/n833 ), .Q(
        n9624) );
  OA22X1 U10414 ( .IN1(n9601), .IN2(n9594), .IN3(n8902), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N14 ) );
  AO221X1 U10415 ( .IN1(n9609), .IN2(n9965), .IN3(n9602), .IN4(n9942), .IN5(
        n10113), .Q(n9594) );
  AO22X1 U10416 ( .IN1(n10086), .IN2(n9784), .IN3(n9783), .IN4(n10085), .Q(
        n10113) );
  INVX0 U10417 ( .INP(n9907), .ZN(n9783) );
  AO221X1 U10418 ( .IN1(n1365), .IN2(n10050), .IN3(n1364), .IN4(n10053), .IN5(
        n10114), .Q(n9907) );
  AO22X1 U10419 ( .IN1(n1371), .IN2(n10046), .IN3(n1380), .IN4(n10048), .Q(
        n10114) );
  INVX0 U10420 ( .INP(n9910), .ZN(n9784) );
  AO221X1 U10421 ( .IN1(n1363), .IN2(n10061), .IN3(n1380), .IN4(n10052), .IN5(
        n10115), .Q(n9910) );
  AO22X1 U10422 ( .IN1(n1372), .IN2(n10049), .IN3(n1368), .IN4(n10059), .Q(
        n10115) );
  INVX0 U10423 ( .INP(n9909), .ZN(n9942) );
  AO222X1 U10424 ( .IN1(n1365), .IN2(n10057), .IN3(\fpu_mul_frac_dp/n765 ), 
        .IN4(n10060), .IN5(n1362), .IN6(n10055), .Q(n9909) );
  MUX21X1 U10425 ( .IN1(n10091), .IN2(n10116), .S(n906), .Q(n10060) );
  AOI222X1 U10426 ( .IN1(n1378), .IN2(n10054), .IN3(n9632), .IN4(n1033), .IN5(
        n1369), .IN6(n10058), .QN(n9965) );
  INVX0 U10427 ( .INP(n9959), .ZN(n9632) );
  MUX21X1 U10428 ( .IN1(n10117), .IN2(n10118), .S(\fpu_mul_frac_dp/n833 ), .Q(
        n9959) );
  INVX0 U10429 ( .INP(n10089), .ZN(n10118) );
  NAND2X0 U10430 ( .IN1(\fpu_mul_frac_dp/n834 ), .IN2(n10119), .QN(n10117) );
  OA22X1 U10431 ( .IN1(n9601), .IN2(n9595), .IN3(n8896), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N13 ) );
  AO221X1 U10432 ( .IN1(n9609), .IN2(n9964), .IN3(n9602), .IN4(n9941), .IN5(
        n10120), .Q(n9595) );
  AO22X1 U10433 ( .IN1(n9795), .IN2(n9605), .IN3(n9607), .IN4(n9796), .Q(
        n10120) );
  INVX0 U10434 ( .INP(n9974), .ZN(n9796) );
  AO221X1 U10435 ( .IN1(n1368), .IN2(n9999), .IN3(n1363), .IN4(n10063), .IN5(
        n10121), .Q(n9974) );
  AO22X1 U10436 ( .IN1(n1378), .IN2(n10009), .IN3(n1370), .IN4(n9997), .Q(
        n10121) );
  AO221X1 U10437 ( .IN1(m4stg_frac[37]), .IN2(n1416), .IN3(m4stg_frac[38]), 
        .IN4(n1427), .IN5(n10122), .Q(n9997) );
  AO22X1 U10438 ( .IN1(m4stg_frac[39]), .IN2(n1437), .IN3(m4stg_frac[40]), 
        .IN4(n1443), .Q(n10122) );
  AO221X1 U10439 ( .IN1(m4stg_frac[41]), .IN2(n1416), .IN3(m4stg_frac[42]), 
        .IN4(n1427), .IN5(n10123), .Q(n10009) );
  AO22X1 U10440 ( .IN1(m4stg_frac[43]), .IN2(n1437), .IN3(m4stg_frac[44]), 
        .IN4(n1443), .Q(n10123) );
  AO222X1 U10441 ( .IN1(m4stg_frac[32]), .IN2(n1446), .IN3(n9384), .IN4(n879), 
        .IN5(m4stg_frac[31]), .IN6(n1431), .Q(n10063) );
  AO221X1 U10442 ( .IN1(m4stg_frac[33]), .IN2(n1416), .IN3(m4stg_frac[34]), 
        .IN4(n1427), .IN5(n10124), .Q(n9999) );
  AO22X1 U10443 ( .IN1(m4stg_frac[35]), .IN2(n1437), .IN3(m4stg_frac[36]), 
        .IN4(n1443), .Q(n10124) );
  INVX0 U10444 ( .INP(n9971), .ZN(n9795) );
  AO221X1 U10445 ( .IN1(n1379), .IN2(n10011), .IN3(n1370), .IN4(n10006), .IN5(
        n10125), .Q(n9971) );
  AO22X1 U10446 ( .IN1(n1367), .IN2(n10005), .IN3(n1362), .IN4(n10008), .Q(
        n10125) );
  AO222X1 U10447 ( .IN1(m4stg_frac[45]), .IN2(n1419), .IN3(
        \fpu_mul_frac_dp/n834 ), .IN4(n9381), .IN5(m4stg_frac[46]), .IN6(n1430), .Q(n10008) );
  AO221X1 U10448 ( .IN1(m4stg_frac[49]), .IN2(n1417), .IN3(m4stg_frac[50]), 
        .IN4(n1427), .IN5(n10126), .Q(n10005) );
  AO22X1 U10449 ( .IN1(m4stg_frac[51]), .IN2(n1437), .IN3(m4stg_frac[52]), 
        .IN4(n1443), .Q(n10126) );
  AO221X1 U10450 ( .IN1(m4stg_frac[53]), .IN2(n1417), .IN3(m4stg_frac[54]), 
        .IN4(n1427), .IN5(n10127), .Q(n10006) );
  AO22X1 U10451 ( .IN1(m4stg_frac[55]), .IN2(n1437), .IN3(m4stg_frac[56]), 
        .IN4(n1444), .Q(n10127) );
  AO221X1 U10452 ( .IN1(m4stg_frac[57]), .IN2(n1417), .IN3(m4stg_frac[58]), 
        .IN4(n1427), .IN5(n10128), .Q(n10011) );
  AO22X1 U10453 ( .IN1(m4stg_frac[59]), .IN2(n1437), .IN3(m4stg_frac[60]), 
        .IN4(n1443), .Q(n10128) );
  INVX0 U10454 ( .INP(n9973), .ZN(n9941) );
  AO222X1 U10455 ( .IN1(n1361), .IN2(n10003), .IN3(\fpu_mul_frac_dp/n765 ), 
        .IN4(n10064), .IN5(n1366), .IN6(n10001), .Q(n9973) );
  AO222X1 U10456 ( .IN1(m4stg_frac[20]), .IN2(n1446), .IN3(n9387), .IN4(n879), 
        .IN5(m4stg_frac[19]), .IN6(n1432), .Q(n10001) );
  MUX21X1 U10457 ( .IN1(n10097), .IN2(n10000), .S(n906), .Q(n10064) );
  AO222X1 U10458 ( .IN1(m4stg_frac[24]), .IN2(n1446), .IN3(n9385), .IN4(n879), 
        .IN5(m4stg_frac[23]), .IN6(n1431), .Q(n10000) );
  MUX21X1 U10459 ( .IN1(n9383), .IN2(n9386), .S(n879), .Q(n10097) );
  AO222X1 U10460 ( .IN1(m4stg_frac[16]), .IN2(n1447), .IN3(n9388), .IN4(n879), 
        .IN5(m4stg_frac[15]), .IN6(n1432), .Q(n10003) );
  AOI222X1 U10461 ( .IN1(n1380), .IN2(n10004), .IN3(n9748), .IN4(n1033), .IN5(
        n1370), .IN6(n9955), .QN(n9964) );
  AO221X1 U10462 ( .IN1(m4stg_frac[5]), .IN2(n1417), .IN3(m4stg_frac[6]), 
        .IN4(n1428), .IN5(n10129), .Q(n9955) );
  AO22X1 U10463 ( .IN1(m4stg_frac[7]), .IN2(n1437), .IN3(m4stg_frac[8]), .IN4(
        n1444), .Q(n10129) );
  INVX0 U10464 ( .INP(n9958), .ZN(n9748) );
  MUX21X1 U10465 ( .IN1(n10130), .IN2(n10131), .S(\fpu_mul_frac_dp/n833 ), .Q(
        n9958) );
  INVX0 U10466 ( .INP(n9957), .ZN(n10131) );
  AO221X1 U10467 ( .IN1(m4stg_frac[1]), .IN2(n1417), .IN3(m4stg_frac[2]), 
        .IN4(n1427), .IN5(n10132), .Q(n9957) );
  AO22X1 U10468 ( .IN1(m4stg_frac[3]), .IN2(n1437), .IN3(m4stg_frac[4]), .IN4(
        n1444), .Q(n10132) );
  NAND2X0 U10469 ( .IN1(m4stg_frac[0]), .IN2(n1447), .QN(n10130) );
  AO221X1 U10470 ( .IN1(m4stg_frac[9]), .IN2(n1417), .IN3(m4stg_frac[10]), 
        .IN4(n1428), .IN5(n10133), .Q(n10004) );
  AO22X1 U10471 ( .IN1(m4stg_frac[11]), .IN2(n1437), .IN3(m4stg_frac[12]), 
        .IN4(n1444), .Q(n10133) );
  OA22X1 U10472 ( .IN1(n9601), .IN2(n9596), .IN3(n8890), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N12 ) );
  INVX0 U10473 ( .INP(n9027), .ZN(n8890) );
  AO221X1 U10474 ( .IN1(n9609), .IN2(n9963), .IN3(n9602), .IN4(n9945), .IN5(
        n10134), .Q(n9596) );
  AO22X1 U10475 ( .IN1(n10086), .IN2(n9806), .IN3(n9805), .IN4(n10085), .Q(
        n10134) );
  NOR2X0 U10476 ( .IN1(n9876), .IN2(n908), .QN(n10085) );
  INVX0 U10477 ( .INP(n9978), .ZN(n9805) );
  AO221X1 U10478 ( .IN1(n1378), .IN2(n10020), .IN3(n1372), .IN4(n10015), .IN5(
        n10135), .Q(n9978) );
  AO22X1 U10479 ( .IN1(n1368), .IN2(n10014), .IN3(n1364), .IN4(n10017), .Q(
        n10135) );
  AO222X1 U10480 ( .IN1(m4stg_frac[44]), .IN2(n1420), .IN3(
        \fpu_mul_frac_dp/n834 ), .IN4(n9382), .IN5(m4stg_frac[45]), .IN6(n1430), .Q(n10017) );
  AO221X1 U10481 ( .IN1(m4stg_frac[48]), .IN2(n1417), .IN3(m4stg_frac[49]), 
        .IN4(n1428), .IN5(n10136), .Q(n10014) );
  AO22X1 U10482 ( .IN1(m4stg_frac[50]), .IN2(n1438), .IN3(m4stg_frac[51]), 
        .IN4(n1444), .Q(n10136) );
  AO221X1 U10483 ( .IN1(m4stg_frac[52]), .IN2(n1417), .IN3(m4stg_frac[53]), 
        .IN4(n1428), .IN5(n10137), .Q(n10015) );
  AO22X1 U10484 ( .IN1(m4stg_frac[54]), .IN2(n1438), .IN3(m4stg_frac[55]), 
        .IN4(n1444), .Q(n10137) );
  AO221X1 U10485 ( .IN1(m4stg_frac[56]), .IN2(n1417), .IN3(m4stg_frac[57]), 
        .IN4(n1428), .IN5(n10138), .Q(n10020) );
  AO22X1 U10486 ( .IN1(m4stg_frac[58]), .IN2(n1438), .IN3(m4stg_frac[59]), 
        .IN4(n1444), .Q(n10138) );
  INVX0 U10487 ( .INP(n9981), .ZN(n9806) );
  AO221X1 U10488 ( .IN1(n1377), .IN2(n10018), .IN3(n1371), .IN4(n10024), .IN5(
        n10139), .Q(n9981) );
  AO22X1 U10489 ( .IN1(n1366), .IN2(n10022), .IN3(n1363), .IN4(n10073), .Q(
        n10139) );
  AO222X1 U10490 ( .IN1(m4stg_frac[28]), .IN2(n1420), .IN3(
        \fpu_mul_frac_dp/n834 ), .IN4(n9389), .IN5(m4stg_frac[29]), .IN6(n1430), .Q(n10073) );
  AO221X1 U10491 ( .IN1(m4stg_frac[32]), .IN2(n1417), .IN3(m4stg_frac[33]), 
        .IN4(n1428), .IN5(n10140), .Q(n10022) );
  AO22X1 U10492 ( .IN1(m4stg_frac[34]), .IN2(n1438), .IN3(m4stg_frac[35]), 
        .IN4(n1444), .Q(n10140) );
  AO221X1 U10493 ( .IN1(m4stg_frac[36]), .IN2(n1417), .IN3(m4stg_frac[37]), 
        .IN4(n1428), .IN5(n10141), .Q(n10024) );
  AO22X1 U10494 ( .IN1(m4stg_frac[38]), .IN2(n1438), .IN3(m4stg_frac[39]), 
        .IN4(n1444), .Q(n10141) );
  AO221X1 U10495 ( .IN1(m4stg_frac[40]), .IN2(n1417), .IN3(m4stg_frac[41]), 
        .IN4(n1428), .IN5(n10142), .Q(n10018) );
  AO22X1 U10496 ( .IN1(m4stg_frac[42]), .IN2(n1438), .IN3(m4stg_frac[43]), 
        .IN4(n1444), .Q(n10142) );
  NOR2X0 U10497 ( .IN1(n9876), .IN2(\fpu_mul_frac_dp/n838 ), .QN(n10086) );
  INVX0 U10498 ( .INP(n9980), .ZN(n9945) );
  MUX21X1 U10499 ( .IN1(n10076), .IN2(n10074), .S(\fpu_mul_frac_dp/n765 ), .Q(
        n9980) );
  MUX21X1 U10500 ( .IN1(n10106), .IN2(n10027), .S(n906), .Q(n10074) );
  AO222X1 U10501 ( .IN1(m4stg_frac[20]), .IN2(n1420), .IN3(
        \fpu_mul_frac_dp/n834 ), .IN4(n9391), .IN5(m4stg_frac[21]), .IN6(n1430), .Q(n10027) );
  MUX21X1 U10502 ( .IN1(n9390), .IN2(n9392), .S(n879), .Q(n10106) );
  MUX21X1 U10503 ( .IN1(n10107), .IN2(n10025), .S(\fpu_mul_frac_dp/n833 ), .Q(
        n10076) );
  AO222X1 U10504 ( .IN1(m4stg_frac[16]), .IN2(n1420), .IN3(
        \fpu_mul_frac_dp/n834 ), .IN4(n9393), .IN5(m4stg_frac[17]), .IN6(n1430), .Q(n10025) );
  MUX21X1 U10505 ( .IN1(n9395), .IN2(n9394), .S(n879), .Q(n10107) );
  AOI222X1 U10506 ( .IN1(n1377), .IN2(n10075), .IN3(n1367), .IN4(n9621), .IN5(
        n1372), .IN6(n9622), .QN(n9963) );
  AO221X1 U10507 ( .IN1(m4stg_frac[4]), .IN2(n1418), .IN3(m4stg_frac[5]), 
        .IN4(n1428), .IN5(n10143), .Q(n9622) );
  AO22X1 U10508 ( .IN1(m4stg_frac[6]), .IN2(n1438), .IN3(m4stg_frac[7]), .IN4(
        n1444), .Q(n10143) );
  AO222X1 U10509 ( .IN1(m4stg_frac[3]), .IN2(n1447), .IN3(n10119), .IN4(n879), 
        .IN5(m4stg_frac[2]), .IN6(n1431), .Q(n9621) );
  AO221X1 U10510 ( .IN1(m4stg_frac[8]), .IN2(n1417), .IN3(m4stg_frac[9]), 
        .IN4(n1429), .IN5(n10144), .Q(n10075) );
  AO22X1 U10511 ( .IN1(m4stg_frac[10]), .IN2(n1438), .IN3(m4stg_frac[11]), 
        .IN4(n1445), .Q(n10144) );
  OA22X1 U10512 ( .IN1(n9601), .IN2(n9597), .IN3(n8884), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N11 ) );
  INVX0 U10513 ( .INP(n8891), .ZN(n8884) );
  AO221X1 U10514 ( .IN1(n9609), .IN2(n9962), .IN3(n9602), .IN4(n9940), .IN5(
        n10145), .Q(n9597) );
  AO22X1 U10515 ( .IN1(n9815), .IN2(n9605), .IN3(n9607), .IN4(n9816), .Q(
        n10145) );
  INVX0 U10516 ( .INP(n9988), .ZN(n9816) );
  AO222X1 U10517 ( .IN1(n1372), .IN2(n10039), .IN3(n10081), .IN4(n1033), .IN5(
        n1380), .IN6(n10029), .Q(n9988) );
  AO221X1 U10518 ( .IN1(m4stg_frac[39]), .IN2(n1418), .IN3(m4stg_frac[40]), 
        .IN4(n1428), .IN5(n10146), .Q(n10029) );
  AO22X1 U10519 ( .IN1(m4stg_frac[41]), .IN2(n1438), .IN3(m4stg_frac[42]), 
        .IN4(n1444), .Q(n10146) );
  MUX21X1 U10520 ( .IN1(n10037), .IN2(n10112), .S(n906), .Q(n10081) );
  MUX21X1 U10521 ( .IN1(n9384), .IN2(n9383), .S(n879), .Q(n10112) );
  MUX21X1 U10522 ( .IN1(m4stg_frac[28]), .IN2(m4stg_frac[27]), .S(n884), .Q(
        n9383) );
  MUX21X1 U10523 ( .IN1(m4stg_frac[29]), .IN2(m4stg_frac[30]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9384) );
  AO221X1 U10524 ( .IN1(m4stg_frac[31]), .IN2(n1417), .IN3(m4stg_frac[32]), 
        .IN4(n1429), .IN5(n10147), .Q(n10037) );
  AO22X1 U10525 ( .IN1(m4stg_frac[33]), .IN2(n1438), .IN3(m4stg_frac[34]), 
        .IN4(n1445), .Q(n10147) );
  AO221X1 U10526 ( .IN1(m4stg_frac[35]), .IN2(n1418), .IN3(m4stg_frac[36]), 
        .IN4(n1428), .IN5(n10148), .Q(n10039) );
  AO22X1 U10527 ( .IN1(m4stg_frac[37]), .IN2(n1438), .IN3(m4stg_frac[38]), 
        .IN4(n1444), .Q(n10148) );
  NOR2X0 U10528 ( .IN1(n9696), .IN2(se_mul), .QN(n9607) );
  AND2X1 U10529 ( .IN1(n9619), .IN2(n1357), .Q(n9605) );
  INVX0 U10530 ( .INP(n9985), .ZN(n9815) );
  AO221X1 U10531 ( .IN1(n1362), .IN2(n10032), .IN3(n1367), .IN4(n10033), .IN5(
        n10149), .Q(n9985) );
  AO22X1 U10532 ( .IN1(n1377), .IN2(n10035), .IN3(n1372), .IN4(n10030), .Q(
        n10149) );
  AO221X1 U10533 ( .IN1(m4stg_frac[51]), .IN2(n1418), .IN3(m4stg_frac[52]), 
        .IN4(n1429), .IN5(n10150), .Q(n10030) );
  AO22X1 U10534 ( .IN1(m4stg_frac[53]), .IN2(n1438), .IN3(m4stg_frac[54]), 
        .IN4(n1445), .Q(n10150) );
  AO221X1 U10535 ( .IN1(m4stg_frac[55]), .IN2(n1418), .IN3(m4stg_frac[56]), 
        .IN4(n1427), .IN5(n10151), .Q(n10035) );
  AO22X1 U10536 ( .IN1(m4stg_frac[57]), .IN2(n1438), .IN3(m4stg_frac[58]), 
        .IN4(n1444), .Q(n10151) );
  AO222X1 U10537 ( .IN1(m4stg_frac[50]), .IN2(n1446), .IN3(n9381), .IN4(n879), 
        .IN5(m4stg_frac[49]), .IN6(n1431), .Q(n10033) );
  MUX21X1 U10538 ( .IN1(m4stg_frac[47]), .IN2(m4stg_frac[48]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9381) );
  AO221X1 U10539 ( .IN1(m4stg_frac[43]), .IN2(n1418), .IN3(m4stg_frac[44]), 
        .IN4(n1429), .IN5(n10152), .Q(n10032) );
  AO22X1 U10540 ( .IN1(m4stg_frac[45]), .IN2(n1438), .IN3(m4stg_frac[46]), 
        .IN4(n1444), .Q(n10152) );
  INVX0 U10541 ( .INP(n9987), .ZN(n9940) );
  AO221X1 U10542 ( .IN1(n1369), .IN2(n10041), .IN3(n1379), .IN4(n10082), .IN5(
        n10153), .Q(n9987) );
  AO22X1 U10543 ( .IN1(n1364), .IN2(n10043), .IN3(n1365), .IN4(n10044), .Q(
        n10153) );
  AO222X1 U10544 ( .IN1(m4stg_frac[15]), .IN2(n1420), .IN3(
        \fpu_mul_frac_dp/n834 ), .IN4(n9387), .IN5(m4stg_frac[16]), .IN6(n1430), .Q(n10044) );
  MUX21X1 U10545 ( .IN1(m4stg_frac[17]), .IN2(m4stg_frac[18]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9387) );
  AO222X1 U10546 ( .IN1(m4stg_frac[11]), .IN2(n1420), .IN3(
        \fpu_mul_frac_dp/n834 ), .IN4(n9388), .IN5(m4stg_frac[12]), .IN6(n1430), .Q(n10043) );
  MUX21X1 U10547 ( .IN1(m4stg_frac[13]), .IN2(m4stg_frac[14]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9388) );
  AO222X1 U10548 ( .IN1(m4stg_frac[23]), .IN2(n1420), .IN3(
        \fpu_mul_frac_dp/n834 ), .IN4(n9386), .IN5(m4stg_frac[24]), .IN6(n1430), .Q(n10082) );
  MUX21X1 U10549 ( .IN1(m4stg_frac[26]), .IN2(m4stg_frac[25]), .S(n884), .Q(
        n9386) );
  AO222X1 U10550 ( .IN1(m4stg_frac[19]), .IN2(n1420), .IN3(
        \fpu_mul_frac_dp/n834 ), .IN4(n9385), .IN5(m4stg_frac[20]), .IN6(n1430), .Q(n10041) );
  MUX21X1 U10551 ( .IN1(m4stg_frac[22]), .IN2(m4stg_frac[21]), .S(n884), .Q(
        n9385) );
  AOI222X1 U10552 ( .IN1(n1378), .IN2(n10040), .IN3(n1365), .IN4(n9970), .IN5(
        n1371), .IN6(n10083), .QN(n9962) );
  AO221X1 U10553 ( .IN1(m4stg_frac[3]), .IN2(n1418), .IN3(m4stg_frac[4]), 
        .IN4(n1429), .IN5(n10154), .Q(n10083) );
  AO22X1 U10554 ( .IN1(m4stg_frac[5]), .IN2(n1438), .IN3(m4stg_frac[6]), .IN4(
        n1445), .Q(n10154) );
  AO222X1 U10555 ( .IN1(m4stg_frac[2]), .IN2(n1447), .IN3(m4stg_frac[0]), 
        .IN4(n1427), .IN5(m4stg_frac[1]), .IN6(n1431), .Q(n9970) );
  AO221X1 U10556 ( .IN1(m4stg_frac[7]), .IN2(n1418), .IN3(m4stg_frac[8]), 
        .IN4(n9347), .IN5(n10155), .Q(n10040) );
  AO22X1 U10557 ( .IN1(m4stg_frac[9]), .IN2(n1433), .IN3(m4stg_frac[10]), 
        .IN4(n1444), .Q(n10155) );
  OA22X1 U10558 ( .IN1(n9601), .IN2(n9598), .IN3(n8878), .IN4(n2929), .Q(
        \fpu_mul_frac_dp/i_m5stg_frac_pre1/N10 ) );
  INVX0 U10559 ( .INP(n9028), .ZN(n8878) );
  AO222X1 U10560 ( .IN1(n10156), .IN2(n10157), .IN3(n9609), .IN4(n9961), .IN5(
        n9602), .IN6(n9934), .Q(n9598) );
  AOI222X1 U10561 ( .IN1(n1361), .IN2(n10054), .IN3(\fpu_mul_frac_dp/n765 ), 
        .IN4(n10092), .IN5(n1367), .IN6(n10055), .QN(n9934) );
  AO222X1 U10562 ( .IN1(m4stg_frac[17]), .IN2(n1447), .IN3(n9395), .IN4(n879), 
        .IN5(m4stg_frac[16]), .IN6(n1431), .Q(n10055) );
  MUX21X1 U10563 ( .IN1(m4stg_frac[14]), .IN2(m4stg_frac[15]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9395) );
  MUX21X1 U10564 ( .IN1(n10116), .IN2(n10057), .S(n906), .Q(n10092) );
  AO222X1 U10565 ( .IN1(m4stg_frac[21]), .IN2(n1446), .IN3(n9393), .IN4(n879), 
        .IN5(m4stg_frac[20]), .IN6(n1432), .Q(n10057) );
  MUX21X1 U10566 ( .IN1(m4stg_frac[18]), .IN2(m4stg_frac[19]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9393) );
  MUX21X1 U10567 ( .IN1(n9392), .IN2(n9391), .S(n879), .Q(n10116) );
  MUX21X1 U10568 ( .IN1(m4stg_frac[22]), .IN2(m4stg_frac[23]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9391) );
  MUX21X1 U10569 ( .IN1(m4stg_frac[24]), .IN2(m4stg_frac[25]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9392) );
  AO222X1 U10570 ( .IN1(m4stg_frac[10]), .IN2(n1420), .IN3(
        \fpu_mul_frac_dp/n834 ), .IN4(n9394), .IN5(m4stg_frac[11]), .IN6(n1430), .Q(n10054) );
  MUX21X1 U10571 ( .IN1(m4stg_frac[12]), .IN2(m4stg_frac[13]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9394) );
  NOR2X0 U10572 ( .IN1(n9654), .IN2(se_mul), .QN(n9602) );
  AOI222X1 U10573 ( .IN1(n1380), .IN2(n10058), .IN3(n10158), .IN4(n1366), 
        .IN5(n1370), .IN6(n10089), .QN(n9961) );
  AO221X1 U10574 ( .IN1(m4stg_frac[2]), .IN2(n1418), .IN3(m4stg_frac[3]), 
        .IN4(n9347), .IN5(n10159), .Q(n10089) );
  AO22X1 U10575 ( .IN1(m4stg_frac[4]), .IN2(n1438), .IN3(m4stg_frac[5]), .IN4(
        n1445), .Q(n10159) );
  AND2X1 U10576 ( .IN1(n10119), .IN2(\fpu_mul_frac_dp/n834 ), .Q(n10158) );
  MUX21X1 U10577 ( .IN1(m4stg_frac[0]), .IN2(m4stg_frac[1]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n10119) );
  AO221X1 U10578 ( .IN1(m4stg_frac[6]), .IN2(n1419), .IN3(m4stg_frac[7]), 
        .IN4(n1429), .IN5(n10160), .Q(n10058) );
  AO22X1 U10579 ( .IN1(m4stg_frac[8]), .IN2(n1437), .IN3(m4stg_frac[9]), .IN4(
        n1445), .Q(n10160) );
  NOR2X0 U10580 ( .IN1(n9655), .IN2(se_mul), .QN(n9609) );
  INVX0 U10581 ( .INP(n9824), .ZN(n10157) );
  MUX21X1 U10582 ( .IN1(n9995), .IN2(n10161), .S(\fpu_mul_frac_dp/n838 ), .Q(
        n9824) );
  AO221X1 U10583 ( .IN1(n1361), .IN2(n10091), .IN3(n1368), .IN4(n10061), .IN5(
        n10162), .Q(n9995) );
  AO22X1 U10584 ( .IN1(n1379), .IN2(n10049), .IN3(n1371), .IN4(n10059), .Q(
        n10162) );
  AO221X1 U10585 ( .IN1(m4stg_frac[34]), .IN2(n1418), .IN3(m4stg_frac[35]), 
        .IN4(n9347), .IN5(n10163), .Q(n10059) );
  AO22X1 U10586 ( .IN1(m4stg_frac[36]), .IN2(n9349), .IN3(m4stg_frac[37]), 
        .IN4(n1445), .Q(n10163) );
  AO221X1 U10587 ( .IN1(m4stg_frac[38]), .IN2(n1419), .IN3(m4stg_frac[39]), 
        .IN4(n1429), .IN5(n10164), .Q(n10049) );
  AO22X1 U10588 ( .IN1(m4stg_frac[40]), .IN2(n9349), .IN3(m4stg_frac[41]), 
        .IN4(n1445), .Q(n10164) );
  AO222X1 U10589 ( .IN1(m4stg_frac[33]), .IN2(n1447), .IN3(n9389), .IN4(n879), 
        .IN5(m4stg_frac[32]), .IN6(n1431), .Q(n10061) );
  MUX21X1 U10590 ( .IN1(m4stg_frac[30]), .IN2(m4stg_frac[31]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9389) );
  AO222X1 U10591 ( .IN1(m4stg_frac[29]), .IN2(n1447), .IN3(n9390), .IN4(n879), 
        .IN5(m4stg_frac[28]), .IN6(n1431), .Q(n10091) );
  MUX21X1 U10592 ( .IN1(m4stg_frac[26]), .IN2(m4stg_frac[27]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9390) );
  INVX0 U10593 ( .INP(n9876), .ZN(n10156) );
  NAND2X0 U10594 ( .IN1(\fpu_mul_frac_dp/n766 ), .IN2(n1359), .QN(n9876) );
  OA21X1 U10595 ( .IN1(n9600), .IN2(n10165), .IN3(n1357), .Q(n9601) );
  INVX0 U10596 ( .INP(m4stg_shl_55), .ZN(n10165) );
  NAND4X0 U10597 ( .IN1(n10166), .IN2(n10167), .IN3(n10168), .IN4(n10169), 
        .QN(m4stg_shl_55) );
  OA22X1 U10598 ( .IN1(n10170), .IN2(n10171), .IN3(n9691), .IN4(n9648), .Q(
        n10169) );
  NAND2X0 U10599 ( .IN1(n10172), .IN2(\fpu_mul_frac_dp/n833 ), .QN(n9648) );
  INVX0 U10600 ( .INP(n9743), .ZN(n9691) );
  AO221X1 U10601 ( .IN1(m4stg_frac[94]), .IN2(n1418), .IN3(m4stg_frac[95]), 
        .IN4(n9347), .IN5(n10173), .Q(n9743) );
  AO22X1 U10602 ( .IN1(m4stg_frac[96]), .IN2(n9349), .IN3(m4stg_frac[97]), 
        .IN4(n1445), .Q(n10173) );
  INVX0 U10603 ( .INP(n9742), .ZN(n10171) );
  NOR2X0 U10604 ( .IN1(n906), .IN2(n10174), .QN(n9742) );
  AOI22X1 U10605 ( .IN1(n879), .IN2(n9663), .IN3(n1432), .IN4(m4stg_frac[104]), 
        .QN(n10170) );
  MUX21X1 U10606 ( .IN1(m4stg_frac[103]), .IN2(m4stg_frac[102]), .S(n884), .Q(
        n9663) );
  OA22X1 U10607 ( .IN1(n10174), .IN2(n9459), .IN3(n10175), .IN4(n9646), .Q(
        n10168) );
  OR2X1 U10608 ( .IN1(n10174), .IN2(\fpu_mul_frac_dp/n833 ), .Q(n9646) );
  INVX0 U10609 ( .INP(n9698), .ZN(n10175) );
  AO221X1 U10610 ( .IN1(m4stg_frac[98]), .IN2(n1419), .IN3(m4stg_frac[99]), 
        .IN4(n1428), .IN5(n10176), .Q(n9698) );
  AO22X1 U10611 ( .IN1(m4stg_frac[100]), .IN2(n9349), .IN3(m4stg_frac[101]), 
        .IN4(n1445), .Q(n10176) );
  NAND3X0 U10612 ( .IN1(n1439), .IN2(\fpu_mul_frac_dp/n833 ), .IN3(
        m4stg_frac_105), .QN(n9459) );
  NAND2X0 U10613 ( .IN1(\fpu_mul_frac_dp/n765 ), .IN2(n9619), .QN(n10174) );
  AOI22X1 U10614 ( .IN1(n9825), .IN2(n9614), .IN3(n9739), .IN4(n9651), .QN(
        n10167) );
  INVX0 U10615 ( .INP(n9693), .ZN(n9651) );
  NAND2X0 U10616 ( .IN1(n10172), .IN2(n906), .QN(n9693) );
  AND2X1 U10617 ( .IN1(n9619), .IN2(n1033), .Q(n10172) );
  NOR2X0 U10618 ( .IN1(n908), .IN2(n1035), .QN(n9619) );
  AO221X1 U10619 ( .IN1(m4stg_frac[90]), .IN2(n1418), .IN3(m4stg_frac[91]), 
        .IN4(n1429), .IN5(n10177), .Q(n9739) );
  AO22X1 U10620 ( .IN1(m4stg_frac[92]), .IN2(n9349), .IN3(m4stg_frac[93]), 
        .IN4(n1445), .Q(n10177) );
  INVX0 U10621 ( .INP(n9696), .ZN(n9614) );
  NAND2X0 U10622 ( .IN1(\fpu_mul_frac_dp/n766 ), .IN2(n908), .QN(n9696) );
  AO221X1 U10623 ( .IN1(n1379), .IN2(n9788), .IN3(n1369), .IN4(n9791), .IN5(
        n10178), .Q(n9825) );
  AO22X1 U10624 ( .IN1(n1367), .IN2(n9787), .IN3(n1361), .IN4(n9858), .Q(
        n10178) );
  AO221X1 U10625 ( .IN1(m4stg_frac[74]), .IN2(n1419), .IN3(m4stg_frac[75]), 
        .IN4(n9347), .IN5(n10179), .Q(n9858) );
  AO22X1 U10626 ( .IN1(m4stg_frac[76]), .IN2(n9349), .IN3(m4stg_frac[77]), 
        .IN4(n1445), .Q(n10179) );
  AO221X1 U10627 ( .IN1(m4stg_frac[78]), .IN2(n1418), .IN3(m4stg_frac[79]), 
        .IN4(n1429), .IN5(n10180), .Q(n9787) );
  AO22X1 U10628 ( .IN1(m4stg_frac[80]), .IN2(n9349), .IN3(m4stg_frac[81]), 
        .IN4(n1445), .Q(n10180) );
  AO221X1 U10629 ( .IN1(m4stg_frac[82]), .IN2(n1419), .IN3(m4stg_frac[83]), 
        .IN4(n9347), .IN5(n10181), .Q(n9791) );
  AO22X1 U10630 ( .IN1(m4stg_frac[84]), .IN2(n9349), .IN3(m4stg_frac[85]), 
        .IN4(n1446), .Q(n10181) );
  AO221X1 U10631 ( .IN1(m4stg_frac[86]), .IN2(n1419), .IN3(m4stg_frac[87]), 
        .IN4(n1429), .IN5(n10182), .Q(n9788) );
  AO22X1 U10632 ( .IN1(m4stg_frac[88]), .IN2(n9349), .IN3(m4stg_frac[89]), 
        .IN4(n1445), .Q(n10182) );
  OA22X1 U10633 ( .IN1(n9993), .IN2(n9654), .IN3(n9992), .IN4(n9655), .Q(
        n10166) );
  NAND2X0 U10634 ( .IN1(n908), .IN2(n1035), .QN(n9655) );
  INVX0 U10635 ( .INP(n10161), .ZN(n9992) );
  AO221X1 U10636 ( .IN1(n1361), .IN2(n10052), .IN3(n1365), .IN4(n10053), .IN5(
        n10183), .Q(n10161) );
  AO22X1 U10637 ( .IN1(n1378), .IN2(n10046), .IN3(n1369), .IN4(n10050), .Q(
        n10183) );
  AO221X1 U10638 ( .IN1(m4stg_frac[50]), .IN2(n1419), .IN3(m4stg_frac[51]), 
        .IN4(n9347), .IN5(n10184), .Q(n10050) );
  AO22X1 U10639 ( .IN1(m4stg_frac[52]), .IN2(n9349), .IN3(m4stg_frac[53]), 
        .IN4(n1446), .Q(n10184) );
  AO221X1 U10640 ( .IN1(m4stg_frac[54]), .IN2(n1419), .IN3(m4stg_frac[55]), 
        .IN4(n1429), .IN5(n10185), .Q(n10046) );
  AO22X1 U10641 ( .IN1(m4stg_frac[56]), .IN2(n9349), .IN3(m4stg_frac[57]), 
        .IN4(n1446), .Q(n10185) );
  AO222X1 U10642 ( .IN1(m4stg_frac[49]), .IN2(n1447), .IN3(n9382), .IN4(n879), 
        .IN5(m4stg_frac[48]), .IN6(n1431), .Q(n10053) );
  MUX21X1 U10643 ( .IN1(m4stg_frac[46]), .IN2(m4stg_frac[47]), .S(
        \fpu_mul_frac_dp/n831 ), .Q(n9382) );
  AO221X1 U10644 ( .IN1(m4stg_frac[42]), .IN2(n1419), .IN3(m4stg_frac[43]), 
        .IN4(n9347), .IN5(n10186), .Q(n10052) );
  AO22X1 U10645 ( .IN1(m4stg_frac[44]), .IN2(n9349), .IN3(m4stg_frac[45]), 
        .IN4(n1446), .Q(n10186) );
  NAND2X0 U10646 ( .IN1(\fpu_mul_frac_dp/n838 ), .IN2(n1035), .QN(n9654) );
  INVX0 U10647 ( .INP(n9823), .ZN(n9993) );
  AO221X1 U10648 ( .IN1(n1378), .IN2(n9856), .IN3(n1370), .IN4(n9885), .IN5(
        n10187), .Q(n9823) );
  AO22X1 U10649 ( .IN1(n1368), .IN2(n9911), .IN3(n1362), .IN4(n10048), .Q(
        n10187) );
  AO221X1 U10650 ( .IN1(m4stg_frac[58]), .IN2(n1419), .IN3(m4stg_frac[59]), 
        .IN4(n9347), .IN5(n10188), .Q(n10048) );
  AO22X1 U10651 ( .IN1(m4stg_frac[60]), .IN2(n9349), .IN3(m4stg_frac[61]), 
        .IN4(n1445), .Q(n10188) );
  AO221X1 U10652 ( .IN1(m4stg_frac[62]), .IN2(n1419), .IN3(m4stg_frac[63]), 
        .IN4(n9347), .IN5(n10189), .Q(n9911) );
  AO22X1 U10653 ( .IN1(m4stg_frac[64]), .IN2(n9349), .IN3(m4stg_frac[65]), 
        .IN4(n1446), .Q(n10189) );
  AO221X1 U10654 ( .IN1(m4stg_frac[66]), .IN2(n1418), .IN3(m4stg_frac[67]), 
        .IN4(n1429), .IN5(n10190), .Q(n9885) );
  AO22X1 U10655 ( .IN1(m4stg_frac[68]), .IN2(n9349), .IN3(m4stg_frac[69]), 
        .IN4(n1445), .Q(n10190) );
  AO221X1 U10656 ( .IN1(m4stg_frac[70]), .IN2(n1411), .IN3(m4stg_frac[71]), 
        .IN4(n1421), .IN5(n10191), .Q(n9856) );
  AO22X1 U10657 ( .IN1(m4stg_frac[72]), .IN2(n1432), .IN3(m4stg_frac[73]), 
        .IN4(n1439), .Q(n10191) );
  NAND2X0 U10658 ( .IN1(\fpu_mul_frac_dp/n834 ), .IN2(\fpu_mul_frac_dp/n831 ), 
        .QN(n9307) );
  INVX0 U10659 ( .INP(n9675), .ZN(n9349) );
  NAND2X0 U10660 ( .IN1(\fpu_mul_frac_dp/n834 ), .IN2(n884), .QN(n9675) );
  INVX0 U10661 ( .INP(n9661), .ZN(n9347) );
  NAND2X0 U10662 ( .IN1(\fpu_mul_frac_dp/n831 ), .IN2(n879), .QN(n9661) );
  NAND2X0 U10663 ( .IN1(\fpu_mul_frac_dp/n833 ), .IN2(\fpu_mul_frac_dp/n765 ), 
        .QN(n9304) );
  NAND2X0 U10664 ( .IN1(m4stg_inc_exp_55), .IN2(n2929), .QN(n9600) );
  NAND2X0 U10665 ( .IN1(fmul_clken_l), .IN2(n1358), .QN(
        \fpu_mul_frac_dp/ckbuf_mul_frac_dp/N1 ) );
  XOR2X1 U10666 ( .IN1(n10192), .IN2(n445), .Q(
        \fpu_mul_exp_dp/m4stg_exp_plus1[9] ) );
  NOR2X0 U10667 ( .IN1(n10193), .IN2(n10194), .QN(
        \fpu_mul_exp_dp/m4stg_exp_plus1[8] ) );
  OA21X1 U10668 ( .IN1(n447), .IN2(n10195), .IN3(n52), .Q(n10194) );
  XOR2X1 U10669 ( .IN1(m4stg_exp[7]), .IN2(n10196), .Q(
        \fpu_mul_exp_dp/m4stg_exp_plus1[7] ) );
  NOR2X0 U10670 ( .IN1(n10196), .IN2(n10197), .QN(
        \fpu_mul_exp_dp/m4stg_exp_plus1[6] ) );
  OA21X1 U10671 ( .IN1(n444), .IN2(n10198), .IN3(n44), .Q(n10197) );
  XOR2X1 U10672 ( .IN1(n10198), .IN2(n444), .Q(
        \fpu_mul_exp_dp/m4stg_exp_plus1[5] ) );
  NOR2X0 U10673 ( .IN1(n10199), .IN2(n10200), .QN(
        \fpu_mul_exp_dp/m4stg_exp_plus1[4] ) );
  OA21X1 U10674 ( .IN1(n446), .IN2(n10201), .IN3(n37), .Q(n10200) );
  XOR2X1 U10675 ( .IN1(m4stg_exp[3]), .IN2(n10202), .Q(
        \fpu_mul_exp_dp/m4stg_exp_plus1[3] ) );
  NOR2X0 U10676 ( .IN1(n10202), .IN2(n10203), .QN(
        \fpu_mul_exp_dp/m4stg_exp_plus1[2] ) );
  OA21X1 U10677 ( .IN1(n442), .IN2(n438), .IN3(n29), .Q(n10203) );
  XOR2X1 U10678 ( .IN1(n442), .IN2(n438), .Q(
        \fpu_mul_exp_dp/m4stg_exp_plus1[1] ) );
  XOR2X1 U10679 ( .IN1(m4stg_exp[11]), .IN2(n10204), .Q(
        \fpu_mul_exp_dp/m4stg_exp_plus1[11] ) );
  NOR2X0 U10680 ( .IN1(n10204), .IN2(n10205), .QN(
        \fpu_mul_exp_dp/m4stg_exp_plus1[10] ) );
  OA21X1 U10681 ( .IN1(n445), .IN2(n10192), .IN3(n60), .Q(n10205) );
  INVX0 U10682 ( .INP(n1630), .ZN(n10204) );
  NAND3X0 U10683 ( .IN1(m4stg_exp[9]), .IN2(m4stg_exp[10]), .IN3(n10193), .QN(
        n1630) );
  INVX0 U10684 ( .INP(n10192), .ZN(n10193) );
  NAND3X0 U10685 ( .IN1(m4stg_exp[7]), .IN2(m4stg_exp[8]), .IN3(n10196), .QN(
        n10192) );
  INVX0 U10686 ( .INP(n10195), .ZN(n10196) );
  NAND3X0 U10687 ( .IN1(m4stg_exp[6]), .IN2(m4stg_exp[5]), .IN3(n10199), .QN(
        n10195) );
  INVX0 U10688 ( .INP(n10198), .ZN(n10199) );
  NAND3X0 U10689 ( .IN1(m4stg_exp[4]), .IN2(m4stg_exp[3]), .IN3(n10202), .QN(
        n10198) );
  INVX0 U10690 ( .INP(n10201), .ZN(n10202) );
  NAND3X0 U10691 ( .IN1(m4stg_exp[0]), .IN2(m4stg_exp[1]), .IN3(m4stg_exp[2]), 
        .QN(n10201) );
  NAND2X0 U10692 ( .IN1(fmul_clken_l_buf1), .IN2(n1360), .QN(
        \fpu_mul_exp_dp/ckbuf_mul_exp_dp/N1 ) );
  AO22X1 U10693 ( .IN1(inq_in1[51]), .IN2(n1601), .IN3(n1403), .IN4(n893), .Q(
        \fpu_mul_ctl/n561 ) );
  AO21X1 U10694 ( .IN1(n1387), .IN2(n894), .IN3(n1633), .Q(\fpu_mul_ctl/n560 )
         );
  AND2X1 U10695 ( .IN1(inq_in1[54]), .IN2(n1593), .Q(n1633) );
  AO22X1 U10696 ( .IN1(inq_in1_53_0_neq_0), .IN2(n1601), .IN3(n1631), .IN4(
        n1336), .Q(\fpu_mul_ctl/n559 ) );
  AO22X1 U10697 ( .IN1(inq_in1_50_0_neq_0), .IN2(n1601), .IN3(n1403), .IN4(
        n1204), .Q(\fpu_mul_ctl/n558 ) );
  AO22X1 U10698 ( .IN1(inq_in1_53_32_neq_0), .IN2(n1601), .IN3(n1631), .IN4(
        n1205), .Q(\fpu_mul_ctl/n557 ) );
  AO22X1 U10699 ( .IN1(inq_in1_exp_eq_0), .IN2(n1601), .IN3(\fpu_mul_ctl/n263 ), .IN4(n1385), .Q(\fpu_mul_ctl/n556 ) );
  AO22X1 U10700 ( .IN1(inq_in1_exp_neq_ffs), .IN2(n1601), .IN3(n1400), .IN4(
        n1037), .Q(\fpu_mul_ctl/n555 ) );
  AO22X1 U10701 ( .IN1(inq_in2[51]), .IN2(n1601), .IN3(n1400), .IN4(n1170), 
        .Q(\fpu_mul_ctl/n554 ) );
  AO21X1 U10702 ( .IN1(n1386), .IN2(n1167), .IN3(n1632), .Q(\fpu_mul_ctl/n553 ) );
  AND2X1 U10703 ( .IN1(inq_in2[54]), .IN2(n1594), .Q(n1632) );
  AO22X1 U10704 ( .IN1(inq_in2_53_0_neq_0), .IN2(n1601), .IN3(n1400), .IN4(
        n1337), .Q(\fpu_mul_ctl/n552 ) );
  AO22X1 U10705 ( .IN1(inq_in2_50_0_neq_0), .IN2(n1601), .IN3(n1400), .IN4(
        n1198), .Q(\fpu_mul_ctl/n551 ) );
  AO22X1 U10706 ( .IN1(inq_in2_53_32_neq_0), .IN2(n1601), .IN3(n1400), .IN4(
        n1197), .Q(\fpu_mul_ctl/n550 ) );
  AO22X1 U10707 ( .IN1(inq_in2_exp_eq_0), .IN2(n1601), .IN3(\fpu_mul_ctl/n264 ), .IN4(n1385), .Q(\fpu_mul_ctl/n549 ) );
  AO22X1 U10708 ( .IN1(inq_in2_exp_neq_ffs), .IN2(n1601), .IN3(n1400), .IN4(
        \fpu_mul_ctl/n253 ), .Q(\fpu_mul_ctl/n548 ) );
  AO22X1 U10709 ( .IN1(n1405), .IN2(n1030), .IN3(n3148), .IN4(n1592), .Q(
        \fpu_mul_ctl/n547 ) );
  AO22X1 U10710 ( .IN1(n1404), .IN2(n1284), .IN3(n3149), .IN4(n1592), .Q(
        \fpu_mul_ctl/n546 ) );
  OAI22X1 U10711 ( .IN1(n1723), .IN2(n1688), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n100 ), .QN(\fpu_mul_ctl/n545 ) );
  NOR2X0 U10712 ( .IN1(n3148), .IN2(n3149), .QN(n1688) );
  AND3X1 U10713 ( .IN1(\fpu_mul_ctl/n264 ), .IN2(\fpu_mul_ctl/n110 ), .IN3(
        \fpu_mul_ctl/n268 ), .Q(n3149) );
  AND3X1 U10714 ( .IN1(\fpu_mul_ctl/n263 ), .IN2(\fpu_mul_ctl/n102 ), .IN3(
        \fpu_mul_ctl/n273 ), .Q(n3148) );
  AO21X1 U10715 ( .IN1(m1stg_sngop), .IN2(n1631), .IN3(n10206), .Q(
        \fpu_mul_ctl/n544 ) );
  AO21X1 U10716 ( .IN1(n1386), .IN2(n1298), .IN3(n10206), .Q(
        \fpu_mul_ctl/n543 ) );
  AO21X1 U10717 ( .IN1(n1386), .IN2(n1056), .IN3(n10206), .Q(
        \fpu_mul_ctl/n542 ) );
  AO21X1 U10718 ( .IN1(n1386), .IN2(n923), .IN3(n10206), .Q(\fpu_mul_ctl/n541 ) );
  AO21X1 U10719 ( .IN1(n1386), .IN2(n910), .IN3(n10206), .Q(\fpu_mul_ctl/n540 ) );
  AND2X1 U10720 ( .IN1(inq_op[0]), .IN2(n1593), .Q(n10206) );
  AO21X1 U10721 ( .IN1(m1stg_dblop), .IN2(n1631), .IN3(n10207), .Q(
        \fpu_mul_ctl/n539 ) );
  AO21X1 U10722 ( .IN1(n1386), .IN2(n1299), .IN3(n10207), .Q(
        \fpu_mul_ctl/n538 ) );
  AO21X1 U10723 ( .IN1(\fpu_mul_ctl/n265 ), .IN2(n1631), .IN3(n10207), .Q(
        \fpu_mul_ctl/n537 ) );
  AO22X1 U10724 ( .IN1(n1405), .IN2(n1344), .IN3(n1593), .IN4(n3143), .Q(
        \fpu_mul_ctl/n536 ) );
  NAND2X0 U10725 ( .IN1(n1887), .IN2(n1881), .QN(n3143) );
  NAND3X0 U10726 ( .IN1(n885), .IN2(n1056), .IN3(n10208), .QN(n1881) );
  NAND2X0 U10727 ( .IN1(\fpu_mul_ctl/n112 ), .IN2(\fpu_mul_ctl/n268 ), .QN(
        n10208) );
  NAND3X0 U10728 ( .IN1(n10209), .IN2(n885), .IN3(\fpu_mul_ctl/n265 ), .QN(
        n1887) );
  NAND2X0 U10729 ( .IN1(\fpu_mul_ctl/n111 ), .IN2(\fpu_mul_ctl/n267 ), .QN(
        n10209) );
  AO22X1 U10730 ( .IN1(n3150), .IN2(n1602), .IN3(n1400), .IN4(n1029), .Q(
        \fpu_mul_ctl/n535 ) );
  AO221X1 U10731 ( .IN1(n1383), .IN2(n1341), .IN3(n3150), .IN4(n1592), .IN5(
        n10210), .Q(\fpu_mul_ctl/n534 ) );
  INVX0 U10732 ( .INP(n3141), .ZN(n3150) );
  NAND2X0 U10733 ( .IN1(\fpu_mul_ctl/n256 ), .IN2(n10211), .QN(n3141) );
  AO22X1 U10734 ( .IN1(n3144), .IN2(n1056), .IN3(n3145), .IN4(
        \fpu_mul_ctl/n265 ), .Q(n10211) );
  NOR2X0 U10735 ( .IN1(n1204), .IN2(n893), .QN(n3145) );
  NOR2X0 U10736 ( .IN1(n1205), .IN2(n894), .QN(n3144) );
  AO21X1 U10737 ( .IN1(n1386), .IN2(n1297), .IN3(n10210), .Q(
        \fpu_mul_ctl/n533 ) );
  AND3X1 U10738 ( .IN1(n3146), .IN2(n885), .IN3(n1608), .Q(n10210) );
  NAND2X0 U10739 ( .IN1(n10212), .IN2(n10213), .QN(n3146) );
  NAND3X0 U10740 ( .IN1(\fpu_mul_ctl/n111 ), .IN2(\fpu_mul_ctl/n267 ), .IN3(
        \fpu_mul_ctl/n265 ), .QN(n10213) );
  NAND3X0 U10741 ( .IN1(\fpu_mul_ctl/n268 ), .IN2(n1056), .IN3(
        \fpu_mul_ctl/n112 ), .QN(n10212) );
  AO21X1 U10742 ( .IN1(n1386), .IN2(n922), .IN3(n10207), .Q(\fpu_mul_ctl/n532 ) );
  AO22X1 U10743 ( .IN1(n1594), .IN2(n3139), .IN3(\fpu_mul_ctl/n730 ), .IN4(
        n1384), .Q(\fpu_mul_ctl/n531 ) );
  INVX0 U10744 ( .INP(n1846), .ZN(n3139) );
  NOR2X0 U10745 ( .IN1(n1854), .IN2(n1853), .QN(n1846) );
  NOR4X0 U10746 ( .IN1(n1037), .IN2(n894), .IN3(\fpu_mul_ctl/n104 ), .IN4(
        \fpu_mul_ctl/n116 ), .QN(n1853) );
  NOR4X0 U10747 ( .IN1(n893), .IN2(n1037), .IN3(\fpu_mul_ctl/n103 ), .IN4(
        \fpu_mul_ctl/n120 ), .QN(n1854) );
  AO22X1 U10748 ( .IN1(n1405), .IN2(n1164), .IN3(n1593), .IN4(n10214), .Q(
        \fpu_mul_ctl/n530 ) );
  NAND2X0 U10749 ( .IN1(n1817), .IN2(n1818), .QN(n10214) );
  NAND4X0 U10750 ( .IN1(\fpu_mul_ctl/n268 ), .IN2(n1197), .IN3(n923), .IN4(
        n885), .QN(n1818) );
  NAND4X0 U10751 ( .IN1(\fpu_mul_ctl/n267 ), .IN2(n1198), .IN3(n922), .IN4(
        n885), .QN(n1817) );
  AO22X1 U10752 ( .IN1(\fpu_mul_ctl/n731 ), .IN2(n1405), .IN3(n10215), .IN4(
        \fpu_mul_ctl/n256 ), .Q(\fpu_mul_ctl/n529 ) );
  NOR2X0 U10753 ( .IN1(n3147), .IN2(n1723), .QN(n10215) );
  OA22X1 U10754 ( .IN1(\fpu_mul_ctl/n120 ), .IN2(\fpu_mul_ctl/n272 ), .IN3(
        \fpu_mul_ctl/n116 ), .IN4(\fpu_mul_ctl/n273 ), .Q(n3147) );
  AO22X1 U10755 ( .IN1(n1594), .IN2(n1847), .IN3(n1400), .IN4(n1328), .Q(
        \fpu_mul_ctl/n528 ) );
  NAND2X0 U10756 ( .IN1(n3082), .IN2(n3153), .QN(n1847) );
  NAND3X0 U10757 ( .IN1(n885), .IN2(n1170), .IN3(n922), .QN(n3153) );
  NAND3X0 U10758 ( .IN1(n885), .IN2(n1167), .IN3(n923), .QN(n3082) );
  AO21X1 U10759 ( .IN1(n1386), .IN2(n886), .IN3(n10207), .Q(\fpu_mul_ctl/n527 ) );
  NOR2X0 U10760 ( .IN1(n10216), .IN2(n1723), .QN(n10207) );
  AO22X1 U10761 ( .IN1(n1594), .IN2(n10216), .IN3(m1stg_dblop_inv), .IN4(n1384), .Q(\fpu_mul_ctl/n526 ) );
  INVX0 U10762 ( .INP(inq_op[1]), .ZN(n10216) );
  AO22X1 U10763 ( .IN1(inq_rnd_mode[1]), .IN2(n1602), .IN3(n1399), .IN4(n1002), 
        .Q(\fpu_mul_ctl/n525 ) );
  AO22X1 U10764 ( .IN1(inq_rnd_mode[0]), .IN2(n1602), .IN3(n1399), .IN4(n1333), 
        .Q(\fpu_mul_ctl/n524 ) );
  AO22X1 U10765 ( .IN1(inq_id[4]), .IN2(n1602), .IN3(n1399), .IN4(n1334), .Q(
        \fpu_mul_ctl/n523 ) );
  AO22X1 U10766 ( .IN1(inq_id[3]), .IN2(n1602), .IN3(n1399), .IN4(n1003), .Q(
        \fpu_mul_ctl/n522 ) );
  AO22X1 U10767 ( .IN1(inq_id[2]), .IN2(n1602), .IN3(n1399), .IN4(n1004), .Q(
        \fpu_mul_ctl/n521 ) );
  AO22X1 U10768 ( .IN1(inq_id[1]), .IN2(n1602), .IN3(n1399), .IN4(n1005), .Q(
        \fpu_mul_ctl/n520 ) );
  AO22X1 U10769 ( .IN1(inq_id[0]), .IN2(n1602), .IN3(n1399), .IN4(n1006), .Q(
        \fpu_mul_ctl/n519 ) );
  AO22X1 U10770 ( .IN1(n1594), .IN2(n1002), .IN3(n1399), .IN4(n1240), .Q(
        \fpu_mul_ctl/n518 ) );
  OAI22X1 U10771 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n135 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n134 ), .QN(\fpu_mul_ctl/n517 ) );
  OAI22X1 U10772 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n142 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n141 ), .QN(\fpu_mul_ctl/n516 ) );
  AO22X1 U10773 ( .IN1(n1594), .IN2(n1003), .IN3(n1399), .IN4(n1241), .Q(
        \fpu_mul_ctl/n515 ) );
  AO22X1 U10774 ( .IN1(n1594), .IN2(n1004), .IN3(n1399), .IN4(n1242), .Q(
        \fpu_mul_ctl/n514 ) );
  AO22X1 U10775 ( .IN1(n1594), .IN2(n1005), .IN3(n1399), .IN4(n1243), .Q(
        \fpu_mul_ctl/n513 ) );
  AO22X1 U10776 ( .IN1(n1594), .IN2(n1006), .IN3(n1399), .IN4(n1244), .Q(
        \fpu_mul_ctl/n512 ) );
  AO22X1 U10777 ( .IN1(n1594), .IN2(n1240), .IN3(n1399), .IN4(n1007), .Q(
        \fpu_mul_ctl/n511 ) );
  OAI22X1 U10778 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n134 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n133 ), .QN(\fpu_mul_ctl/n510 ) );
  OAI22X1 U10779 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n141 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n140 ), .QN(\fpu_mul_ctl/n509 ) );
  AO22X1 U10780 ( .IN1(n1594), .IN2(n1241), .IN3(n1399), .IN4(n1008), .Q(
        \fpu_mul_ctl/n508 ) );
  AO22X1 U10781 ( .IN1(n1594), .IN2(n1242), .IN3(n1398), .IN4(n1009), .Q(
        \fpu_mul_ctl/n507 ) );
  AO22X1 U10782 ( .IN1(n1594), .IN2(n1243), .IN3(n1398), .IN4(n1010), .Q(
        \fpu_mul_ctl/n506 ) );
  AO22X1 U10783 ( .IN1(n1594), .IN2(n1244), .IN3(n1398), .IN4(n1011), .Q(
        \fpu_mul_ctl/n505 ) );
  AO22X1 U10784 ( .IN1(n1595), .IN2(n1007), .IN3(n1398), .IN4(n1245), .Q(
        \fpu_mul_ctl/n504 ) );
  OAI22X1 U10785 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n133 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n132 ), .QN(\fpu_mul_ctl/n503 ) );
  OAI22X1 U10786 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n140 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n139 ), .QN(\fpu_mul_ctl/n502 ) );
  AO22X1 U10787 ( .IN1(n1594), .IN2(n1008), .IN3(n1398), .IN4(n1246), .Q(
        \fpu_mul_ctl/n501 ) );
  AO22X1 U10788 ( .IN1(n1595), .IN2(n1009), .IN3(n1398), .IN4(n1247), .Q(
        \fpu_mul_ctl/n500 ) );
  AO22X1 U10789 ( .IN1(n1594), .IN2(n1010), .IN3(n1398), .IN4(n1248), .Q(
        \fpu_mul_ctl/n499 ) );
  AO22X1 U10790 ( .IN1(n1595), .IN2(n1011), .IN3(n1398), .IN4(n1249), .Q(
        \fpu_mul_ctl/n498 ) );
  AO22X1 U10791 ( .IN1(n1595), .IN2(n1245), .IN3(n1398), .IN4(n1012), .Q(
        \fpu_mul_ctl/n497 ) );
  OAI22X1 U10792 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n132 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n131 ), .QN(\fpu_mul_ctl/n496 ) );
  OAI22X1 U10793 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n139 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n138 ), .QN(\fpu_mul_ctl/n495 ) );
  AO22X1 U10794 ( .IN1(n1595), .IN2(n1246), .IN3(n1398), .IN4(n1013), .Q(
        \fpu_mul_ctl/n494 ) );
  AO22X1 U10795 ( .IN1(n1595), .IN2(n1247), .IN3(n1398), .IN4(n1014), .Q(
        \fpu_mul_ctl/n493 ) );
  AO22X1 U10796 ( .IN1(n1595), .IN2(n1248), .IN3(n1398), .IN4(n1015), .Q(
        \fpu_mul_ctl/n492 ) );
  AO22X1 U10797 ( .IN1(n1595), .IN2(n1249), .IN3(n1398), .IN4(n1016), .Q(
        \fpu_mul_ctl/n491 ) );
  AO22X1 U10798 ( .IN1(n1595), .IN2(n1012), .IN3(n1398), .IN4(n1250), .Q(
        \fpu_mul_ctl/n490 ) );
  OAI22X1 U10799 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n131 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n130 ), .QN(\fpu_mul_ctl/n489 ) );
  OAI22X1 U10800 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n138 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n137 ), .QN(\fpu_mul_ctl/n488 ) );
  AO22X1 U10801 ( .IN1(n1595), .IN2(n1013), .IN3(n1397), .IN4(n1251), .Q(
        \fpu_mul_ctl/n487 ) );
  AO22X1 U10802 ( .IN1(n1595), .IN2(n1014), .IN3(n1397), .IN4(n1252), .Q(
        \fpu_mul_ctl/n486 ) );
  AO22X1 U10803 ( .IN1(n1595), .IN2(n1015), .IN3(n1400), .IN4(n1253), .Q(
        \fpu_mul_ctl/n485 ) );
  AO22X1 U10804 ( .IN1(n1595), .IN2(n1016), .IN3(n1397), .IN4(n1254), .Q(
        \fpu_mul_ctl/n484 ) );
  AO22X1 U10805 ( .IN1(n1595), .IN2(n1250), .IN3(n1397), .IN4(n926), .Q(
        \fpu_mul_ctl/n483 ) );
  OAI22X1 U10806 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n130 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n732 ), .QN(\fpu_mul_ctl/n482 ) );
  OAI22X1 U10807 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n137 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n136 ), .QN(\fpu_mul_ctl/n481 ) );
  AO22X1 U10808 ( .IN1(n1595), .IN2(n1251), .IN3(n1397), .IN4(n931), .Q(
        \fpu_mul_ctl/n480 ) );
  AO22X1 U10809 ( .IN1(n1595), .IN2(n1252), .IN3(n1397), .IN4(n982), .Q(
        \fpu_mul_ctl/n479 ) );
  AO22X1 U10810 ( .IN1(n1596), .IN2(n1253), .IN3(n1397), .IN4(n983), .Q(
        \fpu_mul_ctl/n478 ) );
  AO22X1 U10811 ( .IN1(n1598), .IN2(n1254), .IN3(n1397), .IN4(n984), .Q(
        \fpu_mul_ctl/n477 ) );
  AO22X1 U10812 ( .IN1(m2stg_fsmuld), .IN2(n10217), .IN3(n10218), .IN4(n10219), 
        .Q(\fpu_mul_ctl/n476 ) );
  NOR2X0 U10813 ( .IN1(\fpu_mul_ctl/n257 ), .IN2(n10220), .QN(n10218) );
  AO22X1 U10814 ( .IN1(m2stg_fmuld), .IN2(n10217), .IN3(n10219), .IN4(n1702), 
        .Q(\fpu_mul_ctl/n475 ) );
  AO22X1 U10815 ( .IN1(m2stg_fmuls), .IN2(n10217), .IN3(n10221), .IN4(n10219), 
        .Q(\fpu_mul_ctl/n474 ) );
  NOR2X0 U10816 ( .IN1(n1055), .IN2(n10220), .QN(n10221) );
  AO22X1 U10817 ( .IN1(n10217), .IN2(n1017), .IN3(n10219), .IN4(n3134), .Q(
        \fpu_mul_ctl/n473 ) );
  AO21X1 U10818 ( .IN1(n1680), .IN2(n1055), .IN3(n1702), .Q(n3134) );
  AO22X1 U10819 ( .IN1(n10217), .IN2(n954), .IN3(n10219), .IN4(n2928), .Q(
        \fpu_mul_ctl/n472 ) );
  AO22X1 U10820 ( .IN1(n10217), .IN2(n1255), .IN3(m2stg_fmuld), .IN4(n10219), 
        .Q(\fpu_mul_ctl/n471 ) );
  AO22X1 U10821 ( .IN1(n10217), .IN2(n1018), .IN3(n10219), .IN4(m2stg_fmuls), 
        .Q(\fpu_mul_ctl/n470 ) );
  AO22X1 U10822 ( .IN1(n10217), .IN2(n1256), .IN3(n10219), .IN4(n1017), .Q(
        \fpu_mul_ctl/n469 ) );
  AO22X1 U10823 ( .IN1(n10217), .IN2(n1139), .IN3(n10219), .IN4(n954), .Q(
        \fpu_mul_ctl/n468 ) );
  AO22X1 U10824 ( .IN1(n10217), .IN2(n1019), .IN3(n10219), .IN4(n1255), .Q(
        \fpu_mul_ctl/n467 ) );
  AO22X1 U10825 ( .IN1(n10217), .IN2(n1257), .IN3(n10219), .IN4(n1018), .Q(
        \fpu_mul_ctl/n466 ) );
  AO22X1 U10826 ( .IN1(n10217), .IN2(n1020), .IN3(n10219), .IN4(n1256), .Q(
        \fpu_mul_ctl/n465 ) );
  AO22X1 U10827 ( .IN1(n10217), .IN2(n901), .IN3(n10219), .IN4(n1139), .Q(
        \fpu_mul_ctl/n464 ) );
  AO22X1 U10828 ( .IN1(n10217), .IN2(n1258), .IN3(n10219), .IN4(n1019), .Q(
        \fpu_mul_ctl/n463 ) );
  AO22X1 U10829 ( .IN1(n10217), .IN2(n1021), .IN3(n10219), .IN4(n1257), .Q(
        \fpu_mul_ctl/n462 ) );
  AO22X1 U10830 ( .IN1(n10217), .IN2(n1259), .IN3(n10219), .IN4(n1020), .Q(
        \fpu_mul_ctl/n461 ) );
  AO22X1 U10831 ( .IN1(n10217), .IN2(n883), .IN3(n10219), .IN4(n901), .Q(
        \fpu_mul_ctl/n460 ) );
  AO22X1 U10832 ( .IN1(n10217), .IN2(n966), .IN3(n10219), .IN4(n1258), .Q(
        \fpu_mul_ctl/n459 ) );
  AO22X1 U10833 ( .IN1(m5stg_fmulda), .IN2(n10217), .IN3(n10219), .IN4(n966), 
        .Q(\fpu_mul_ctl/n458 ) );
  AO22X1 U10834 ( .IN1(n10217), .IN2(n1260), .IN3(n10219), .IN4(n1021), .Q(
        \fpu_mul_ctl/n457 ) );
  AO22X1 U10835 ( .IN1(n10217), .IN2(n1022), .IN3(n10219), .IN4(n1259), .Q(
        \fpu_mul_ctl/n456 ) );
  AO22X1 U10836 ( .IN1(n10217), .IN2(n1138), .IN3(n10219), .IN4(n883), .Q(
        \fpu_mul_ctl/n455 ) );
  AO22X1 U10837 ( .IN1(m5stg_fmuld), .IN2(n10217), .IN3(n10219), .IN4(n966), 
        .Q(\fpu_mul_ctl/n454 ) );
  AO22X1 U10838 ( .IN1(m5stg_fmuls), .IN2(n10217), .IN3(n10219), .IN4(n1260), 
        .Q(\fpu_mul_ctl/n453 ) );
  AO22X1 U10839 ( .IN1(n10217), .IN2(n1261), .IN3(n10219), .IN4(n1022), .Q(
        \fpu_mul_ctl/n452 ) );
  AO22X1 U10840 ( .IN1(n10217), .IN2(\fpu_mul_ctl/m5stg_opdec[4] ), .IN3(
        n10219), .IN4(n1138), .Q(\fpu_mul_ctl/n451 ) );
  AO22X1 U10841 ( .IN1(m6stg_fmuls), .IN2(n10217), .IN3(n10219), .IN4(
        m5stg_fmuls), .Q(\fpu_mul_ctl/n450 ) );
  AO22X1 U10842 ( .IN1(m6stg_fmul_dbl_dst), .IN2(n10217), .IN3(n10219), .IN4(
        n1261), .Q(\fpu_mul_ctl/n449 ) );
  AND2X1 U10843 ( .IN1(\fpu_mul_ctl/n735 ), .IN2(\fpu_mul_ctl/n105 ), .Q(
        n10219) );
  AO22X1 U10844 ( .IN1(n1598), .IN2(m6stg_id_in[9]), .IN3(n1397), .IN4(n1262), 
        .Q(\fpu_mul_ctl/n448 ) );
  AO22X1 U10845 ( .IN1(n1798), .IN2(n1262), .IN3(n10222), .IN4(n10223), .Q(
        m6stg_id_in[9]) );
  AO22X1 U10846 ( .IN1(n10224), .IN2(n1216), .IN3(n10225), .IN4(n1592), .Q(
        \fpu_mul_ctl/n447 ) );
  NOR2X0 U10847 ( .IN1(\fpu_mul_ctl/n163 ), .IN2(n1798), .QN(n10225) );
  AO22X1 U10848 ( .IN1(n10224), .IN2(n1217), .IN3(n10226), .IN4(n1592), .Q(
        \fpu_mul_ctl/n446 ) );
  NOR2X0 U10849 ( .IN1(\fpu_mul_ctl/n156 ), .IN2(n1798), .QN(n10226) );
  AO21X1 U10850 ( .IN1(n1798), .IN2(n1360), .IN3(n1383), .Q(n10224) );
  AO22X1 U10851 ( .IN1(n1598), .IN2(m6stg_id_in[2]), .IN3(n1397), .IN4(n1263), 
        .Q(\fpu_mul_ctl/n445 ) );
  AO22X1 U10852 ( .IN1(n1798), .IN2(n1263), .IN3(n10227), .IN4(
        \fpu_mul_ctl/n136 ), .Q(m6stg_id_in[2]) );
  NOR2X0 U10853 ( .IN1(n10228), .IN2(n931), .QN(n10227) );
  AO22X1 U10854 ( .IN1(n1598), .IN2(m6stg_id_in[3]), .IN3(n1397), .IN4(n1264), 
        .Q(\fpu_mul_ctl/n444 ) );
  AO22X1 U10855 ( .IN1(n1798), .IN2(n1264), .IN3(n10229), .IN4(
        \fpu_mul_ctl/n136 ), .Q(m6stg_id_in[3]) );
  NOR2X0 U10856 ( .IN1(n10230), .IN2(n931), .QN(n10229) );
  AO22X1 U10857 ( .IN1(n1598), .IN2(m6stg_id_in[4]), .IN3(n1397), .IN4(n1265), 
        .Q(\fpu_mul_ctl/n443 ) );
  AO22X1 U10858 ( .IN1(n1798), .IN2(n1265), .IN3(n10231), .IN4(
        \fpu_mul_ctl/n136 ), .Q(m6stg_id_in[4]) );
  NOR2X0 U10859 ( .IN1(\fpu_mul_ctl/n143 ), .IN2(n10228), .QN(n10231) );
  AO22X1 U10860 ( .IN1(n1598), .IN2(m6stg_id_in[5]), .IN3(n1397), .IN4(n1266), 
        .Q(\fpu_mul_ctl/n442 ) );
  AO22X1 U10861 ( .IN1(n1798), .IN2(n1266), .IN3(n10232), .IN4(
        \fpu_mul_ctl/n136 ), .Q(m6stg_id_in[5]) );
  NOR2X0 U10862 ( .IN1(\fpu_mul_ctl/n143 ), .IN2(n10230), .QN(n10232) );
  AO22X1 U10863 ( .IN1(n1598), .IN2(m6stg_id_in[6]), .IN3(n1397), .IN4(n1267), 
        .Q(\fpu_mul_ctl/n441 ) );
  AO22X1 U10864 ( .IN1(n1798), .IN2(n1267), .IN3(n10233), .IN4(
        \fpu_mul_ctl/n143 ), .Q(m6stg_id_in[6]) );
  NOR2X0 U10865 ( .IN1(\fpu_mul_ctl/n136 ), .IN2(n10228), .QN(n10233) );
  INVX0 U10866 ( .INP(n10234), .ZN(n10228) );
  AO22X1 U10867 ( .IN1(n1598), .IN2(m6stg_id_in[7]), .IN3(n1396), .IN4(n1268), 
        .Q(\fpu_mul_ctl/n440 ) );
  AO22X1 U10868 ( .IN1(n1798), .IN2(n1268), .IN3(n10235), .IN4(
        \fpu_mul_ctl/n143 ), .Q(m6stg_id_in[7]) );
  NOR2X0 U10869 ( .IN1(\fpu_mul_ctl/n136 ), .IN2(n10230), .QN(n10235) );
  INVX0 U10870 ( .INP(n10223), .ZN(n10230) );
  NOR2X0 U10871 ( .IN1(n1798), .IN2(\fpu_mul_ctl/n260 ), .QN(n10223) );
  AO22X1 U10872 ( .IN1(n1598), .IN2(m6stg_id_in[8]), .IN3(n1396), .IN4(n1269), 
        .Q(\fpu_mul_ctl/n439 ) );
  AO22X1 U10873 ( .IN1(n1798), .IN2(n1269), .IN3(n10222), .IN4(n10234), .Q(
        m6stg_id_in[8]) );
  NOR2X0 U10874 ( .IN1(n982), .IN2(n1798), .QN(n10234) );
  NOR2X0 U10875 ( .IN1(\fpu_mul_ctl/n143 ), .IN2(\fpu_mul_ctl/n136 ), .QN(
        n10222) );
  AO22X1 U10876 ( .IN1(inq_in1[63]), .IN2(n1599), .IN3(n1396), .IN4(n1270), 
        .Q(\fpu_mul_ctl/n438 ) );
  AO22X1 U10877 ( .IN1(inq_in2[63]), .IN2(n1602), .IN3(n1396), .IN4(n1335), 
        .Q(\fpu_mul_ctl/n437 ) );
  AO22X1 U10878 ( .IN1(n1598), .IN2(n1270), .IN3(n1396), .IN4(n980), .Q(
        \fpu_mul_ctl/n436 ) );
  OAI22X1 U10879 ( .IN1(n1723), .IN2(\fpu_mul_ctl/n52 ), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n50 ), .QN(\fpu_mul_ctl/n435 ) );
  AO21X1 U10880 ( .IN1(n1386), .IN2(n1281), .IN3(n1689), .Q(\fpu_mul_ctl/n434 ) );
  AO22X1 U10881 ( .IN1(n10236), .IN2(n10237), .IN3(n1396), .IN4(n1023), .Q(
        \fpu_mul_ctl/n433 ) );
  MUX21X1 U10882 ( .IN1(n10238), .IN2(n10239), .S(n10240), .Q(n10237) );
  AOI221X1 U10883 ( .IN1(\fpu_mul_ctl/n730 ), .IN2(\fpu_mul_ctl/n262 ), .IN3(
        \fpu_mul_ctl/n731 ), .IN4(\fpu_mul_ctl/n107 ), .IN5(\fpu_mul_ctl/n50 ), 
        .QN(n10240) );
  NAND3X0 U10884 ( .IN1(\fpu_mul_ctl/n262 ), .IN2(n980), .IN3(
        \fpu_mul_ctl/n106 ), .QN(n10239) );
  NOR3X0 U10885 ( .IN1(n1164), .IN2(\fpu_mul_ctl/n51 ), .IN3(n10241), .QN(
        n10238) );
  NOR2X0 U10886 ( .IN1(\fpu_mul_ctl/n730 ), .IN2(\fpu_mul_ctl/n106 ), .QN(
        n10241) );
  OA21X1 U10887 ( .IN1(\fpu_mul_ctl/n98 ), .IN2(\fpu_mul_ctl/n100 ), .IN3(
        n1608), .Q(n10236) );
  AO22X1 U10888 ( .IN1(n1631), .IN2(n1289), .IN3(n1593), .IN4(n10242), .Q(
        \fpu_mul_ctl/n432 ) );
  NAND4X0 U10889 ( .IN1(\fpu_mul_ctl/n262 ), .IN2(n10243), .IN3(n10244), .IN4(
        n1332), .QN(n10242) );
  NAND2X0 U10890 ( .IN1(n1030), .IN2(n1297), .QN(n10244) );
  NAND2X0 U10891 ( .IN1(n1284), .IN2(n1029), .QN(n10243) );
  AO22X1 U10892 ( .IN1(n1598), .IN2(n1281), .IN3(n1396), .IN4(n1024), .Q(
        \fpu_mul_ctl/n431 ) );
  AO22X1 U10893 ( .IN1(n1598), .IN2(n1023), .IN3(n1396), .IN4(n1271), .Q(
        \fpu_mul_ctl/n430 ) );
  AO22X1 U10894 ( .IN1(n1598), .IN2(n1289), .IN3(n1396), .IN4(n1025), .Q(
        \fpu_mul_ctl/n429 ) );
  AO22X1 U10895 ( .IN1(n1598), .IN2(n1024), .IN3(n1396), .IN4(n1272), .Q(
        \fpu_mul_ctl/n428 ) );
  AO22X1 U10896 ( .IN1(n1598), .IN2(n1271), .IN3(n1396), .IN4(n1026), .Q(
        \fpu_mul_ctl/n427 ) );
  AO22X1 U10897 ( .IN1(n1598), .IN2(n1025), .IN3(n1396), .IN4(n1273), .Q(
        \fpu_mul_ctl/n426 ) );
  AO22X1 U10898 ( .IN1(n1598), .IN2(n1272), .IN3(n1396), .IN4(n1027), .Q(
        \fpu_mul_ctl/n425 ) );
  AO22X1 U10899 ( .IN1(n1599), .IN2(n1026), .IN3(n1396), .IN4(n1274), .Q(
        \fpu_mul_ctl/n424 ) );
  AO22X1 U10900 ( .IN1(n1599), .IN2(n1273), .IN3(n1395), .IN4(n1028), .Q(
        \fpu_mul_ctl/n423 ) );
  AO22X1 U10901 ( .IN1(n1599), .IN2(n1027), .IN3(n1395), .IN4(n1275), .Q(
        \fpu_mul_ctl/n422 ) );
  AO22X1 U10902 ( .IN1(n1599), .IN2(n1274), .IN3(n1395), .IN4(n988), .Q(
        \fpu_mul_ctl/n421 ) );
  AO22X1 U10903 ( .IN1(n1599), .IN2(n1028), .IN3(n1395), .IN4(n1276), .Q(
        \fpu_mul_ctl/n420 ) );
  AO22X1 U10904 ( .IN1(n1599), .IN2(n1275), .IN3(n1395), .IN4(n981), .Q(
        \fpu_mul_ctl/n419 ) );
  AO22X1 U10905 ( .IN1(n1599), .IN2(n988), .IN3(mul_sign_out), .IN4(n1384), 
        .Q(\fpu_mul_ctl/n418 ) );
  AO22X1 U10906 ( .IN1(n1599), .IN2(n1276), .IN3(mul_exc_out[4]), .IN4(n1384), 
        .Q(\fpu_mul_ctl/n417 ) );
  AO22X1 U10907 ( .IN1(n1631), .IN2(n1346), .IN3(n10245), .IN4(n10246), .Q(
        \fpu_mul_ctl/n416 ) );
  NOR4X0 U10908 ( .IN1(n10247), .IN2(n10248), .IN3(\fpu_mul_ctl/n271 ), .IN4(
        m5stg_exp[12]), .QN(n10246) );
  NAND3X0 U10909 ( .IN1(m5stg_exp[4]), .IN2(m5stg_exp[5]), .IN3(m5stg_exp[3]), 
        .QN(n10247) );
  NOR4X0 U10910 ( .IN1(n10249), .IN2(n1723), .IN3(n10250), .IN4(n1780), .QN(
        n10245) );
  NAND2X0 U10911 ( .IN1(n9163), .IN2(n10251), .QN(n10249) );
  AND3X1 U10912 ( .IN1(n10252), .IN2(n10253), .IN3(n1751), .Q(n9163) );
  XOR2X1 U10913 ( .IN1(\fpu_mul_ctl/n732 ), .IN2(n10254), .Q(n1751) );
  NOR2X0 U10914 ( .IN1(\fpu_mul_ctl/n123 ), .IN2(\fpu_mul_ctl/n733 ), .QN(
        n10254) );
  AO22X1 U10915 ( .IN1(m5stg_fmuls), .IN2(n10255), .IN3(m5stg_fmuld), .IN4(
        n10256), .Q(n10253) );
  AO22X1 U10916 ( .IN1(n10257), .IN2(n926), .IN3(n10258), .IN4(n9744), .Q(
        n10256) );
  NAND3X0 U10917 ( .IN1(n9841), .IN2(n9913), .IN3(n8855), .QN(n10258) );
  INVX0 U10918 ( .INP(n8867), .ZN(n8855) );
  AO21X1 U10919 ( .IN1(n10259), .IN2(n926), .IN3(n9019), .Q(n10255) );
  OR3X1 U10920 ( .IN1(n9032), .IN2(n10259), .IN3(n926), .Q(n10252) );
  OAI21X1 U10921 ( .IN1(n1625), .IN2(\fpu_mul_ctl/n31 ), .IN3(n1778), .QN(
        \fpu_mul_ctl/n415 ) );
  NAND2X0 U10922 ( .IN1(n9164), .IN2(n1608), .QN(n1778) );
  INVX0 U10923 ( .INP(n1773), .ZN(n9164) );
  NAND3X0 U10924 ( .IN1(n10260), .IN2(n981), .IN3(n10261), .QN(n1773) );
  AO222X1 U10925 ( .IN1(m5stg_fmuls), .IN2(n10262), .IN3(n10263), .IN4(n10251), 
        .IN5(m5stg_fmuld), .IN6(m5stg_exp[11]), .Q(n10261) );
  AOI21X1 U10926 ( .IN1(n1219), .IN2(n10264), .IN3(n1793), .QN(n10251) );
  NAND4X0 U10927 ( .IN1(m5stg_fmuld), .IN2(m5stg_exp[10]), .IN3(m5stg_exp[8]), 
        .IN4(m5stg_exp[9]), .QN(n10264) );
  AND2X1 U10928 ( .IN1(m5stg_exp[7]), .IN2(n1791), .Q(n10263) );
  NOR2X0 U10929 ( .IN1(n1788), .IN2(n1790), .QN(n1791) );
  NAND2X0 U10930 ( .IN1(n1786), .IN2(m5stg_exp[4]), .QN(n1788) );
  NOR2X0 U10931 ( .IN1(n1783), .IN2(n1785), .QN(n1786) );
  INVX0 U10932 ( .INP(m5stg_exp[3]), .ZN(n1785) );
  NAND3X0 U10933 ( .IN1(m5stg_exp[1]), .IN2(m5stg_exp[2]), .IN3(m5stg_exp[0]), 
        .QN(n1783) );
  INVX0 U10934 ( .INP(n10265), .ZN(n10262) );
  INVX0 U10935 ( .INP(m5stg_exp[12]), .ZN(n10260) );
  OAI22X1 U10936 ( .IN1(n1625), .IN2(\fpu_mul_ctl/n30 ), .IN3(n1774), .IN4(
        n1723), .QN(\fpu_mul_ctl/n414 ) );
  NAND3X0 U10937 ( .IN1(n9156), .IN2(n9656), .IN3(n9157), .QN(n1774) );
  AND3X1 U10938 ( .IN1(n9151), .IN2(n9145), .IN3(n9146), .Q(n9157) );
  AND3X1 U10939 ( .IN1(n9134), .IN2(n9140), .IN3(n9135), .Q(n9146) );
  AND4X1 U10940 ( .IN1(n9113), .IN2(n9123), .IN3(n10266), .IN4(n9118), .Q(
        n9135) );
  AND2X1 U10941 ( .IN1(n9112), .IN2(n9129), .Q(n10266) );
  AND3X1 U10942 ( .IN1(n9101), .IN2(n9107), .IN3(n9102), .Q(n9113) );
  AND3X1 U10943 ( .IN1(n9090), .IN2(n9096), .IN3(n9091), .Q(n9102) );
  AND3X1 U10944 ( .IN1(n9084), .IN2(n9085), .IN3(n9079), .Q(n9091) );
  AND3X1 U10945 ( .IN1(n9073), .IN2(n9072), .IN3(n9067), .Q(n9079) );
  AND3X1 U10946 ( .IN1(n9060), .IN2(n9061), .IN3(n9055), .Q(n9067) );
  AND3X1 U10947 ( .IN1(n9049), .IN2(n9048), .IN3(n9043), .Q(n9055) );
  OAI22X1 U10948 ( .IN1(n9037), .IN2(n9036), .IN3(n1219), .IN4(n10267), .QN(
        n9043) );
  AND2X1 U10949 ( .IN1(n9036), .IN2(n9037), .Q(n10267) );
  INVX0 U10950 ( .INP(n9032), .ZN(n9036) );
  NAND3X0 U10951 ( .IN1(n9019), .IN2(n9013), .IN3(n9014), .QN(n9037) );
  AND4X1 U10952 ( .IN1(n8992), .IN2(n8997), .IN3(n10268), .IN4(n9002), .Q(
        n9014) );
  AND2X1 U10953 ( .IN1(n9008), .IN2(n8991), .Q(n10268) );
  AND3X1 U10954 ( .IN1(n8986), .IN2(n8980), .IN3(n8981), .Q(n8992) );
  AND3X1 U10955 ( .IN1(n8975), .IN2(n9020), .IN3(n8969), .Q(n8981) );
  AND3X1 U10956 ( .IN1(n9021), .IN2(n8963), .IN3(n8957), .Q(n8969) );
  AND3X1 U10957 ( .IN1(n8951), .IN2(n9022), .IN3(n8945), .Q(n8957) );
  AND3X1 U10958 ( .IN1(n9023), .IN2(n8939), .IN3(n8933), .Q(n8945) );
  AND3X1 U10959 ( .IN1(n8927), .IN2(n9024), .IN3(n8921), .Q(n8933) );
  AND3X1 U10960 ( .IN1(n9025), .IN2(n8915), .IN3(n8909), .Q(n8921) );
  AND3X1 U10961 ( .IN1(n8903), .IN2(n9026), .IN3(n8897), .Q(n8909) );
  AND3X1 U10962 ( .IN1(n8891), .IN2(n9027), .IN3(n8885), .Q(n8897) );
  AND3X1 U10963 ( .IN1(n8879), .IN2(n9028), .IN3(n8873), .Q(n8885) );
  AND4X1 U10964 ( .IN1(m5stg_fmulda), .IN2(n8867), .IN3(n9029), .IN4(n8866), 
        .Q(n8873) );
  AO22X1 U10965 ( .IN1(mul_exc_out[2]), .IN2(n1405), .IN3(n10269), .IN4(n1592), 
        .Q(\fpu_mul_ctl/n413 ) );
  OA21X1 U10966 ( .IN1(m5stg_exp[12]), .IN2(n10270), .IN3(n10271), .Q(n10269)
         );
  NAND4X0 U10967 ( .IN1(n10272), .IN2(n10273), .IN3(n10274), .IN4(n10275), 
        .QN(n10271) );
  NOR4X0 U10968 ( .IN1(n10276), .IN2(n9048), .IN3(n9032), .IN4(n9049), .QN(
        n10275) );
  NAND4X0 U10969 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[33] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[33] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[33] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[33] ), .QN(n9049) );
  NAND4X0 U10970 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[32] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[32] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[32] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[32] ), .QN(n9032) );
  NAND4X0 U10971 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[34] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[34] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[34] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[34] ), .QN(n9048) );
  OR3X1 U10972 ( .IN1(n9060), .IN2(n9061), .IN3(n9073), .Q(n10276) );
  NAND4X0 U10973 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[37] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[37] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[37] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[37] ), .QN(n9073) );
  NAND4X0 U10974 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[35] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[35] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[35] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[35] ), .QN(n9061) );
  NAND4X0 U10975 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[36] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[36] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[36] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[36] ), .QN(n9060) );
  NOR4X0 U10976 ( .IN1(n10277), .IN2(n9084), .IN3(n9072), .IN4(n9085), .QN(
        n10274) );
  NAND4X0 U10977 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[39] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[39] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[39] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[39] ), .QN(n9085) );
  NAND4X0 U10978 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[38] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[38] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[38] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[38] ), .QN(n9072) );
  NAND4X0 U10979 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[40] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[40] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[40] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[40] ), .QN(n9084) );
  OR3X1 U10980 ( .IN1(n9096), .IN2(n9090), .IN3(n9101), .Q(n10277) );
  NAND4X0 U10981 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[43] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[43] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[43] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[43] ), .QN(n9101) );
  NAND4X0 U10982 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[41] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[41] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[41] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[41] ), .QN(n9090) );
  NAND4X0 U10983 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[42] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[42] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[42] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[42] ), .QN(n9096) );
  NOR4X0 U10984 ( .IN1(n10278), .IN2(n9118), .IN3(n9107), .IN4(n9112), .QN(
        n10273) );
  NAND4X0 U10985 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[45] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[45] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[45] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[45] ), .QN(n9112) );
  NAND4X0 U10986 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[44] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[44] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[44] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[44] ), .QN(n9107) );
  NAND4X0 U10987 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[46] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[46] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[46] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[46] ), .QN(n9118) );
  OR3X1 U10988 ( .IN1(n9129), .IN2(n9123), .IN3(n9134), .Q(n10278) );
  NAND4X0 U10989 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[49] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[49] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[49] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[49] ), .QN(n9134) );
  NAND4X0 U10990 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[47] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[47] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[47] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[47] ), .QN(n9123) );
  NAND4X0 U10991 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[48] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[48] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[48] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[48] ), .QN(n9129) );
  NOR4X0 U10992 ( .IN1(n10279), .IN2(n9151), .IN3(n9140), .IN4(n9145), .QN(
        n10272) );
  NAND4X0 U10993 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[51] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[51] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[51] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[51] ), .QN(n9145) );
  NAND4X0 U10994 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[50] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[50] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[50] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[50] ), .QN(n9140) );
  NAND4X0 U10995 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[52] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[52] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[52] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[52] ), .QN(n9151) );
  OR3X1 U10996 ( .IN1(n9656), .IN2(n9156), .IN3(n10280), .Q(n10279) );
  NAND4X0 U10997 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[53] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[53] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[53] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[53] ), .QN(n9156) );
  NAND4X0 U10998 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre3[54] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre2[54] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[54] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre4[54] ), .QN(n9656) );
  NOR4X0 U10999 ( .IN1(n10281), .IN2(n10282), .IN3(m5stg_exp[4]), .IN4(
        m5stg_exp[3]), .QN(n10270) );
  NAND2X0 U11000 ( .IN1(n10283), .IN2(n30), .QN(m5stg_exp[3]) );
  MUX21X1 U11001 ( .IN1(n32), .IN2(n162), .S(n10284), .Q(n10283) );
  NAND2X0 U11002 ( .IN1(n10285), .IN2(n34), .QN(m5stg_exp[4]) );
  MUX21X1 U11003 ( .IN1(n36), .IN2(n160), .S(n10284), .Q(n10285) );
  NAND3X0 U11004 ( .IN1(n1793), .IN2(n10248), .IN3(n1790), .QN(n10282) );
  INVX0 U11005 ( .INP(m5stg_exp[5]), .ZN(n1790) );
  NAND2X0 U11006 ( .IN1(n10286), .IN2(n38), .QN(m5stg_exp[5]) );
  MUX21X1 U11007 ( .IN1(n40), .IN2(n158), .S(n10284), .Q(n10286) );
  INVX0 U11008 ( .INP(m5stg_exp[7]), .ZN(n10248) );
  NAND2X0 U11009 ( .IN1(n10287), .IN2(n45), .QN(m5stg_exp[7]) );
  MUX21X1 U11010 ( .IN1(n47), .IN2(n180), .S(n10284), .Q(n10287) );
  INVX0 U11011 ( .INP(m5stg_exp[6]), .ZN(n1793) );
  NAND2X0 U11012 ( .IN1(n10288), .IN2(n12), .QN(m5stg_exp[6]) );
  MUX21X1 U11013 ( .IN1(n43), .IN2(n156), .S(n10284), .Q(n10288) );
  NAND4X0 U11014 ( .IN1(n10265), .IN2(n1756), .IN3(n1780), .IN4(n10250), .QN(
        n10281) );
  INVX0 U11015 ( .INP(m5stg_exp[2]), .ZN(n10250) );
  NAND2X0 U11016 ( .IN1(n10289), .IN2(n26), .QN(m5stg_exp[2]) );
  MUX21X1 U11017 ( .IN1(n28), .IN2(n164), .S(n10284), .Q(n10289) );
  INVX0 U11018 ( .INP(m5stg_exp[1]), .ZN(n1780) );
  NAND2X0 U11019 ( .IN1(n10290), .IN2(n22), .QN(m5stg_exp[1]) );
  MUX21X1 U11020 ( .IN1(n24), .IN2(n166), .S(n10284), .Q(n10290) );
  INVX0 U11021 ( .INP(m5stg_exp[0]), .ZN(n1756) );
  NAND2X0 U11022 ( .IN1(n10291), .IN2(n18), .QN(m5stg_exp[0]) );
  MUX21X1 U11023 ( .IN1(n20), .IN2(n168), .S(n10284), .Q(n10291) );
  NOR4X0 U11024 ( .IN1(m5stg_exp[10]), .IN2(m5stg_exp[11]), .IN3(m5stg_exp[8]), 
        .IN4(m5stg_exp[9]), .QN(n10265) );
  NAND2X0 U11025 ( .IN1(n10292), .IN2(n53), .QN(m5stg_exp[9]) );
  MUX21X1 U11026 ( .IN1(n55), .IN2(n176), .S(n10284), .Q(n10292) );
  NAND2X0 U11027 ( .IN1(n10293), .IN2(n49), .QN(m5stg_exp[8]) );
  MUX21X1 U11028 ( .IN1(n51), .IN2(n178), .S(n10284), .Q(n10293) );
  NAND2X0 U11029 ( .IN1(n10294), .IN2(n61), .QN(m5stg_exp[11]) );
  MUX21X1 U11030 ( .IN1(n63), .IN2(n172), .S(n10284), .Q(n10294) );
  NAND2X0 U11031 ( .IN1(n10295), .IN2(n57), .QN(m5stg_exp[10]) );
  MUX21X1 U11032 ( .IN1(n59), .IN2(n174), .S(n10284), .Q(n10295) );
  AO21X1 U11033 ( .IN1(n10284), .IN2(\fpu_mul_exp_dp/m5stg_exp_pre1[12] ), 
        .IN3(n877), .Q(m5stg_exp[12]) );
  AO221X1 U11034 ( .IN1(\fpu_mul_exp_dp/m5stg_shl_54 ), .IN2(
        \fpu_mul_exp_dp/m5stg_inc_exp_54 ), .IN3(
        \fpu_mul_exp_dp/m5stg_inc_exp_55 ), .IN4(\fpu_mul_exp_dp/m5stg_shl_55 ), .IN5(\fpu_mul_exp_dp/m5stg_inc_exp_105 ), .Q(n10284) );
  AO22X1 U11035 ( .IN1(n1404), .IN2(n1345), .IN3(n1593), .IN4(n10296), .Q(
        \fpu_mul_ctl/n412 ) );
  AO22X1 U11036 ( .IN1(m5stg_fmuls), .IN2(n10280), .IN3(m5stg_fmuld), .IN4(
        n10257), .Q(n10296) );
  OR2X1 U11037 ( .IN1(n10259), .IN2(n9019), .Q(n10280) );
  NAND4X0 U11038 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre4[31] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre3[31] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre2[31] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre1[31] ), .QN(n9019) );
  NAND4X0 U11039 ( .IN1(n10297), .IN2(n10298), .IN3(n10299), .IN4(n10300), 
        .QN(n10259) );
  NOR2X0 U11040 ( .IN1(n10301), .IN2(n10302), .QN(n10300) );
  NAND4X0 U11041 ( .IN1(n8926), .IN2(n8932), .IN3(n8938), .IN4(n8944), .QN(
        n10302) );
  INVX0 U11042 ( .INP(n8951), .ZN(n8944) );
  NAND4X0 U11043 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[18] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[18] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[18] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[18] ), .QN(n8951) );
  INVX0 U11044 ( .INP(n9023), .ZN(n8938) );
  NAND4X0 U11045 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[17] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[17] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[17] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[17] ), .QN(n9023) );
  INVX0 U11046 ( .INP(n8939), .ZN(n8932) );
  NAND4X0 U11047 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[16] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[16] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[16] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[16] ), .QN(n8939) );
  INVX0 U11048 ( .INP(n9024), .ZN(n8926) );
  NAND4X0 U11049 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[15] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[15] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[15] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[15] ), .QN(n9024) );
  OR4X1 U11050 ( .IN1(n9025), .IN2(n8927), .IN3(n10257), .IN4(n8867), .Q(
        n10301) );
  NAND4X0 U11051 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[3] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[3] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[3] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[3] ), .QN(n8867) );
  NAND3X0 U11052 ( .IN1(n9841), .IN2(n9913), .IN3(n10303), .QN(n10257) );
  INVX0 U11053 ( .INP(n9744), .ZN(n10303) );
  NAND4X0 U11054 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[2] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[2] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[2] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[2] ), .QN(n9744) );
  AND3X1 U11055 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre4[0] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre3[0] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre1[0] ), .Q(n9913) );
  AND4X1 U11056 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[1] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[1] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[1] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[1] ), .Q(n9841) );
  NAND4X0 U11057 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[14] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[14] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[14] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[14] ), .QN(n8927) );
  NAND4X0 U11058 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[13] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[13] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[13] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[13] ), .QN(n9025) );
  NOR4X0 U11059 ( .IN1(n10304), .IN2(n9020), .IN3(n8986), .IN4(n8980), .QN(
        n10299) );
  NAND4X0 U11060 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[24] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[24] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[24] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[24] ), .QN(n8980) );
  NAND4X0 U11061 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[25] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[25] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[25] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[25] ), .QN(n8986) );
  NAND4X0 U11062 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[23] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[23] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[23] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[23] ), .QN(n9020) );
  NAND4X0 U11063 ( .IN1(n8950), .IN2(n8956), .IN3(n8962), .IN4(n8968), .QN(
        n10304) );
  INVX0 U11064 ( .INP(n8975), .ZN(n8968) );
  NAND4X0 U11065 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[22] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[22] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[22] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[22] ), .QN(n8975) );
  INVX0 U11066 ( .INP(n9021), .ZN(n8962) );
  NAND4X0 U11067 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[21] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[21] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[21] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[21] ), .QN(n9021) );
  INVX0 U11068 ( .INP(n8963), .ZN(n8956) );
  NAND4X0 U11069 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[20] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[20] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[20] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[20] ), .QN(n8963) );
  INVX0 U11070 ( .INP(n9022), .ZN(n8950) );
  NAND4X0 U11071 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[19] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[19] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[19] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[19] ), .QN(n9022) );
  NOR4X0 U11072 ( .IN1(n10305), .IN2(n9008), .IN3(n8866), .IN4(n9013), .QN(
        n10298) );
  NAND4X0 U11073 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[30] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[30] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[30] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[30] ), .QN(n9013) );
  NAND4X0 U11074 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[5] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[5] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[5] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[5] ), .QN(n8866) );
  NAND4X0 U11075 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[29] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[29] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[29] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[29] ), .QN(n9008) );
  OR4X1 U11076 ( .IN1(n8991), .IN2(n9002), .IN3(n8997), .IN4(n9029), .Q(n10305) );
  NAND4X0 U11077 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[4] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[4] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[4] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[4] ), .QN(n9029) );
  NAND4X0 U11078 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[27] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[27] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[27] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[27] ), .QN(n8997) );
  NAND4X0 U11079 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[28] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[28] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[28] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[28] ), .QN(n9002) );
  NAND4X0 U11080 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[26] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[26] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[26] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[26] ), .QN(n8991) );
  NOR4X0 U11081 ( .IN1(n10306), .IN2(n9027), .IN3(n9028), .IN4(n8891), .QN(
        n10297) );
  NAND4X0 U11082 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[8] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[8] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[8] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[8] ), .QN(n8891) );
  NAND4X0 U11083 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[7] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[7] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[7] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[7] ), .QN(n9028) );
  NAND4X0 U11084 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[9] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[9] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[9] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[9] ), .QN(n9027) );
  NAND4X0 U11085 ( .IN1(n8872), .IN2(n8908), .IN3(n8902), .IN4(n8896), .QN(
        n10306) );
  INVX0 U11086 ( .INP(n8903), .ZN(n8896) );
  NAND4X0 U11087 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[10] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[10] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[10] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[10] ), .QN(n8903) );
  INVX0 U11088 ( .INP(n9026), .ZN(n8902) );
  NAND4X0 U11089 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[11] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[11] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[11] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[11] ), .QN(n9026) );
  INVX0 U11090 ( .INP(n8915), .ZN(n8908) );
  NAND4X0 U11091 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[12] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[12] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[12] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[12] ), .QN(n8915) );
  INVX0 U11092 ( .INP(n8879), .ZN(n8872) );
  NAND4X0 U11093 ( .IN1(\fpu_mul_frac_dp/m5stg_frac_pre1[6] ), .IN2(
        \fpu_mul_frac_dp/m5stg_frac_pre4[6] ), .IN3(
        \fpu_mul_frac_dp/m5stg_frac_pre3[6] ), .IN4(
        \fpu_mul_frac_dp/m5stg_frac_pre2[6] ), .QN(n8879) );
  AO22X1 U11094 ( .IN1(n10307), .IN2(n10308), .IN3(n1395), .IN4(n974), .Q(
        \fpu_mul_ctl/n411 ) );
  AO221X1 U11095 ( .IN1(n10309), .IN2(n10310), .IN3(n10311), .IN4(n10312), 
        .IN5(n10313), .Q(n10308) );
  MUX21X1 U11096 ( .IN1(n10314), .IN2(n10315), .S(n10316), .Q(n10313) );
  NOR2X0 U11097 ( .IN1(n10317), .IN2(n10318), .QN(n10315) );
  OA21X1 U11098 ( .IN1(n10319), .IN2(n10320), .IN3(n10321), .Q(n10317) );
  INVX0 U11099 ( .INP(n10322), .ZN(n10320) );
  OA21X1 U11100 ( .IN1(n10323), .IN2(n10324), .IN3(n10325), .Q(n10319) );
  INVX0 U11101 ( .INP(n10326), .ZN(n10324) );
  OA21X1 U11102 ( .IN1(n10327), .IN2(n10328), .IN3(n10329), .Q(n10323) );
  INVX0 U11103 ( .INP(n10330), .ZN(n10328) );
  OA21X1 U11104 ( .IN1(n10331), .IN2(n10332), .IN3(n10333), .Q(n10314) );
  INVX0 U11105 ( .INP(n10334), .ZN(n10332) );
  NOR2X0 U11106 ( .IN1(n10335), .IN2(n10336), .QN(n10331) );
  INVX0 U11107 ( .INP(n10337), .ZN(n10336) );
  OA221X1 U11108 ( .IN1(n10338), .IN2(n10339), .IN3(n10340), .IN4(n10339), 
        .IN5(n10341), .Q(n10335) );
  MUX21X1 U11109 ( .IN1(n10342), .IN2(n10343), .S(n10344), .Q(n10311) );
  NAND2X0 U11110 ( .IN1(m1stg_dblop), .IN2(n10345), .QN(n10343) );
  AO21X1 U11111 ( .IN1(\fpu_mul_frac_dp/n792 ), .IN2(n956), .IN3(n1180), .Q(
        n10345) );
  NOR2X0 U11112 ( .IN1(n10346), .IN2(n10347), .QN(n10342) );
  OA221X1 U11113 ( .IN1(n10348), .IN2(n10349), .IN3(n10350), .IN4(n1121), 
        .IN5(n10351), .Q(n10347) );
  OA21X1 U11114 ( .IN1(\fpu_mul_frac_dp/n781 ), .IN2(n952), .IN3(
        \fpu_mul_frac_dp/n802 ), .Q(n10350) );
  NOR2X0 U11115 ( .IN1(\fpu_mul_frac_dp/n756 ), .IN2(n943), .QN(n10348) );
  OA21X1 U11116 ( .IN1(n10352), .IN2(n882), .IN3(n10353), .Q(n10346) );
  OA21X1 U11117 ( .IN1(n10354), .IN2(n899), .IN3(\fpu_mul_frac_dp/n805 ), .Q(
        n10352) );
  OA21X1 U11118 ( .IN1(\fpu_mul_frac_dp/n795 ), .IN2(n1202), .IN3(
        \fpu_mul_frac_dp/n778 ), .Q(n10354) );
  OA22X1 U11119 ( .IN1(n10355), .IN2(n10356), .IN3(n10357), .IN4(n10358), .Q(
        n10309) );
  MUX21X1 U11120 ( .IN1(n10359), .IN2(n10360), .S(n10361), .Q(n10358) );
  OA21X1 U11121 ( .IN1(n10362), .IN2(\fpu_mul_frac_dp/n763 ), .IN3(
        \fpu_mul_frac_dp/n786 ), .Q(n10360) );
  OA21X1 U11122 ( .IN1(n10363), .IN2(\fpu_mul_frac_dp/n796 ), .IN3(
        \fpu_mul_frac_dp/n785 ), .Q(n10359) );
  OA21X1 U11123 ( .IN1(n10364), .IN2(n10365), .IN3(n10366), .Q(n10356) );
  INVX0 U11124 ( .INP(n10367), .ZN(n10365) );
  NOR2X0 U11125 ( .IN1(n10368), .IN2(n10369), .QN(n10364) );
  OA21X1 U11126 ( .IN1(\fpu_mul_frac_dp/n357 ), .IN2(n1031), .IN3(
        \fpu_mul_frac_dp/n354 ), .Q(n10368) );
  OA21X1 U11127 ( .IN1(n10370), .IN2(n10371), .IN3(n10372), .Q(n10355) );
  NAND4X0 U11128 ( .IN1(n10373), .IN2(n10374), .IN3(n10375), .IN4(n10376), 
        .QN(\fpu_mul_ctl/n410 ) );
  OA222X1 U11129 ( .IN1(\fpu_mul_ctl/n26 ), .IN2(n1625), .IN3(n10377), .IN4(
        n10378), .IN5(n10379), .IN6(n10380), .Q(n10376) );
  OA22X1 U11130 ( .IN1(n10381), .IN2(n10382), .IN3(n10383), .IN4(n10384), .Q(
        n10379) );
  AO21X1 U11131 ( .IN1(n10385), .IN2(n10386), .IN3(n10371), .Q(n10384) );
  INVX0 U11132 ( .INP(n10387), .ZN(n10371) );
  AO21X1 U11133 ( .IN1(n10362), .IN2(n10388), .IN3(n10363), .Q(n10386) );
  OA22X1 U11134 ( .IN1(n1171), .IN2(n10389), .IN3(n10349), .IN4(n943), .Q(
        n10377) );
  OR2X1 U11135 ( .IN1(n1121), .IN2(n10390), .Q(n10389) );
  OA21X1 U11136 ( .IN1(n10391), .IN2(n10392), .IN3(n10393), .Q(n10375) );
  NAND4X0 U11137 ( .IN1(n10394), .IN2(\fpu_mul_frac_dp/n805 ), .IN3(
        \fpu_mul_frac_dp/n759 ), .IN4(n10395), .QN(n10393) );
  NAND3X0 U11138 ( .IN1(\fpu_mul_frac_dp/n751 ), .IN2(n10396), .IN3(
        \fpu_mul_frac_dp/n778 ), .QN(n10395) );
  NAND3X0 U11139 ( .IN1(\fpu_mul_frac_dp/n795 ), .IN2(n10397), .IN3(
        \fpu_mul_frac_dp/n807 ), .QN(n10396) );
  AO21X1 U11140 ( .IN1(n10398), .IN2(n10399), .IN3(n10400), .Q(n10392) );
  NAND3X0 U11141 ( .IN1(n10338), .IN2(n10401), .IN3(n10402), .QN(n10399) );
  NAND4X0 U11142 ( .IN1(n10403), .IN2(\fpu_mul_frac_dp/n764 ), .IN3(n10404), 
        .IN4(\fpu_mul_frac_dp/n792 ), .QN(n10374) );
  OA21X1 U11143 ( .IN1(n1208), .IN2(n956), .IN3(m1stg_dblop), .Q(n10404) );
  INVX0 U11144 ( .INP(n10405), .ZN(n10403) );
  NAND4X0 U11145 ( .IN1(n10406), .IN2(n10325), .IN3(n10322), .IN4(n10407), 
        .QN(n10373) );
  AO21X1 U11146 ( .IN1(n10330), .IN2(n10327), .IN3(n10408), .Q(n10407) );
  NAND4X0 U11147 ( .IN1(n10409), .IN2(n10410), .IN3(n10411), .IN4(n10412), 
        .QN(\fpu_mul_ctl/n409 ) );
  NAND4X0 U11148 ( .IN1(n10413), .IN2(\fpu_mul_frac_dp/n802 ), .IN3(
        \fpu_mul_frac_dp/n760 ), .IN4(n10390), .QN(n10412) );
  NAND3X0 U11149 ( .IN1(n10414), .IN2(n10415), .IN3(n10307), .QN(n10411) );
  NAND3X0 U11150 ( .IN1(n10416), .IN2(n10417), .IN3(n10418), .QN(n10415) );
  NAND3X0 U11151 ( .IN1(n10398), .IN2(n10419), .IN3(n10420), .QN(n10418) );
  NAND4X0 U11152 ( .IN1(n10402), .IN2(n10421), .IN3(n10338), .IN4(n10422), 
        .QN(n10419) );
  NAND4X0 U11153 ( .IN1(n10325), .IN2(n10322), .IN3(n10423), .IN4(n10424), 
        .QN(n10422) );
  INVX0 U11154 ( .INP(n10401), .ZN(n10421) );
  NAND4X0 U11155 ( .IN1(n10316), .IN2(n10318), .IN3(n10425), .IN4(n10426), 
        .QN(n10416) );
  NOR2X0 U11156 ( .IN1(n10427), .IN2(n10428), .QN(n10425) );
  AO21X1 U11157 ( .IN1(n10429), .IN2(n10397), .IN3(n10430), .Q(n10414) );
  AO21X1 U11158 ( .IN1(m1stg_dblop), .IN2(n10431), .IN3(n10405), .Q(n10410) );
  NAND4X0 U11159 ( .IN1(\fpu_mul_frac_dp/n827 ), .IN2(\fpu_mul_frac_dp/n382 ), 
        .IN3(\fpu_mul_frac_dp/n764 ), .IN4(\fpu_mul_frac_dp/n792 ), .QN(n10431) );
  OR2X1 U11160 ( .IN1(n1625), .IN2(\fpu_mul_ctl/n25 ), .Q(n10409) );
  OAI221X1 U11161 ( .IN1(n10380), .IN2(n10357), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n24 ), .IN5(n10432), .QN(\fpu_mul_ctl/n408 ) );
  NOR2X0 U11162 ( .IN1(n10413), .IN2(n10406), .QN(n10432) );
  AND3X1 U11163 ( .IN1(n10316), .IN2(n10424), .IN3(n10307), .Q(n10406) );
  INVX0 U11164 ( .INP(n10378), .ZN(n10413) );
  NAND2X0 U11165 ( .IN1(n10394), .IN2(n10351), .QN(n10378) );
  NOR2X0 U11166 ( .IN1(n10433), .IN2(n10344), .QN(n10394) );
  NAND3X0 U11167 ( .IN1(n10405), .IN2(n10380), .IN3(n10434), .QN(
        \fpu_mul_ctl/n407 ) );
  OR2X1 U11168 ( .IN1(n1625), .IN2(\fpu_mul_ctl/n23 ), .Q(n10434) );
  NAND2X0 U11169 ( .IN1(n10307), .IN2(n10310), .QN(n10380) );
  AND3X1 U11170 ( .IN1(n10318), .IN2(n10430), .IN3(n10316), .Q(n10310) );
  INVX0 U11171 ( .INP(n10312), .ZN(n10430) );
  NAND2X0 U11172 ( .IN1(n10435), .IN2(n10344), .QN(n10405) );
  NAND2X0 U11173 ( .IN1(m1stg_dblop), .IN2(n10436), .QN(n10344) );
  NAND4X0 U11174 ( .IN1(\fpu_mul_frac_dp/n806 ), .IN2(\fpu_mul_frac_dp/n787 ), 
        .IN3(n10437), .IN4(\fpu_mul_frac_dp/n756 ), .QN(n10436) );
  NOR2X0 U11175 ( .IN1(n10349), .IN2(n10397), .QN(n10437) );
  INVX0 U11176 ( .INP(n10351), .ZN(n10397) );
  NOR2X0 U11177 ( .IN1(n10353), .IN2(\fpu_mul_frac_dp/n836 ), .QN(n10351) );
  NAND4X0 U11178 ( .IN1(\fpu_mul_frac_dp/n821 ), .IN2(\fpu_mul_frac_dp/n807 ), 
        .IN3(\fpu_mul_frac_dp/n795 ), .IN4(n10429), .QN(n10353) );
  NOR4X0 U11179 ( .IN1(n960), .IN2(n1159), .IN3(n882), .IN4(n899), .QN(n10429)
         );
  NAND4X0 U11180 ( .IN1(\fpu_mul_frac_dp/n828 ), .IN2(\fpu_mul_frac_dp/n802 ), 
        .IN3(\fpu_mul_frac_dp/n760 ), .IN4(n10390), .QN(n10349) );
  NOR2X0 U11181 ( .IN1(n1186), .IN2(n952), .QN(n10390) );
  INVX0 U11182 ( .INP(n10433), .ZN(n10435) );
  OAI21X1 U11183 ( .IN1(n1625), .IN2(\fpu_mul_ctl/n22 ), .IN3(n10433), .QN(
        \fpu_mul_ctl/n406 ) );
  NAND2X0 U11184 ( .IN1(n10307), .IN2(n10312), .QN(n10433) );
  NOR3X0 U11185 ( .IN1(n10438), .IN2(n10362), .IN3(n10417), .QN(n10312) );
  NAND4X0 U11186 ( .IN1(n10316), .IN2(n10318), .IN3(n10361), .IN4(n10427), 
        .QN(n10417) );
  INVX0 U11187 ( .INP(n10357), .ZN(n10427) );
  NAND3X0 U11188 ( .IN1(n10387), .IN2(n10385), .IN3(n10372), .QN(n10357) );
  INVX0 U11189 ( .INP(n10383), .ZN(n10372) );
  NAND3X0 U11190 ( .IN1(n10426), .IN2(n10381), .IN3(n10439), .QN(n10383) );
  OA22X1 U11191 ( .IN1(\fpu_mul_frac_dp/n358 ), .IN2(n1031), .IN3(
        \fpu_mul_frac_dp/n355 ), .IN4(n1032), .Q(n10439) );
  INVX0 U11192 ( .INP(n10428), .ZN(n10381) );
  AO221X1 U11193 ( .IN1(m1stg_dblop_inv), .IN2(n1182), .IN3(m1stg_dblop), 
        .IN4(n967), .IN5(n10369), .Q(n10428) );
  AO22X1 U11194 ( .IN1(m1stg_dblop_inv), .IN2(n947), .IN3(m1stg_dblop), .IN4(
        n1183), .Q(n10369) );
  INVX0 U11195 ( .INP(n10382), .ZN(n10426) );
  NAND2X0 U11196 ( .IN1(n10367), .IN2(n10366), .QN(n10382) );
  OA22X1 U11197 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n351 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n354 ), .Q(n10366) );
  OA22X1 U11198 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n352 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n355 ), .Q(n10367) );
  OA21X1 U11199 ( .IN1(n1207), .IN2(n1031), .IN3(n10370), .Q(n10385) );
  OA22X1 U11200 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n357 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n360 ), .Q(n10370) );
  OA22X1 U11201 ( .IN1(n1031), .IN2(\fpu_mul_frac_dp/n359 ), .IN3(n1032), 
        .IN4(\fpu_mul_frac_dp/n356 ), .Q(n10387) );
  OA21X1 U11202 ( .IN1(n1031), .IN2(n10388), .IN3(n10440), .Q(n10361) );
  INVX0 U11203 ( .INP(n10363), .ZN(n10440) );
  OA21X1 U11204 ( .IN1(n1220), .IN2(n986), .IN3(m1stg_dblop), .Q(n10363) );
  NOR2X0 U11205 ( .IN1(n1201), .IN2(n978), .QN(n10388) );
  INVX0 U11206 ( .INP(n10424), .ZN(n10318) );
  AO221X1 U11207 ( .IN1(m1stg_dblop_inv), .IN2(n1187), .IN3(m1stg_dblop), 
        .IN4(n947), .IN5(n10321), .Q(n10424) );
  NAND4X0 U11208 ( .IN1(n10322), .IN2(n10330), .IN3(n10325), .IN4(n10441), 
        .QN(n10321) );
  OA221X1 U11209 ( .IN1(\fpu_mul_frac_dp/n352 ), .IN2(n1031), .IN3(
        \fpu_mul_frac_dp/n349 ), .IN4(n1032), .IN5(n10442), .Q(n10441) );
  AND2X1 U11210 ( .IN1(n10423), .IN2(n10327), .Q(n10442) );
  OA22X1 U11211 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n348 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n351 ), .Q(n10327) );
  INVX0 U11212 ( .INP(n10408), .ZN(n10423) );
  NAND2X0 U11213 ( .IN1(n10329), .IN2(n10326), .QN(n10408) );
  OA22X1 U11214 ( .IN1(n1031), .IN2(\fpu_mul_frac_dp/n348 ), .IN3(n1032), 
        .IN4(\fpu_mul_frac_dp/n345 ), .Q(n10326) );
  OA22X1 U11215 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n346 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n349 ), .Q(n10329) );
  OA22X1 U11216 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n344 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n347 ), .Q(n10325) );
  OA22X1 U11217 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n347 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n350 ), .Q(n10330) );
  OA22X1 U11218 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n343 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n346 ), .Q(n10322) );
  AND4X1 U11219 ( .IN1(n10420), .IN2(n10398), .IN3(n10338), .IN4(n10443), .Q(
        n10316) );
  NOR2X0 U11220 ( .IN1(n10401), .IN2(n10339), .QN(n10443) );
  INVX0 U11221 ( .INP(n10402), .ZN(n10339) );
  OA22X1 U11222 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n339 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n342 ), .Q(n10402) );
  AO221X1 U11223 ( .IN1(m1stg_dblop_inv), .IN2(n1193), .IN3(m1stg_dblop), 
        .IN4(n973), .IN5(n10340), .Q(n10401) );
  AO22X1 U11224 ( .IN1(m1stg_dblop_inv), .IN2(n1195), .IN3(m1stg_dblop), .IN4(
        n977), .Q(n10340) );
  OA22X1 U11225 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n340 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n343 ), .Q(n10338) );
  AND2X1 U11226 ( .IN1(n10341), .IN2(n10337), .Q(n10398) );
  OA22X1 U11227 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n337 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n340 ), .Q(n10337) );
  OA22X1 U11228 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n338 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n341 ), .Q(n10341) );
  INVX0 U11229 ( .INP(n10400), .ZN(n10420) );
  NAND2X0 U11230 ( .IN1(n10333), .IN2(n10334), .QN(n10400) );
  OA22X1 U11231 ( .IN1(n1031), .IN2(\fpu_mul_frac_dp/n339 ), .IN3(n1032), 
        .IN4(\fpu_mul_frac_dp/n336 ), .Q(n10334) );
  OA22X1 U11232 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n335 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n338 ), .Q(n10333) );
  OA21X1 U11233 ( .IN1(n1221), .IN2(n987), .IN3(m1stg_dblop), .Q(n10362) );
  OA21X1 U11234 ( .IN1(n1222), .IN2(n985), .IN3(m1stg_dblop), .Q(n10438) );
  INVX0 U11235 ( .INP(n10391), .ZN(n10307) );
  NAND2X0 U11236 ( .IN1(n10444), .IN2(\fpu_mul_ctl/n263 ), .QN(n10391) );
  AO22X1 U11237 ( .IN1(n10445), .IN2(n10446), .IN3(n1395), .IN4(n1181), .Q(
        \fpu_mul_ctl/n405 ) );
  AO221X1 U11238 ( .IN1(n10447), .IN2(n10448), .IN3(n10449), .IN4(n10450), 
        .IN5(n10451), .Q(n10446) );
  MUX21X1 U11239 ( .IN1(n10452), .IN2(n10453), .S(n10454), .Q(n10451) );
  NAND2X0 U11240 ( .IN1(n10455), .IN2(n10456), .QN(n10453) );
  NAND4X0 U11241 ( .IN1(n10457), .IN2(\fpu_mul_frac_dp/n762 ), .IN3(n10458), 
        .IN4(n10459), .QN(n10456) );
  NAND2X0 U11242 ( .IN1(\fpu_mul_frac_dp/n749 ), .IN2(n941), .QN(n10458) );
  MUX21X1 U11243 ( .IN1(n10460), .IN2(n10461), .S(n10462), .Q(n10455) );
  NAND2X0 U11244 ( .IN1(\fpu_mul_frac_dp/n788 ), .IN2(n10463), .QN(n10461) );
  AO21X1 U11245 ( .IN1(\fpu_mul_frac_dp/n808 ), .IN2(n898), .IN3(n881), .Q(
        n10463) );
  OA21X1 U11246 ( .IN1(n10464), .IN2(n932), .IN3(n10465), .Q(n10460) );
  OA21X1 U11247 ( .IN1(n10466), .IN2(n930), .IN3(\fpu_mul_frac_dp/n804 ), .Q(
        n10464) );
  OA21X1 U11248 ( .IN1(\fpu_mul_frac_dp/n817 ), .IN2(n892), .IN3(
        \fpu_mul_frac_dp/n758 ), .Q(n10466) );
  NAND4X0 U11249 ( .IN1(n10467), .IN2(n10468), .IN3(n10469), .IN4(n10470), 
        .QN(n10452) );
  OA22X1 U11250 ( .IN1(n10471), .IN2(n10472), .IN3(n10473), .IN4(n10474), .Q(
        n10470) );
  NAND2X0 U11251 ( .IN1(\fpu_mul_frac_dp/n791 ), .IN2(n10475), .QN(n10474) );
  AO21X1 U11252 ( .IN1(n10476), .IN2(\fpu_mul_frac_dp/n793 ), .IN3(n897), .Q(
        n10475) );
  OA21X1 U11253 ( .IN1(n10477), .IN2(n10478), .IN3(n10479), .Q(n10471) );
  INVX0 U11254 ( .INP(n10480), .ZN(n10478) );
  OA21X1 U11255 ( .IN1(n10481), .IN2(n10482), .IN3(n10483), .Q(n10477) );
  INVX0 U11256 ( .INP(n10484), .ZN(n10482) );
  OA21X1 U11257 ( .IN1(n10485), .IN2(n10486), .IN3(n10487), .Q(n10481) );
  INVX0 U11258 ( .INP(n10488), .ZN(n10486) );
  OR2X1 U11259 ( .IN1(n10489), .IN2(n10490), .Q(n10469) );
  AO221X1 U11260 ( .IN1(n10491), .IN2(n10492), .IN3(n10493), .IN4(n10494), 
        .IN5(n10495), .Q(n10468) );
  NAND3X0 U11261 ( .IN1(n10496), .IN2(n10497), .IN3(n10498), .QN(n10494) );
  NAND2X0 U11262 ( .IN1(n10499), .IN2(n10500), .QN(n10498) );
  NAND4X0 U11263 ( .IN1(n10501), .IN2(\fpu_mul_frac_dp/n775 ), .IN3(n10502), 
        .IN4(n10503), .QN(n10467) );
  NAND2X0 U11264 ( .IN1(\fpu_mul_frac_dp/n809 ), .IN2(n940), .QN(n10502) );
  NAND2X0 U11265 ( .IN1(m1stg_dblop), .IN2(n10504), .QN(n10450) );
  AO21X1 U11266 ( .IN1(\fpu_mul_frac_dp/n790 ), .IN2(n939), .IN3(n896), .Q(
        n10504) );
  INVX0 U11267 ( .INP(n10505), .ZN(n10449) );
  INVX0 U11268 ( .INP(n10506), .ZN(n10448) );
  NOR2X0 U11269 ( .IN1(n10507), .IN2(n10508), .QN(n10447) );
  OA22X1 U11270 ( .IN1(n10509), .IN2(n10510), .IN3(n10511), .IN4(n10512), .Q(
        n10508) );
  OA21X1 U11271 ( .IN1(n10513), .IN2(n10514), .IN3(n10515), .Q(n10511) );
  INVX0 U11272 ( .INP(n10516), .ZN(n10514) );
  NAND2X0 U11273 ( .IN1(n10517), .IN2(n10518), .QN(n10510) );
  OAI21X1 U11274 ( .IN1(n887), .IN2(n10519), .IN3(n10520), .QN(n10518) );
  INVX0 U11275 ( .INP(n10521), .ZN(n10509) );
  OAI22X1 U11276 ( .IN1(n10522), .IN2(n10523), .IN3(\fpu_mul_ctl/n20 ), .IN4(
        n1625), .QN(\fpu_mul_ctl/n404 ) );
  OA221X1 U11277 ( .IN1(n10524), .IN2(n10525), .IN3(n10526), .IN4(n10506), 
        .IN5(n10527), .Q(n10522) );
  AO221X1 U11278 ( .IN1(n10528), .IN2(n10529), .IN3(n10530), .IN4(n10531), 
        .IN5(n10532), .Q(n10527) );
  NAND2X0 U11279 ( .IN1(\fpu_mul_frac_dp/n814 ), .IN2(\fpu_mul_frac_dp/n790 ), 
        .QN(n10531) );
  NAND3X0 U11280 ( .IN1(\fpu_mul_frac_dp/n780 ), .IN2(n10533), .IN3(
        \fpu_mul_frac_dp/n804 ), .QN(n10529) );
  NAND3X0 U11281 ( .IN1(\fpu_mul_frac_dp/n750 ), .IN2(n10534), .IN3(
        \fpu_mul_frac_dp/n758 ), .QN(n10533) );
  NAND3X0 U11282 ( .IN1(\fpu_mul_frac_dp/n783 ), .IN2(n10535), .IN3(
        \fpu_mul_frac_dp/n817 ), .QN(n10534) );
  NAND2X0 U11283 ( .IN1(n10536), .IN2(n10537), .QN(n10528) );
  NAND3X0 U11284 ( .IN1(\fpu_mul_frac_dp/n777 ), .IN2(n10538), .IN3(
        \fpu_mul_frac_dp/n808 ), .QN(n10537) );
  NAND2X0 U11285 ( .IN1(\fpu_mul_frac_dp/n762 ), .IN2(\fpu_mul_frac_dp/n749 ), 
        .QN(n10538) );
  OA21X1 U11286 ( .IN1(n10512), .IN2(n10539), .IN3(n10540), .Q(n10526) );
  NAND4X0 U11287 ( .IN1(n10521), .IN2(n10520), .IN3(n10517), .IN4(n10541), 
        .QN(n10540) );
  NAND2X0 U11288 ( .IN1(n10542), .IN2(n10543), .QN(n10541) );
  MUX21X1 U11289 ( .IN1(n10544), .IN2(n10545), .S(n10476), .Q(n10542) );
  NAND2X0 U11290 ( .IN1(\fpu_mul_frac_dp/n819 ), .IN2(\fpu_mul_frac_dp/n791 ), 
        .QN(n10545) );
  NAND2X0 U11291 ( .IN1(\fpu_mul_frac_dp/n809 ), .IN2(\fpu_mul_frac_dp/n775 ), 
        .QN(n10544) );
  AO21X1 U11292 ( .IN1(n10513), .IN2(n10516), .IN3(n10546), .Q(n10539) );
  INVX0 U11293 ( .INP(n10515), .ZN(n10546) );
  INVX0 U11294 ( .INP(n10547), .ZN(n10512) );
  OA22X1 U11295 ( .IN1(n10548), .IN2(n10549), .IN3(n10550), .IN4(n10489), .Q(
        n10525) );
  NAND3X0 U11296 ( .IN1(n10551), .IN2(n10552), .IN3(n10491), .QN(n10489) );
  INVX0 U11297 ( .INP(n10490), .ZN(n10550) );
  AO21X1 U11298 ( .IN1(n10553), .IN2(n10554), .IN3(n10495), .Q(n10549) );
  INVX0 U11299 ( .INP(n10555), .ZN(n10495) );
  NAND4X0 U11300 ( .IN1(n10492), .IN2(n10483), .IN3(n10480), .IN4(n10556), 
        .QN(n10554) );
  NAND3X0 U11301 ( .IN1(n10484), .IN2(n10557), .IN3(n10487), .QN(n10556) );
  NAND2X0 U11302 ( .IN1(n10485), .IN2(n10488), .QN(n10557) );
  INVX0 U11303 ( .INP(n10493), .ZN(n10548) );
  AO22X1 U11304 ( .IN1(n1631), .IN2(n1321), .IN3(n10558), .IN4(n10445), .Q(
        \fpu_mul_ctl/n403 ) );
  NOR2X0 U11305 ( .IN1(n10559), .IN2(n10560), .QN(n10558) );
  OA221X1 U11306 ( .IN1(n10462), .IN2(n10561), .IN3(n10562), .IN4(n10563), 
        .IN5(n10564), .Q(n10560) );
  INVX0 U11307 ( .INP(n10532), .ZN(n10564) );
  AO21X1 U11308 ( .IN1(n10565), .IN2(n10530), .IN3(n10566), .Q(n10532) );
  NAND2X0 U11309 ( .IN1(m1stg_dblop), .IN2(n10567), .QN(n10565) );
  NAND4X0 U11310 ( .IN1(\fpu_mul_frac_dp/n816 ), .IN2(\fpu_mul_frac_dp/n334 ), 
        .IN3(\fpu_mul_frac_dp/n814 ), .IN4(\fpu_mul_frac_dp/n790 ), .QN(n10567) );
  OA221X1 U11311 ( .IN1(n10476), .IN2(n10473), .IN3(n10568), .IN4(n10472), 
        .IN5(n10569), .Q(n10559) );
  OA22X1 U11312 ( .IN1(n10570), .IN2(n10571), .IN3(n10492), .IN4(n10572), .Q(
        n10569) );
  NAND2X0 U11313 ( .IN1(n10517), .IN2(n10573), .QN(n10571) );
  INVX0 U11314 ( .INP(n10524), .ZN(n10570) );
  INVX0 U11315 ( .INP(n10503), .ZN(n10476) );
  OAI22X1 U11316 ( .IN1(\fpu_mul_ctl/n18 ), .IN2(n1625), .IN3(n10574), .IN4(
        n10523), .QN(\fpu_mul_ctl/n402 ) );
  OA21X1 U11317 ( .IN1(n10575), .IN2(n10473), .IN3(n10472), .Q(n10574) );
  NAND3X0 U11318 ( .IN1(n10492), .IN2(n10576), .IN3(n10491), .QN(n10472) );
  INVX0 U11319 ( .INP(n10572), .ZN(n10491) );
  INVX0 U11320 ( .INP(n10552), .ZN(n10492) );
  OA21X1 U11321 ( .IN1(n10535), .IN2(n10530), .IN3(n10454), .Q(n10575) );
  AO22X1 U11322 ( .IN1(n1404), .IN2(n1322), .IN3(n10445), .IN4(n10577), .Q(
        \fpu_mul_ctl/n401 ) );
  NAND2X0 U11323 ( .IN1(n10506), .IN2(n10505), .QN(n10577) );
  NAND2X0 U11324 ( .IN1(n10454), .IN2(n10530), .QN(n10505) );
  AO21X1 U11325 ( .IN1(n10562), .IN2(n10457), .IN3(n1031), .Q(n10530) );
  INVX0 U11326 ( .INP(n10563), .ZN(n10457) );
  NAND3X0 U11327 ( .IN1(\fpu_mul_frac_dp/n777 ), .IN2(n10536), .IN3(
        \fpu_mul_frac_dp/n808 ), .QN(n10563) );
  NOR3X0 U11328 ( .IN1(n881), .IN2(n10535), .IN3(n925), .QN(n10536) );
  INVX0 U11329 ( .INP(n10462), .ZN(n10535) );
  NOR2X0 U11330 ( .IN1(n1113), .IN2(n10465), .QN(n10462) );
  OR4X1 U11331 ( .IN1(n1054), .IN2(n927), .IN3(n892), .IN4(n10561), .Q(n10465)
         );
  NAND4X0 U11332 ( .IN1(\fpu_mul_frac_dp/n804 ), .IN2(\fpu_mul_frac_dp/n780 ), 
        .IN3(\fpu_mul_frac_dp/n758 ), .IN4(\fpu_mul_frac_dp/n750 ), .QN(n10561) );
  INVX0 U11333 ( .INP(n10459), .ZN(n10562) );
  NAND4X0 U11334 ( .IN1(\fpu_mul_frac_dp/n801 ), .IN2(\fpu_mul_frac_dp/n784 ), 
        .IN3(\fpu_mul_frac_dp/n762 ), .IN4(\fpu_mul_frac_dp/n749 ), .QN(n10459) );
  NAND2X0 U11335 ( .IN1(n10524), .IN2(n10566), .QN(n10506) );
  AO22X1 U11336 ( .IN1(n10445), .IN2(n10454), .IN3(n1395), .IN4(n1162), .Q(
        \fpu_mul_ctl/n400 ) );
  INVX0 U11337 ( .INP(n10566), .ZN(n10454) );
  NAND3X0 U11338 ( .IN1(n10578), .IN2(n10503), .IN3(n10501), .QN(n10566) );
  INVX0 U11339 ( .INP(n10473), .ZN(n10501) );
  NAND2X0 U11340 ( .IN1(n10524), .IN2(n10507), .QN(n10473) );
  INVX0 U11341 ( .INP(n10573), .ZN(n10507) );
  NAND4X0 U11342 ( .IN1(n10521), .IN2(n10520), .IN3(n10517), .IN4(n10543), 
        .QN(n10573) );
  AOI221X1 U11343 ( .IN1(m1stg_dblop_inv), .IN2(n887), .IN3(
        \fpu_mul_frac_dp/n837 ), .IN4(m1stg_dblop), .IN5(n10519), .QN(n10543)
         );
  NOR2X0 U11344 ( .IN1(n1031), .IN2(\fpu_mul_frac_dp/n311 ), .QN(n10519) );
  AND4X1 U11345 ( .IN1(n10547), .IN2(n10513), .IN3(n10516), .IN4(n10515), .Q(
        n10517) );
  OA22X1 U11346 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n303 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n306 ), .Q(n10515) );
  OA22X1 U11347 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n776 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n307 ), .Q(n10516) );
  OA22X1 U11348 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n305 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n820 ), .Q(n10513) );
  OA22X1 U11349 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n812 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n305 ), .Q(n10547) );
  OA22X1 U11350 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n307 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n310 ), .Q(n10520) );
  OA22X1 U11351 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n306 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n309 ), .Q(n10521) );
  NOR3X0 U11352 ( .IN1(n10552), .IN2(n10576), .IN3(n10572), .QN(n10524) );
  NAND3X0 U11353 ( .IN1(n10493), .IN2(n10555), .IN3(n10553), .QN(n10572) );
  AND3X1 U11354 ( .IN1(n10496), .IN2(n10497), .IN3(n10499), .Q(n10553) );
  OA22X1 U11355 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n289 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n761 ), .Q(n10499) );
  NAND2X0 U11356 ( .IN1(m1stg_dblop_inv), .IN2(n942), .QN(n10497) );
  NAND2X0 U11357 ( .IN1(m1stg_dblop), .IN2(n891), .QN(n10496) );
  OA22X1 U11358 ( .IN1(n1031), .IN2(\fpu_mul_frac_dp/n289 ), .IN3(n1032), 
        .IN4(\fpu_mul_frac_dp/n286 ), .Q(n10555) );
  OA22X1 U11359 ( .IN1(n1031), .IN2(\fpu_mul_frac_dp/n818 ), .IN3(n1032), 
        .IN4(\fpu_mul_frac_dp/n287 ), .Q(n10493) );
  AO221X1 U11360 ( .IN1(m1stg_dblop_inv), .IN2(n889), .IN3(m1stg_dblop), .IN4(
        n909), .IN5(n10479), .Q(n10576) );
  NAND4X0 U11361 ( .IN1(n10485), .IN2(n10579), .IN3(n10580), .IN4(n10488), 
        .QN(n10479) );
  OA22X1 U11362 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n803 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n754 ), .Q(n10488) );
  OA22X1 U11363 ( .IN1(\fpu_mul_frac_dp/n300 ), .IN2(n1032), .IN3(
        \fpu_mul_frac_dp/n303 ), .IN4(n1031), .Q(n10580) );
  INVX0 U11364 ( .INP(n10568), .ZN(n10579) );
  NAND4X0 U11365 ( .IN1(n10487), .IN2(n10483), .IN3(n10480), .IN4(n10484), 
        .QN(n10568) );
  OA22X1 U11366 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n800 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n782 ), .Q(n10484) );
  OA22X1 U11367 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n811 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n779 ), .Q(n10480) );
  OA22X1 U11368 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n815 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n803 ), .Q(n10483) );
  OA22X1 U11369 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n779 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n300 ), .Q(n10487) );
  OA22X1 U11370 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n782 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n812 ), .Q(n10485) );
  AO221X1 U11371 ( .IN1(m1stg_dblop_inv), .IN2(n890), .IN3(m1stg_dblop), .IN4(
        n880), .IN5(n10500), .Q(n10552) );
  NAND3X0 U11372 ( .IN1(n10490), .IN2(n10551), .IN3(n10581), .QN(n10500) );
  OA22X1 U11373 ( .IN1(\fpu_mul_frac_dp/n761 ), .IN2(n1032), .IN3(
        \fpu_mul_frac_dp/n815 ), .IN4(n1031), .Q(n10581) );
  OA22X1 U11374 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n818 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n753 ), .Q(n10551) );
  OA22X1 U11375 ( .IN1(n1032), .IN2(\fpu_mul_frac_dp/n789 ), .IN3(n1031), 
        .IN4(\fpu_mul_frac_dp/n811 ), .Q(n10490) );
  NAND2X0 U11376 ( .IN1(m1stg_dblop), .IN2(n10582), .QN(n10503) );
  NAND4X0 U11377 ( .IN1(\fpu_mul_frac_dp/n826 ), .IN2(\fpu_mul_frac_dp/n819 ), 
        .IN3(\fpu_mul_frac_dp/n793 ), .IN4(\fpu_mul_frac_dp/n791 ), .QN(n10582) );
  NAND2X0 U11378 ( .IN1(m1stg_dblop), .IN2(n10583), .QN(n10578) );
  NAND4X0 U11379 ( .IN1(\fpu_mul_frac_dp/n822 ), .IN2(\fpu_mul_frac_dp/n809 ), 
        .IN3(\fpu_mul_frac_dp/n794 ), .IN4(\fpu_mul_frac_dp/n775 ), .QN(n10583) );
  INVX0 U11380 ( .INP(n10523), .ZN(n10445) );
  NAND2X0 U11381 ( .IN1(n10444), .IN2(\fpu_mul_ctl/n264 ), .QN(n10523) );
  OA21X1 U11382 ( .IN1(n886), .IN2(n910), .IN3(n1689), .Q(n10444) );
  NOR2X0 U11383 ( .IN1(n1679), .IN2(n1723), .QN(n1689) );
  NAND2X0 U11384 ( .IN1(n1882), .IN2(n1876), .QN(n1679) );
  NAND2X0 U11385 ( .IN1(n10584), .IN2(n1298), .QN(n1876) );
  NAND2X0 U11386 ( .IN1(n10584), .IN2(n1299), .QN(n1882) );
  NAND2X0 U11387 ( .IN1(\fpu_mul_ctl/n253 ), .IN2(n1037), .QN(n10584) );
  AO22X1 U11388 ( .IN1(n1404), .IN2(n1290), .IN3(n1593), .IN4(n10585), .Q(
        \fpu_mul_ctl/n399 ) );
  OAI21X1 U11389 ( .IN1(n974), .IN2(n1181), .IN3(n10586), .QN(n10585) );
  AO22X1 U11390 ( .IN1(n1631), .IN2(n1291), .IN3(n10587), .IN4(n1592), .Q(
        \fpu_mul_ctl/n398 ) );
  XOR3X1 U11391 ( .IN1(\fpu_mul_ctl/n26 ), .IN2(\fpu_mul_ctl/n20 ), .IN3(
        n10586), .Q(n10587) );
  AO22X1 U11392 ( .IN1(n1404), .IN2(n1292), .IN3(n1593), .IN4(n10588), .Q(
        \fpu_mul_ctl/n397 ) );
  XOR3X1 U11393 ( .IN1(\fpu_mul_ctl/n25 ), .IN2(\fpu_mul_ctl/n19 ), .IN3(
        n10589), .Q(n10588) );
  AO22X1 U11394 ( .IN1(n1405), .IN2(n1293), .IN3(n1593), .IN4(n10590), .Q(
        \fpu_mul_ctl/n396 ) );
  XOR3X1 U11395 ( .IN1(\fpu_mul_ctl/n18 ), .IN2(\fpu_mul_ctl/n24 ), .IN3(
        n10591), .Q(n10590) );
  AO22X1 U11396 ( .IN1(n1631), .IN2(n1294), .IN3(n1593), .IN4(n10592), .Q(
        \fpu_mul_ctl/n395 ) );
  XOR3X1 U11397 ( .IN1(\fpu_mul_ctl/n23 ), .IN2(\fpu_mul_ctl/n17 ), .IN3(
        n10593), .Q(n10592) );
  AO22X1 U11398 ( .IN1(n1404), .IN2(n1295), .IN3(n1593), .IN4(n10594), .Q(
        \fpu_mul_ctl/n394 ) );
  XOR2X1 U11399 ( .IN1(\fpu_mul_ctl/n22 ), .IN2(n10595), .Q(n10594) );
  OA21X1 U11400 ( .IN1(n10596), .IN2(n1162), .IN3(n10597), .Q(n10595) );
  AO22X1 U11401 ( .IN1(n1404), .IN2(n1296), .IN3(n1593), .IN4(n10598), .Q(
        \fpu_mul_ctl/n393 ) );
  AO22X1 U11402 ( .IN1(\fpu_mul_ctl/n16 ), .IN2(n10599), .IN3(
        \fpu_mul_ctl/n22 ), .IN4(n10597), .Q(n10598) );
  NAND2X0 U11403 ( .IN1(n1162), .IN2(n10596), .QN(n10597) );
  INVX0 U11404 ( .INP(n10599), .ZN(n10596) );
  OA22X1 U11405 ( .IN1(n10593), .IN2(\fpu_mul_ctl/n17 ), .IN3(n10600), .IN4(
        \fpu_mul_ctl/n23 ), .Q(n10599) );
  AND2X1 U11406 ( .IN1(n10593), .IN2(\fpu_mul_ctl/n17 ), .Q(n10600) );
  OA22X1 U11407 ( .IN1(n10591), .IN2(\fpu_mul_ctl/n18 ), .IN3(n10601), .IN4(
        \fpu_mul_ctl/n24 ), .Q(n10593) );
  AND2X1 U11408 ( .IN1(n10591), .IN2(\fpu_mul_ctl/n18 ), .Q(n10601) );
  OA22X1 U11409 ( .IN1(n10589), .IN2(\fpu_mul_ctl/n19 ), .IN3(n10602), .IN4(
        \fpu_mul_ctl/n25 ), .Q(n10591) );
  AND2X1 U11410 ( .IN1(n10589), .IN2(\fpu_mul_ctl/n19 ), .Q(n10602) );
  OA22X1 U11411 ( .IN1(n10586), .IN2(\fpu_mul_ctl/n20 ), .IN3(n10603), .IN4(
        \fpu_mul_ctl/n26 ), .Q(n10589) );
  AND2X1 U11412 ( .IN1(\fpu_mul_ctl/n20 ), .IN2(n10586), .Q(n10603) );
  NAND2X0 U11413 ( .IN1(n974), .IN2(n1181), .QN(n10586) );
  AO22X1 U11414 ( .IN1(n1599), .IN2(n1290), .IN3(m3bstg_ld0_inv[0]), .IN4(
        n1384), .Q(\fpu_mul_ctl/n392 ) );
  AO22X1 U11415 ( .IN1(n1599), .IN2(n1291), .IN3(m3bstg_ld0_inv[1]), .IN4(
        n1383), .Q(\fpu_mul_ctl/n391 ) );
  AO22X1 U11416 ( .IN1(n1599), .IN2(n1292), .IN3(m3bstg_ld0_inv[2]), .IN4(
        n1384), .Q(\fpu_mul_ctl/n390 ) );
  AO22X1 U11417 ( .IN1(n1599), .IN2(n1293), .IN3(m3bstg_ld0_inv[3]), .IN4(
        n1383), .Q(\fpu_mul_ctl/n389 ) );
  AO22X1 U11418 ( .IN1(n1599), .IN2(n1294), .IN3(m3bstg_ld0_inv[4]), .IN4(
        n1384), .Q(\fpu_mul_ctl/n388 ) );
  AO22X1 U11419 ( .IN1(n1596), .IN2(n1295), .IN3(m3bstg_ld0_inv[5]), .IN4(
        n1383), .Q(\fpu_mul_ctl/n387 ) );
  AO22X1 U11420 ( .IN1(n1598), .IN2(n1296), .IN3(m3bstg_ld0_inv[6]), .IN4(
        n1383), .Q(\fpu_mul_ctl/n386 ) );
  INVX0 U11421 ( .INP(n1723), .ZN(n604) );
  OAI22X1 U11422 ( .IN1(n10604), .IN2(n1723), .IN3(n1625), .IN4(
        \fpu_mul_ctl/n1 ), .QN(\fpu_mul_ctl/n385 ) );
  OAI22X1 U11423 ( .IN1(n8819), .IN2(n1723), .IN3(n1625), .IN4(
        m4stg_inc_exp_55), .QN(\fpu_mul_ctl/n384 ) );
  NAND2X0 U11424 ( .IN1(n1359), .IN2(n2929), .QN(n1723) );
  INVX0 U11425 ( .INP(n603), .ZN(n2929) );
  NAND2X0 U11426 ( .IN1(n8847), .IN2(n8838), .QN(n8819) );
  NAND2X0 U11427 ( .IN1(n1749), .IN2(n10604), .QN(n8838) );
  NAND4X0 U11428 ( .IN1(n10605), .IN2(n10606), .IN3(n10607), .IN4(n10608), 
        .QN(n10604) );
  NOR4X0 U11429 ( .IN1(n10609), .IN2(n10610), .IN3(n10611), .IN4(n10612), .QN(
        n10608) );
  XOR2X1 U11430 ( .IN1(n98), .IN2(m3stg_ld0_inv[0]), .Q(n10612) );
  XOR2X1 U11431 ( .IN1(n118), .IN2(m3stg_ld0_inv[5]), .Q(n10611) );
  XOR2X1 U11432 ( .IN1(n888), .IN2(n1059), .Q(n10610) );
  XOR2X1 U11433 ( .IN1(n106), .IN2(m3stg_ld0_inv[2]), .Q(n10609) );
  NOR3X0 U11434 ( .IN1(n10613), .IN2(n10614), .IN3(n1119), .QN(n10607) );
  XOR2X1 U11435 ( .IN1(n110), .IN2(m3stg_ld0_inv[3]), .Q(n10613) );
  XOR2X1 U11436 ( .IN1(m3stg_ld0_inv[6]), .IN2(n1114), .Q(n10606) );
  XOR2X1 U11437 ( .IN1(n1051), .IN2(n452), .Q(n10605) );
  XNOR2X1 U11438 ( .IN1(n10615), .IN2(n147), .Q(n1749) );
  NAND2X0 U11439 ( .IN1(n143), .IN2(n1747), .QN(n10615) );
  NOR2X0 U11440 ( .IN1(n1152), .IN2(n1745), .QN(n1747) );
  NAND2X0 U11441 ( .IN1(n135), .IN2(n1744), .QN(n1745) );
  INVX0 U11442 ( .INP(n1742), .ZN(n1744) );
  NAND2X0 U11443 ( .IN1(n453), .IN2(n1740), .QN(n1742) );
  NOR2X0 U11444 ( .IN1(n1153), .IN2(n1739), .QN(n1740) );
  AO22X1 U11445 ( .IN1(m3stg_ld0_inv[6]), .IN2(n1737), .IN3(n10616), .IN4(
        n1122), .Q(n1739) );
  OR2X1 U11446 ( .IN1(n1737), .IN2(m3stg_ld0_inv[6]), .Q(n10616) );
  AO22X1 U11447 ( .IN1(m3stg_ld0_inv[5]), .IN2(n10617), .IN3(n10618), .IN4(
        n1213), .Q(n1737) );
  NAND2X0 U11448 ( .IN1(n1735), .IN2(n1279), .QN(n10618) );
  INVX0 U11449 ( .INP(n10617), .ZN(n1735) );
  AO22X1 U11450 ( .IN1(m3stg_ld0_inv[4]), .IN2(n1733), .IN3(n10619), .IN4(
        n1211), .Q(n10617) );
  OR2X1 U11451 ( .IN1(n1733), .IN2(m3stg_ld0_inv[4]), .Q(n10619) );
  AO22X1 U11452 ( .IN1(m3stg_ld0_inv[3]), .IN2(n10620), .IN3(n10621), .IN4(
        n1214), .Q(n1733) );
  NAND2X0 U11453 ( .IN1(n1731), .IN2(n1280), .QN(n10621) );
  INVX0 U11454 ( .INP(n10620), .ZN(n1731) );
  AO22X1 U11455 ( .IN1(m3stg_ld0_inv[2]), .IN2(n1729), .IN3(n10622), .IN4(
        n1212), .Q(n10620) );
  NAND2X0 U11456 ( .IN1(n10623), .IN2(n1150), .QN(n10622) );
  INVX0 U11457 ( .INP(n10623), .ZN(n1729) );
  OA22X1 U11458 ( .IN1(n1051), .IN2(n1726), .IN3(n10624), .IN4(n103), .Q(
        n10623) );
  AND2X1 U11459 ( .IN1(n1726), .IN2(n1051), .Q(n10624) );
  NOR2X0 U11460 ( .IN1(n1154), .IN2(m3stg_ld0_inv[0]), .QN(n1726) );
  NAND2X0 U11461 ( .IN1(n146), .IN2(n10625), .QN(n8847) );
  NAND4X0 U11462 ( .IN1(n8845), .IN2(n10626), .IN3(n118), .IN4(n122), .QN(
        n10625) );
  INVX0 U11463 ( .INP(n10614), .ZN(n10626) );
  NAND4X0 U11464 ( .IN1(n142), .IN2(n138), .IN3(n10627), .IN4(n134), .QN(
        n10614) );
  NOR2X0 U11465 ( .IN1(n900), .IN2(n1203), .QN(n10627) );
  AND2X1 U11466 ( .IN1(n8827), .IN2(n114), .Q(n8845) );
  NOR2X0 U11467 ( .IN1(n8837), .IN2(n895), .QN(n8827) );
  NAND2X0 U11468 ( .IN1(n10628), .IN2(n110), .QN(n8837) );
  INVX0 U11469 ( .INP(n8830), .ZN(n10628) );
  NAND2X0 U11470 ( .IN1(n106), .IN2(n452), .QN(n8830) );
  NOR4X0 U11471 ( .IN1(\fpu_mul_ctl/n261 ), .IN2(n2928), .IN3(n1138), .IN4(
        n954), .QN(\fpu_mul_ctl/n380 ) );
  INVX0 U11472 ( .INP(n3131), .ZN(n2928) );
  NOR2X0 U11473 ( .IN1(n1702), .IN2(n1680), .QN(n3131) );
  INVX0 U11474 ( .INP(n10220), .ZN(n1680) );
  NAND3X0 U11475 ( .IN1(n10629), .IN2(n1206), .IN3(\fpu_mul_ctl/n269 ), .QN(
        n10220) );
  AND4X1 U11476 ( .IN1(\fpu_mul_ctl/n270 ), .IN2(\fpu_mul_ctl/n257 ), .IN3(
        n10629), .IN4(n1282), .Q(n1702) );
  AND4X1 U11477 ( .IN1(\fpu_mul_ctl/n96 ), .IN2(\fpu_mul_ctl/n94 ), .IN3(
        n10630), .IN4(\fpu_mul_ctl/n93 ), .Q(n10629) );
  NOR2X0 U11478 ( .IN1(\fpu_mul_ctl/n97 ), .IN2(\fpu_mul_ctl/n95 ), .QN(n10630) );
  NOR4X0 U11479 ( .IN1(\fpu_mul_ctl/m5stg_opdec[4] ), .IN2(n883), .IN3(n901), 
        .IN4(n1139), .QN(\fpu_mul_ctl/n379 ) );
  AO22X1 U11480 ( .IN1(n10217), .IN2(n1343), .IN3(inq_op[6]), .IN4(n10631), 
        .Q(\fpu_mul_ctl/i_m1stg_op/N9 ) );
  AO22X1 U11481 ( .IN1(n10217), .IN2(n1055), .IN3(inq_op[5]), .IN4(n10631), 
        .Q(\fpu_mul_ctl/i_m1stg_op/N8 ) );
  AO22X1 U11482 ( .IN1(n10217), .IN2(n1347), .IN3(inq_op[4]), .IN4(n10631), 
        .Q(\fpu_mul_ctl/i_m1stg_op/N7 ) );
  AO22X1 U11483 ( .IN1(n10217), .IN2(n1342), .IN3(inq_op[3]), .IN4(n10631), 
        .Q(\fpu_mul_ctl/i_m1stg_op/N6 ) );
  AO22X1 U11484 ( .IN1(n10217), .IN2(n1351), .IN3(inq_op[2]), .IN4(n10631), 
        .Q(\fpu_mul_ctl/i_m1stg_op/N5 ) );
  AO22X1 U11485 ( .IN1(n10217), .IN2(n1282), .IN3(n10631), .IN4(inq_op[1]), 
        .Q(\fpu_mul_ctl/i_m1stg_op/N4 ) );
  AO22X1 U11486 ( .IN1(n10217), .IN2(n1206), .IN3(n10631), .IN4(inq_op[0]), 
        .Q(\fpu_mul_ctl/i_m1stg_op/N3 ) );
  AO22X1 U11487 ( .IN1(n10217), .IN2(n1350), .IN3(inq_op[7]), .IN4(n10631), 
        .Q(\fpu_mul_ctl/i_m1stg_op/N10 ) );
  AO21X1 U11488 ( .IN1(n10217), .IN2(n1215), .IN3(n10631), .Q(
        \fpu_mul_ctl/i_m1stg_mul/N3 ) );
  AND3X1 U11489 ( .IN1(m1stg_step), .IN2(\fpu_mul_ctl/n735 ), .IN3(inq_mul), 
        .Q(n10631) );
  NOR2X0 U11490 ( .IN1(mul_rst_l), .IN2(se_mul), .QN(\fpu_mul_ctl/n735 ) );
  NOR2X0 U11491 ( .IN1(n1215), .IN2(n1798), .QN(m1stg_step) );
  NOR2X0 U11492 ( .IN1(mul_dest_rdya), .IN2(n1223), .QN(n1798) );
  INVX0 U11493 ( .INP(\fpu_mul_ctl/n105 ), .ZN(n10217) );
  NAND2X0 U11494 ( .IN1(n1405), .IN2(n1209), .QN(\fpu_mul_ctl/n105 ) );
  INVX0 U11495 ( .INP(n1625), .ZN(n1631) );
  NAND2X0 U11496 ( .IN1(n603), .IN2(n1357), .QN(n1625) );
  NOR2X0 U11497 ( .IN1(mul_dest_rdy), .IN2(n1223), .QN(n603) );
  AND2X1 U11498 ( .IN1(grst_l), .IN2(n1358), .Q(\fpu_mul_ctl/dffrl_mul_ctl/N4 ) );
endmodule

