
module fpu_out ( d8stg_fdiv_in, m6stg_fmul_in, a6stg_fadd_in, div_id_out_in, 
        m6stg_id_in, add_id_out_in, div_exc_out, d8stg_fdivd, d8stg_fdivs, 
        div_sign_out, div_exp_out, div_frac_out, mul_exc_out, 
        m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out, mul_exp_out, 
        mul_frac_out, add_exc_out, a6stg_fcmpop, add_cc_out, add_fcc_out, 
        a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst, a6stg_int_dst, 
        add_sign_out, add_exp_out, add_frac_out, arst_l, grst_l, rclk, 
        fp_cpx_req_cq, add_dest_rdy, mul_dest_rdy, div_dest_rdy, 
        fp_cpx_data_ca, se, si, so );
  input [9:0] div_id_out_in;
  input [9:0] m6stg_id_in;
  input [9:0] add_id_out_in;
  input [4:0] div_exc_out;
  input [10:0] div_exp_out;
  input [51:0] div_frac_out;
  input [4:0] mul_exc_out;
  input [10:0] mul_exp_out;
  input [51:0] mul_frac_out;
  input [4:0] add_exc_out;
  input [1:0] add_cc_out;
  input [1:0] add_fcc_out;
  input [10:0] add_exp_out;
  input [63:0] add_frac_out;
  output [7:0] fp_cpx_req_cq;
  output [144:0] fp_cpx_data_ca;
  input d8stg_fdiv_in, m6stg_fmul_in, a6stg_fadd_in, d8stg_fdivd, d8stg_fdivs,
         div_sign_out, m6stg_fmul_dbl_dst, m6stg_fmuls, mul_sign_out,
         a6stg_fcmpop, a6stg_dbl_dst, a6stg_sng_dst, a6stg_long_dst,
         a6stg_int_dst, add_sign_out, arst_l, grst_l, rclk, se, si;
  output add_dest_rdy, mul_dest_rdy, div_dest_rdy, so;
  wire   \fpu_out_ctl/out_ctl_rst_l , \fpu_out_ctl/dffrl_out_ctl/N4 ,
         \fpu_out_ctl/i_fp_cpx_req_cq/N10 , \fpu_out_ctl/i_fp_cpx_req_cq/N9 ,
         \fpu_out_ctl/i_fp_cpx_req_cq/N8 , \fpu_out_ctl/i_fp_cpx_req_cq/N7 ,
         \fpu_out_ctl/i_fp_cpx_req_cq/N6 , \fpu_out_ctl/i_fp_cpx_req_cq/N5 ,
         \fpu_out_ctl/i_fp_cpx_req_cq/N4 , \fpu_out_ctl/i_fp_cpx_req_cq/N3 ,
         \fpu_out_ctl/i_req_thread/N4 , \fpu_out_ctl/i_req_thread/N3 ,
         \fpu_out_ctl/i_dest_rdy/N3 , \fpu_out_ctl/i_mul_dest_rdy/N3 ,
         \fpu_out_dp/i_fp_cpx_data_ca_84_77/N9 ,
         \fpu_out_dp/i_fp_cpx_data_ca_84_77/N4 ,
         \fpu_out_dp/i_fp_cpx_data_ca_84_77/N3 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N79 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N78 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N77 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N76 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N75 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N72 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N71 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N70 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N69 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N68 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N66 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N65 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N64 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N63 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N62 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N61 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N60 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N59 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N58 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N57 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N56 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N55 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N54 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N53 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N52 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N51 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N50 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N49 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N48 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N47 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N46 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N45 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N44 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N43 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N42 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N41 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N40 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N39 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N38 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N37 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N36 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N35 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N34 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N33 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N32 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N31 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N30 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N29 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N28 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N27 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N26 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N25 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N24 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N23 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N22 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N21 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N20 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N19 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N18 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N17 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N16 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N15 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N14 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N13 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N12 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N11 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N10 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N9 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N8 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N7 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N6 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N5 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N4 ,
         \fpu_out_dp/i_fp_cpx_data_ca_76_0/N3 , n101, n102, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564;
  wire   [1:0] req_thread;
  assign fp_cpx_data_ca[143] = fp_cpx_data_ca[144];
  assign so = 1'b0;
  assign fp_cpx_data_ca[139] = 1'b0;
  assign fp_cpx_data_ca[138] = 1'b0;
  assign fp_cpx_data_ca[137] = 1'b0;
  assign fp_cpx_data_ca[133] = 1'b0;
  assign fp_cpx_data_ca[132] = 1'b0;
  assign fp_cpx_data_ca[131] = 1'b0;
  assign fp_cpx_data_ca[130] = 1'b0;
  assign fp_cpx_data_ca[129] = 1'b0;
  assign fp_cpx_data_ca[128] = 1'b0;
  assign fp_cpx_data_ca[127] = 1'b0;
  assign fp_cpx_data_ca[126] = 1'b0;
  assign fp_cpx_data_ca[125] = 1'b0;
  assign fp_cpx_data_ca[124] = 1'b0;
  assign fp_cpx_data_ca[123] = 1'b0;
  assign fp_cpx_data_ca[122] = 1'b0;
  assign fp_cpx_data_ca[121] = 1'b0;
  assign fp_cpx_data_ca[120] = 1'b0;
  assign fp_cpx_data_ca[119] = 1'b0;
  assign fp_cpx_data_ca[118] = 1'b0;
  assign fp_cpx_data_ca[117] = 1'b0;
  assign fp_cpx_data_ca[116] = 1'b0;
  assign fp_cpx_data_ca[115] = 1'b0;
  assign fp_cpx_data_ca[114] = 1'b0;
  assign fp_cpx_data_ca[113] = 1'b0;
  assign fp_cpx_data_ca[112] = 1'b0;
  assign fp_cpx_data_ca[111] = 1'b0;
  assign fp_cpx_data_ca[110] = 1'b0;
  assign fp_cpx_data_ca[109] = 1'b0;
  assign fp_cpx_data_ca[108] = 1'b0;
  assign fp_cpx_data_ca[107] = 1'b0;
  assign fp_cpx_data_ca[106] = 1'b0;
  assign fp_cpx_data_ca[105] = 1'b0;
  assign fp_cpx_data_ca[104] = 1'b0;
  assign fp_cpx_data_ca[103] = 1'b0;
  assign fp_cpx_data_ca[102] = 1'b0;
  assign fp_cpx_data_ca[101] = 1'b0;
  assign fp_cpx_data_ca[100] = 1'b0;
  assign fp_cpx_data_ca[99] = 1'b0;
  assign fp_cpx_data_ca[98] = 1'b0;
  assign fp_cpx_data_ca[97] = 1'b0;
  assign fp_cpx_data_ca[96] = 1'b0;
  assign fp_cpx_data_ca[95] = 1'b0;
  assign fp_cpx_data_ca[94] = 1'b0;
  assign fp_cpx_data_ca[93] = 1'b0;
  assign fp_cpx_data_ca[92] = 1'b0;
  assign fp_cpx_data_ca[91] = 1'b0;
  assign fp_cpx_data_ca[90] = 1'b0;
  assign fp_cpx_data_ca[89] = 1'b0;
  assign fp_cpx_data_ca[88] = 1'b0;
  assign fp_cpx_data_ca[87] = 1'b0;
  assign fp_cpx_data_ca[86] = 1'b0;
  assign fp_cpx_data_ca[85] = 1'b0;
  assign fp_cpx_data_ca[84] = 1'b0;
  assign fp_cpx_data_ca[83] = 1'b0;
  assign fp_cpx_data_ca[82] = 1'b0;
  assign fp_cpx_data_ca[81] = 1'b0;
  assign fp_cpx_data_ca[80] = 1'b0;
  assign fp_cpx_data_ca[79] = 1'b0;
  assign fp_cpx_data_ca[78] = 1'b0;
  assign fp_cpx_data_ca[77] = 1'b0;
  assign fp_cpx_data_ca[64] = 1'b0;
  assign fp_cpx_data_ca[70] = 1'b0;
  assign fp_cpx_data_ca[71] = 1'b0;
  assign fp_cpx_data_ca[136] = 1'b0;
  assign fp_cpx_data_ca[140] = 1'b0;
  assign fp_cpx_data_ca[141] = 1'b0;
  assign fp_cpx_data_ca[142] = 1'b0;

  DFFARX1 \fpu_out_ctl/dffrl_out_ctl/q_reg[0]  ( .D(
        \fpu_out_ctl/dffrl_out_ctl/N4 ), .CLK(rclk), .RSTB(arst_l), .Q(
        \fpu_out_ctl/out_ctl_rst_l ) );
  DFFX1 \fpu_out_ctl/i_add_req/q_reg[0]  ( .D(n283), .CLK(rclk), .Q(n396), 
        .QN(n102) );
  DFFX1 \fpu_out_ctl/i_fp_cpx_req_cq/q_reg[0]  ( .D(
        \fpu_out_ctl/i_fp_cpx_req_cq/N3 ), .CLK(rclk), .Q(fp_cpx_req_cq[0]) );
  DFFX1 \fpu_out_ctl/i_fp_cpx_req_cq/q_reg[1]  ( .D(
        \fpu_out_ctl/i_fp_cpx_req_cq/N4 ), .CLK(rclk), .Q(fp_cpx_req_cq[1]) );
  DFFX1 \fpu_out_ctl/i_fp_cpx_req_cq/q_reg[2]  ( .D(
        \fpu_out_ctl/i_fp_cpx_req_cq/N5 ), .CLK(rclk), .Q(fp_cpx_req_cq[2]) );
  DFFX1 \fpu_out_ctl/i_fp_cpx_req_cq/q_reg[3]  ( .D(
        \fpu_out_ctl/i_fp_cpx_req_cq/N6 ), .CLK(rclk), .Q(fp_cpx_req_cq[3]) );
  DFFX1 \fpu_out_ctl/i_fp_cpx_req_cq/q_reg[4]  ( .D(
        \fpu_out_ctl/i_fp_cpx_req_cq/N7 ), .CLK(rclk), .Q(fp_cpx_req_cq[4]) );
  DFFX1 \fpu_out_ctl/i_fp_cpx_req_cq/q_reg[5]  ( .D(
        \fpu_out_ctl/i_fp_cpx_req_cq/N8 ), .CLK(rclk), .Q(fp_cpx_req_cq[5]) );
  DFFX1 \fpu_out_ctl/i_fp_cpx_req_cq/q_reg[6]  ( .D(
        \fpu_out_ctl/i_fp_cpx_req_cq/N9 ), .CLK(rclk), .Q(fp_cpx_req_cq[6]) );
  DFFX1 \fpu_out_ctl/i_fp_cpx_req_cq/q_reg[7]  ( .D(
        \fpu_out_ctl/i_fp_cpx_req_cq/N10 ), .CLK(rclk), .Q(fp_cpx_req_cq[7])
         );
  DFFX1 \fpu_out_ctl/i_req_thread/q_reg[0]  ( .D(\fpu_out_ctl/i_req_thread/N3 ), .CLK(rclk), .Q(req_thread[0]) );
  DFFX1 \fpu_out_ctl/i_req_thread/q_reg[1]  ( .D(\fpu_out_ctl/i_req_thread/N4 ), .CLK(rclk), .Q(req_thread[1]) );
  DFFX1 \fpu_out_ctl/i_add_dest_rdy/q_reg[0]  ( .D(\fpu_out_ctl/i_dest_rdy/N3 ), .CLK(rclk), .Q(add_dest_rdy) );
  DFFX1 \fpu_out_ctl/i_mul_dest_rdy/q_reg[0]  ( .D(
        \fpu_out_ctl/i_mul_dest_rdy/N3 ), .CLK(rclk), .Q(mul_dest_rdy) );
  DFFSSRX1 \fpu_out_ctl/i_div_dest_rdy/q_reg[0]  ( .D(n101), .RSTB(
        d8stg_fdiv_in), .SETB(1'b1), .CLK(rclk), .Q(div_dest_rdy) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_84_77/q_reg[0]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_84_77/N3 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[134]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_84_77/q_reg[1]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_84_77/N4 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[135]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_84_77/q_reg[7]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_84_77/N9 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[144]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[0]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N3 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[0]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[1]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N4 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[1]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[2]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N5 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[2]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[3]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N6 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[3]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[4]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N7 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[4]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[5]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N8 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[5]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[6]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N9 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[6]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[7]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N10 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[7]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[8]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N11 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[8]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[9]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N12 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[9]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[10]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N13 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[10]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[11]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N14 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[11]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[12]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N15 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[12]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[13]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N16 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[13]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[14]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N17 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[14]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[15]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N18 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[15]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[16]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N19 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[16]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[17]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N20 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[17]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[18]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N21 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[18]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[19]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N22 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[19]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[20]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N23 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[20]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[21]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N24 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[21]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[22]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N25 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[22]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[23]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N26 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[23]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[24]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N27 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[24]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[25]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N28 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[25]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[26]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N29 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[26]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[27]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N30 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[27]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[28]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N31 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[28]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[29]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N32 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[29]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[30]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N33 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[30]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[31]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N34 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[31]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[32]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N35 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[32]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[33]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N36 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[33]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[34]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N37 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[34]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[35]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N38 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[35]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[36]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N39 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[36]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[37]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N40 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[37]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[38]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N41 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[38]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[39]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N42 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[39]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[40]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N43 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[40]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[41]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N44 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[41]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[42]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N45 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[42]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[43]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N46 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[43]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[44]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N47 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[44]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[45]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N48 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[45]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[46]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N49 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[46]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[47]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N50 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[47]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[48]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N51 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[48]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[49]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N52 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[49]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[50]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N53 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[50]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[51]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N54 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[51]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[52]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N55 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[52]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[53]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N56 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[53]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[54]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N57 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[54]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[55]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N58 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[55]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[56]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N59 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[56]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[57]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N60 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[57]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[58]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N61 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[58]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[59]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N62 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[59]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[60]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N63 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[60]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[61]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N64 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[61]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[62]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N65 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[62]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[63]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N66 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[63]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[65]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N68 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[65]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[66]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N69 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[66]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[67]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N70 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[67]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[68]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N71 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[68]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[69]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N72 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[69]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[72]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N75 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[72]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[73]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N76 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[73]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[74]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N77 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[74]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[75]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N78 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[75]) );
  DFFX1 \fpu_out_dp/i_fp_cpx_data_ca_76_0/q_reg[76]  ( .D(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N79 ), .CLK(rclk), .Q(
        fp_cpx_data_ca[76]) );
  OA221X1 U280 ( .IN1(1'b0), .IN2(\fpu_out_ctl/out_ctl_rst_l ), .IN3(n386), 
        .IN4(n102), .IN5(n387), .Q(n283) );
  INVX0 U281 ( .INP(n562), .ZN(n559) );
  INVX0 U282 ( .INP(n560), .ZN(n558) );
  INVX0 U283 ( .INP(n561), .ZN(n557) );
  NAND2X1 U284 ( .IN1(n559), .IN2(m6stg_fmuls), .QN(n555) );
  INVX0 U285 ( .INP(n555), .ZN(n397) );
  INVX2 U286 ( .INP(n556), .ZN(n389) );
  NOR2X0 U287 ( .IN1(se), .IN2(n563), .QN(n398) );
  INVX0 U288 ( .INP(d8stg_fdiv_in), .ZN(n563) );
  INVX0 U289 ( .INP(se), .ZN(n101) );
  NOR2X0 U290 ( .IN1(se), .IN2(n564), .QN(\fpu_out_ctl/i_mul_dest_rdy/N3 ) );
  NAND2X0 U291 ( .IN1(n396), .IN2(a6stg_fadd_in), .QN(n284) );
  NAND3X0 U292 ( .IN1(n284), .IN2(m6stg_fmul_in), .IN3(n563), .QN(n564) );
  NAND2X0 U293 ( .IN1(n102), .IN2(m6stg_fmul_in), .QN(n285) );
  AND4X1 U294 ( .IN1(n101), .IN2(n563), .IN3(a6stg_fadd_in), .IN4(n285), .Q(
        \fpu_out_ctl/i_dest_rdy/N3 ) );
  NAND2X0 U295 ( .IN1(n555), .IN2(n556), .QN(n286) );
  OR2X1 U296 ( .IN1(n392), .IN2(n390), .Q(n287) );
  AO222X1 U297 ( .IN1(n286), .IN2(mul_sign_out), .IN3(n287), .IN4(add_sign_out), .IN5(add_frac_out[63]), .IN6(n395), .Q(n288) );
  AO221X1 U298 ( .IN1(div_sign_out), .IN2(n391), .IN3(div_sign_out), .IN4(n394), .IN5(n288), .Q(\fpu_out_dp/i_fp_cpx_data_ca_76_0/N66 ) );
  NAND2X0 U299 ( .IN1(n392), .IN2(add_frac_out[42]), .QN(n289) );
  NAND2X0 U300 ( .IN1(n393), .IN2(add_frac_out[31]), .QN(n290) );
  NAND2X0 U301 ( .IN1(n389), .IN2(mul_frac_out[31]), .QN(n291) );
  NAND2X0 U302 ( .IN1(n391), .IN2(div_frac_out[31]), .QN(n292) );
  NAND4X0 U303 ( .IN1(n289), .IN2(n290), .IN3(n291), .IN4(n292), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N34 ) );
  NAND2X0 U304 ( .IN1(n392), .IN2(add_frac_out[38]), .QN(n293) );
  NAND2X0 U305 ( .IN1(n393), .IN2(add_frac_out[27]), .QN(n294) );
  NAND2X0 U306 ( .IN1(n389), .IN2(mul_frac_out[27]), .QN(n295) );
  NAND2X0 U307 ( .IN1(n391), .IN2(div_frac_out[27]), .QN(n296) );
  NAND4X0 U308 ( .IN1(n293), .IN2(n294), .IN3(n295), .IN4(n296), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N30 ) );
  NAND2X0 U309 ( .IN1(n392), .IN2(add_frac_out[37]), .QN(n297) );
  NAND2X0 U310 ( .IN1(n393), .IN2(add_frac_out[26]), .QN(n298) );
  NAND2X0 U311 ( .IN1(n389), .IN2(mul_frac_out[26]), .QN(n299) );
  NAND2X0 U312 ( .IN1(n391), .IN2(div_frac_out[26]), .QN(n300) );
  NAND4X0 U313 ( .IN1(n297), .IN2(n298), .IN3(n299), .IN4(n300), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N29 ) );
  NAND2X0 U314 ( .IN1(n392), .IN2(add_frac_out[36]), .QN(n301) );
  NAND2X0 U315 ( .IN1(n393), .IN2(add_frac_out[25]), .QN(n302) );
  NAND2X0 U316 ( .IN1(n389), .IN2(mul_frac_out[25]), .QN(n303) );
  NAND2X0 U317 ( .IN1(n391), .IN2(div_frac_out[25]), .QN(n304) );
  NAND4X0 U318 ( .IN1(n301), .IN2(n302), .IN3(n303), .IN4(n304), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N28 ) );
  NAND2X0 U319 ( .IN1(n392), .IN2(add_frac_out[35]), .QN(n305) );
  NAND2X0 U320 ( .IN1(n393), .IN2(add_frac_out[24]), .QN(n306) );
  NAND2X0 U321 ( .IN1(n389), .IN2(mul_frac_out[24]), .QN(n307) );
  NAND2X0 U322 ( .IN1(n391), .IN2(div_frac_out[24]), .QN(n308) );
  NAND4X0 U323 ( .IN1(n305), .IN2(n306), .IN3(n307), .IN4(n308), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N27 ) );
  NAND2X0 U324 ( .IN1(n392), .IN2(add_frac_out[34]), .QN(n309) );
  NAND2X0 U325 ( .IN1(n393), .IN2(add_frac_out[23]), .QN(n310) );
  NAND2X0 U326 ( .IN1(n389), .IN2(mul_frac_out[23]), .QN(n311) );
  NAND2X0 U327 ( .IN1(n391), .IN2(div_frac_out[23]), .QN(n312) );
  NAND4X0 U328 ( .IN1(n309), .IN2(n310), .IN3(n311), .IN4(n312), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N26 ) );
  NAND2X0 U329 ( .IN1(n392), .IN2(add_frac_out[33]), .QN(n313) );
  NAND2X0 U330 ( .IN1(n393), .IN2(add_frac_out[22]), .QN(n314) );
  NAND2X0 U331 ( .IN1(n389), .IN2(mul_frac_out[22]), .QN(n315) );
  NAND2X0 U332 ( .IN1(n391), .IN2(div_frac_out[22]), .QN(n316) );
  NAND4X0 U333 ( .IN1(n313), .IN2(n314), .IN3(n315), .IN4(n316), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N25 ) );
  NAND2X0 U334 ( .IN1(n392), .IN2(add_frac_out[32]), .QN(n317) );
  NAND2X0 U335 ( .IN1(n393), .IN2(add_frac_out[21]), .QN(n318) );
  NAND2X0 U336 ( .IN1(n389), .IN2(mul_frac_out[21]), .QN(n319) );
  NAND2X0 U337 ( .IN1(n391), .IN2(div_frac_out[21]), .QN(n320) );
  NAND4X0 U338 ( .IN1(n317), .IN2(n318), .IN3(n319), .IN4(n320), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N24 ) );
  NAND2X0 U339 ( .IN1(n392), .IN2(add_frac_out[31]), .QN(n321) );
  NAND2X0 U340 ( .IN1(n393), .IN2(add_frac_out[20]), .QN(n322) );
  NAND2X0 U341 ( .IN1(n389), .IN2(mul_frac_out[20]), .QN(n323) );
  NAND2X0 U342 ( .IN1(n391), .IN2(div_frac_out[20]), .QN(n324) );
  NAND4X0 U343 ( .IN1(n321), .IN2(n322), .IN3(n323), .IN4(n324), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N23 ) );
  NAND2X0 U344 ( .IN1(n392), .IN2(add_frac_out[25]), .QN(n325) );
  NAND2X0 U345 ( .IN1(n393), .IN2(add_frac_out[14]), .QN(n326) );
  NAND2X0 U346 ( .IN1(n389), .IN2(mul_frac_out[14]), .QN(n327) );
  NAND2X0 U347 ( .IN1(n391), .IN2(div_frac_out[14]), .QN(n328) );
  NAND4X0 U348 ( .IN1(n325), .IN2(n326), .IN3(n327), .IN4(n328), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N17 ) );
  NAND2X0 U349 ( .IN1(n392), .IN2(add_frac_out[24]), .QN(n329) );
  NAND2X0 U350 ( .IN1(n393), .IN2(add_frac_out[13]), .QN(n330) );
  NAND2X0 U351 ( .IN1(n389), .IN2(mul_frac_out[13]), .QN(n331) );
  NAND2X0 U352 ( .IN1(n391), .IN2(div_frac_out[13]), .QN(n332) );
  NAND4X0 U353 ( .IN1(n329), .IN2(n330), .IN3(n331), .IN4(n332), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N16 ) );
  NAND2X0 U354 ( .IN1(n392), .IN2(add_frac_out[23]), .QN(n333) );
  NAND2X0 U355 ( .IN1(n393), .IN2(add_frac_out[12]), .QN(n334) );
  NAND2X0 U356 ( .IN1(n389), .IN2(mul_frac_out[12]), .QN(n335) );
  NAND2X0 U357 ( .IN1(n391), .IN2(div_frac_out[12]), .QN(n336) );
  NAND4X0 U358 ( .IN1(n333), .IN2(n334), .IN3(n335), .IN4(n336), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N15 ) );
  NAND2X0 U359 ( .IN1(n392), .IN2(add_frac_out[22]), .QN(n337) );
  NAND2X0 U360 ( .IN1(n393), .IN2(add_frac_out[11]), .QN(n338) );
  NAND2X0 U361 ( .IN1(n389), .IN2(mul_frac_out[11]), .QN(n339) );
  NAND2X0 U362 ( .IN1(n391), .IN2(div_frac_out[11]), .QN(n340) );
  NAND4X0 U363 ( .IN1(n337), .IN2(n338), .IN3(n339), .IN4(n340), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N14 ) );
  NAND2X0 U364 ( .IN1(n392), .IN2(add_frac_out[21]), .QN(n341) );
  NAND2X0 U365 ( .IN1(n393), .IN2(add_frac_out[10]), .QN(n342) );
  NAND2X0 U366 ( .IN1(n389), .IN2(mul_frac_out[10]), .QN(n343) );
  NAND2X0 U367 ( .IN1(n391), .IN2(div_frac_out[10]), .QN(n344) );
  NAND4X0 U368 ( .IN1(n341), .IN2(n342), .IN3(n343), .IN4(n344), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N13 ) );
  NAND2X0 U369 ( .IN1(n392), .IN2(add_frac_out[20]), .QN(n345) );
  NAND2X0 U370 ( .IN1(n393), .IN2(add_frac_out[9]), .QN(n346) );
  NAND2X0 U371 ( .IN1(n389), .IN2(mul_frac_out[9]), .QN(n347) );
  NAND2X0 U372 ( .IN1(n391), .IN2(div_frac_out[9]), .QN(n348) );
  NAND4X0 U373 ( .IN1(n345), .IN2(n346), .IN3(n347), .IN4(n348), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N12 ) );
  NAND2X0 U374 ( .IN1(n392), .IN2(add_frac_out[19]), .QN(n349) );
  NAND2X0 U375 ( .IN1(n393), .IN2(add_frac_out[8]), .QN(n350) );
  NAND2X0 U376 ( .IN1(n389), .IN2(mul_frac_out[8]), .QN(n351) );
  NAND2X0 U377 ( .IN1(n391), .IN2(div_frac_out[8]), .QN(n352) );
  NAND4X0 U378 ( .IN1(n349), .IN2(n350), .IN3(n351), .IN4(n352), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N11 ) );
  NAND2X0 U379 ( .IN1(n392), .IN2(add_frac_out[18]), .QN(n353) );
  NAND2X0 U380 ( .IN1(n393), .IN2(add_frac_out[7]), .QN(n354) );
  NAND2X0 U381 ( .IN1(n389), .IN2(mul_frac_out[7]), .QN(n355) );
  NAND2X0 U382 ( .IN1(n391), .IN2(div_frac_out[7]), .QN(n356) );
  NAND4X0 U383 ( .IN1(n353), .IN2(n354), .IN3(n355), .IN4(n356), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N10 ) );
  NAND2X0 U384 ( .IN1(n392), .IN2(add_frac_out[17]), .QN(n357) );
  NAND2X0 U385 ( .IN1(n393), .IN2(add_frac_out[6]), .QN(n358) );
  NAND2X0 U386 ( .IN1(n389), .IN2(mul_frac_out[6]), .QN(n359) );
  NAND2X0 U387 ( .IN1(n391), .IN2(div_frac_out[6]), .QN(n360) );
  NAND4X0 U388 ( .IN1(n357), .IN2(n358), .IN3(n359), .IN4(n360), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N9 ) );
  NAND2X0 U389 ( .IN1(n392), .IN2(add_frac_out[16]), .QN(n361) );
  NAND2X0 U390 ( .IN1(n393), .IN2(add_frac_out[5]), .QN(n362) );
  NAND2X0 U391 ( .IN1(n389), .IN2(mul_frac_out[5]), .QN(n363) );
  NAND2X0 U392 ( .IN1(n391), .IN2(div_frac_out[5]), .QN(n364) );
  NAND4X0 U393 ( .IN1(n361), .IN2(n362), .IN3(n363), .IN4(n364), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N8 ) );
  NAND2X0 U394 ( .IN1(n392), .IN2(add_frac_out[15]), .QN(n365) );
  NAND2X0 U395 ( .IN1(n393), .IN2(add_frac_out[4]), .QN(n366) );
  NAND2X0 U396 ( .IN1(n389), .IN2(mul_frac_out[4]), .QN(n367) );
  NAND2X0 U397 ( .IN1(n391), .IN2(div_frac_out[4]), .QN(n368) );
  NAND4X0 U398 ( .IN1(n365), .IN2(n366), .IN3(n367), .IN4(n368), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N7 ) );
  NAND2X0 U399 ( .IN1(n392), .IN2(add_frac_out[14]), .QN(n369) );
  NAND2X0 U400 ( .IN1(n393), .IN2(add_frac_out[3]), .QN(n370) );
  NAND2X0 U401 ( .IN1(n389), .IN2(mul_frac_out[3]), .QN(n371) );
  NAND2X0 U402 ( .IN1(n391), .IN2(div_frac_out[3]), .QN(n372) );
  NAND4X0 U403 ( .IN1(n369), .IN2(n370), .IN3(n371), .IN4(n372), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N6 ) );
  NAND2X0 U404 ( .IN1(n392), .IN2(add_frac_out[13]), .QN(n373) );
  NAND2X0 U405 ( .IN1(n393), .IN2(add_frac_out[2]), .QN(n374) );
  NAND2X0 U406 ( .IN1(n389), .IN2(mul_frac_out[2]), .QN(n375) );
  NAND2X0 U407 ( .IN1(n391), .IN2(div_frac_out[2]), .QN(n376) );
  NAND4X0 U408 ( .IN1(n373), .IN2(n374), .IN3(n375), .IN4(n376), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N5 ) );
  NAND2X0 U409 ( .IN1(n392), .IN2(add_frac_out[12]), .QN(n377) );
  NAND2X0 U410 ( .IN1(n393), .IN2(add_frac_out[1]), .QN(n378) );
  NAND2X0 U411 ( .IN1(n389), .IN2(mul_frac_out[1]), .QN(n379) );
  NAND2X0 U412 ( .IN1(n391), .IN2(div_frac_out[1]), .QN(n380) );
  NAND4X0 U413 ( .IN1(n377), .IN2(n378), .IN3(n379), .IN4(n380), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N4 ) );
  NAND2X0 U414 ( .IN1(n392), .IN2(add_frac_out[11]), .QN(n381) );
  NAND2X0 U415 ( .IN1(n393), .IN2(add_frac_out[0]), .QN(n382) );
  NAND2X0 U416 ( .IN1(n389), .IN2(mul_frac_out[0]), .QN(n383) );
  NAND2X0 U417 ( .IN1(n391), .IN2(div_frac_out[0]), .QN(n384) );
  NAND4X0 U418 ( .IN1(n381), .IN2(n382), .IN3(n383), .IN4(n384), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N3 ) );
  NAND2X0 U419 ( .IN1(n563), .IN2(a6stg_fadd_in), .QN(n385) );
  AND3X1 U420 ( .IN1(n101), .IN2(n564), .IN3(n385), .Q(n386) );
  OR3X1 U421 ( .IN1(\fpu_out_ctl/i_dest_rdy/N3 ), .IN2(
        \fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN3(n396), .Q(n387) );
  NAND2X1 U423 ( .IN1(mul_dest_rdy), .IN2(n101), .QN(n562) );
  NAND2X1 U424 ( .IN1(add_dest_rdy), .IN2(n101), .QN(n561) );
  NAND2X1 U425 ( .IN1(div_dest_rdy), .IN2(n101), .QN(n560) );
  AND2X1 U426 ( .IN1(n557), .IN2(a6stg_long_dst), .Q(n393) );
  OA21X1 U427 ( .IN1(a6stg_long_dst), .IN2(a6stg_int_dst), .IN3(n557), .Q(n395) );
  AND2X1 U428 ( .IN1(n557), .IN2(a6stg_dbl_dst), .Q(n392) );
  AND2X1 U429 ( .IN1(n557), .IN2(a6stg_sng_dst), .Q(n390) );
  AND2X1 U430 ( .IN1(n558), .IN2(d8stg_fdivd), .Q(n391) );
  AND2X1 U431 ( .IN1(n558), .IN2(d8stg_fdivs), .Q(n394) );
  NAND2X1 U432 ( .IN1(n393), .IN2(add_frac_out[15]), .QN(n399) );
  NAND2X1 U433 ( .IN1(n392), .IN2(add_frac_out[26]), .QN(n400) );
  NAND2X1 U434 ( .IN1(n391), .IN2(div_frac_out[15]), .QN(n401) );
  NAND2X1 U435 ( .IN1(n389), .IN2(mul_frac_out[15]), .QN(n402) );
  NAND2X1 U436 ( .IN1(n393), .IN2(add_frac_out[16]), .QN(n403) );
  NAND2X1 U437 ( .IN1(n392), .IN2(add_frac_out[27]), .QN(n404) );
  NAND2X1 U438 ( .IN1(n391), .IN2(div_frac_out[16]), .QN(n405) );
  NAND2X1 U439 ( .IN1(n389), .IN2(mul_frac_out[16]), .QN(n406) );
  NAND2X1 U440 ( .IN1(n393), .IN2(add_frac_out[17]), .QN(n407) );
  NAND2X1 U441 ( .IN1(n392), .IN2(add_frac_out[28]), .QN(n408) );
  NAND2X1 U442 ( .IN1(n391), .IN2(div_frac_out[17]), .QN(n409) );
  NAND2X1 U443 ( .IN1(n389), .IN2(mul_frac_out[17]), .QN(n410) );
  NAND2X1 U444 ( .IN1(add_frac_out[18]), .IN2(n393), .QN(n411) );
  NAND2X1 U445 ( .IN1(n392), .IN2(add_frac_out[29]), .QN(n412) );
  NAND2X1 U446 ( .IN1(n391), .IN2(div_frac_out[18]), .QN(n413) );
  NAND2X1 U447 ( .IN1(n389), .IN2(mul_frac_out[18]), .QN(n414) );
  NAND2X1 U448 ( .IN1(n393), .IN2(add_frac_out[19]), .QN(n415) );
  NAND2X1 U449 ( .IN1(n392), .IN2(add_frac_out[30]), .QN(n416) );
  NAND2X1 U450 ( .IN1(n391), .IN2(div_frac_out[19]), .QN(n417) );
  NAND2X1 U451 ( .IN1(n389), .IN2(mul_frac_out[19]), .QN(n418) );
  NAND2X1 U452 ( .IN1(n393), .IN2(add_frac_out[28]), .QN(n419) );
  NAND2X1 U453 ( .IN1(n392), .IN2(add_frac_out[39]), .QN(n420) );
  NAND2X1 U454 ( .IN1(n391), .IN2(div_frac_out[28]), .QN(n421) );
  NAND2X1 U455 ( .IN1(n389), .IN2(mul_frac_out[28]), .QN(n422) );
  NAND2X1 U456 ( .IN1(n393), .IN2(add_frac_out[29]), .QN(n423) );
  NAND2X1 U457 ( .IN1(add_frac_out[40]), .IN2(n392), .QN(n424) );
  NAND2X1 U458 ( .IN1(div_frac_out[29]), .IN2(n391), .QN(n425) );
  NAND2X1 U459 ( .IN1(n389), .IN2(mul_frac_out[29]), .QN(n426) );
  NAND2X1 U460 ( .IN1(n393), .IN2(add_frac_out[30]), .QN(n427) );
  NAND2X1 U461 ( .IN1(n392), .IN2(add_frac_out[41]), .QN(n428) );
  NAND2X1 U462 ( .IN1(n391), .IN2(div_frac_out[30]), .QN(n429) );
  NAND2X1 U463 ( .IN1(n389), .IN2(mul_frac_out[30]), .QN(n430) );
  NAND2X1 U464 ( .IN1(n389), .IN2(mul_frac_out[32]), .QN(n431) );
  NAND2X1 U465 ( .IN1(n389), .IN2(mul_frac_out[33]), .QN(n435) );
  NAND2X1 U466 ( .IN1(n389), .IN2(mul_frac_out[34]), .QN(n439) );
  NAND2X1 U467 ( .IN1(n389), .IN2(mul_frac_out[35]), .QN(n443) );
  NAND2X1 U468 ( .IN1(n389), .IN2(mul_frac_out[36]), .QN(n447) );
  NAND2X1 U469 ( .IN1(n389), .IN2(mul_frac_out[37]), .QN(n451) );
  NAND2X1 U470 ( .IN1(n389), .IN2(mul_frac_out[38]), .QN(n455) );
  NAND2X1 U471 ( .IN1(n389), .IN2(mul_frac_out[39]), .QN(n459) );
  NAND2X1 U472 ( .IN1(n389), .IN2(mul_frac_out[40]), .QN(n463) );
  NAND2X1 U473 ( .IN1(n389), .IN2(mul_frac_out[41]), .QN(n467) );
  NAND2X1 U474 ( .IN1(n389), .IN2(mul_frac_out[42]), .QN(n471) );
  NAND2X1 U475 ( .IN1(n389), .IN2(mul_frac_out[43]), .QN(n475) );
  NAND2X1 U476 ( .IN1(n389), .IN2(mul_frac_out[44]), .QN(n479) );
  NAND2X1 U477 ( .IN1(n389), .IN2(mul_frac_out[45]), .QN(n483) );
  NAND2X1 U478 ( .IN1(n389), .IN2(mul_frac_out[46]), .QN(n487) );
  NAND2X1 U479 ( .IN1(n389), .IN2(mul_frac_out[47]), .QN(n491) );
  NAND2X1 U480 ( .IN1(n389), .IN2(mul_frac_out[48]), .QN(n495) );
  NAND2X1 U481 ( .IN1(n389), .IN2(mul_frac_out[49]), .QN(n499) );
  NAND2X1 U482 ( .IN1(n389), .IN2(mul_frac_out[50]), .QN(n503) );
  NAND2X1 U483 ( .IN1(n389), .IN2(mul_frac_out[51]), .QN(n507) );
  NAND2X1 U484 ( .IN1(n389), .IN2(mul_exp_out[0]), .QN(n511) );
  NAND2X1 U485 ( .IN1(n389), .IN2(mul_exp_out[1]), .QN(n515) );
  NAND2X1 U486 ( .IN1(n389), .IN2(mul_exp_out[2]), .QN(n519) );
  NAND2X1 U487 ( .IN1(n389), .IN2(mul_exp_out[3]), .QN(n523) );
  NAND2X1 U488 ( .IN1(n389), .IN2(mul_exp_out[4]), .QN(n527) );
  NAND2X1 U489 ( .IN1(n389), .IN2(mul_exp_out[5]), .QN(n531) );
  NAND2X1 U490 ( .IN1(n389), .IN2(mul_exp_out[6]), .QN(n535) );
  NAND2X1 U491 ( .IN1(n389), .IN2(mul_exp_out[7]), .QN(n539) );
  NAND2X1 U492 ( .IN1(n389), .IN2(mul_exp_out[8]), .QN(n543) );
  NAND2X1 U493 ( .IN1(n389), .IN2(mul_exp_out[9]), .QN(n547) );
  NAND2X1 U494 ( .IN1(n389), .IN2(mul_exp_out[10]), .QN(n551) );
  NAND2X1 U495 ( .IN1(n559), .IN2(m6stg_fmul_dbl_dst), .QN(n556) );
  AND2X1 U496 ( .IN1(grst_l), .IN2(n101), .Q(\fpu_out_ctl/dffrl_out_ctl/N4 )
         );
  AO222X1 U497 ( .IN1(\fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN2(m6stg_id_in[9]), 
        .IN3(n398), .IN4(div_id_out_in[9]), .IN5(\fpu_out_ctl/i_dest_rdy/N3 ), 
        .IN6(add_id_out_in[9]), .Q(\fpu_out_ctl/i_fp_cpx_req_cq/N10 ) );
  AO222X1 U498 ( .IN1(\fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN2(m6stg_id_in[2]), 
        .IN3(\fpu_out_ctl/i_dest_rdy/N3 ), .IN4(add_id_out_in[2]), .IN5(
        div_id_out_in[2]), .IN6(n398), .Q(\fpu_out_ctl/i_fp_cpx_req_cq/N3 ) );
  AO222X1 U499 ( .IN1(\fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN2(m6stg_id_in[3]), 
        .IN3(\fpu_out_ctl/i_dest_rdy/N3 ), .IN4(add_id_out_in[3]), .IN5(
        div_id_out_in[3]), .IN6(n398), .Q(\fpu_out_ctl/i_fp_cpx_req_cq/N4 ) );
  AO222X1 U500 ( .IN1(\fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN2(m6stg_id_in[4]), 
        .IN3(\fpu_out_ctl/i_dest_rdy/N3 ), .IN4(add_id_out_in[4]), .IN5(
        div_id_out_in[4]), .IN6(n398), .Q(\fpu_out_ctl/i_fp_cpx_req_cq/N5 ) );
  AO222X1 U501 ( .IN1(\fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN2(m6stg_id_in[5]), 
        .IN3(\fpu_out_ctl/i_dest_rdy/N3 ), .IN4(add_id_out_in[5]), .IN5(
        div_id_out_in[5]), .IN6(n398), .Q(\fpu_out_ctl/i_fp_cpx_req_cq/N6 ) );
  AO222X1 U502 ( .IN1(\fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN2(m6stg_id_in[6]), 
        .IN3(\fpu_out_ctl/i_dest_rdy/N3 ), .IN4(add_id_out_in[6]), .IN5(
        div_id_out_in[6]), .IN6(n398), .Q(\fpu_out_ctl/i_fp_cpx_req_cq/N7 ) );
  AO222X1 U503 ( .IN1(\fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN2(m6stg_id_in[7]), 
        .IN3(\fpu_out_ctl/i_dest_rdy/N3 ), .IN4(add_id_out_in[7]), .IN5(
        div_id_out_in[7]), .IN6(n398), .Q(\fpu_out_ctl/i_fp_cpx_req_cq/N8 ) );
  AO222X1 U504 ( .IN1(\fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN2(m6stg_id_in[8]), 
        .IN3(\fpu_out_ctl/i_dest_rdy/N3 ), .IN4(add_id_out_in[8]), .IN5(
        div_id_out_in[8]), .IN6(n398), .Q(\fpu_out_ctl/i_fp_cpx_req_cq/N9 ) );
  AO222X1 U505 ( .IN1(\fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN2(m6stg_id_in[0]), 
        .IN3(\fpu_out_ctl/i_dest_rdy/N3 ), .IN4(add_id_out_in[0]), .IN5(
        div_id_out_in[0]), .IN6(n398), .Q(\fpu_out_ctl/i_req_thread/N3 ) );
  AO222X1 U506 ( .IN1(\fpu_out_ctl/i_mul_dest_rdy/N3 ), .IN2(m6stg_id_in[1]), 
        .IN3(\fpu_out_ctl/i_dest_rdy/N3 ), .IN4(add_id_out_in[1]), .IN5(
        div_id_out_in[1]), .IN6(n398), .Q(\fpu_out_ctl/i_req_thread/N4 ) );
  NAND4X0 U507 ( .IN1(n402), .IN2(n401), .IN3(n400), .IN4(n399), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N18 ) );
  NAND4X0 U508 ( .IN1(n406), .IN2(n405), .IN3(n404), .IN4(n403), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N19 ) );
  NAND4X0 U509 ( .IN1(n410), .IN2(n409), .IN3(n408), .IN4(n407), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N20 ) );
  NAND4X0 U510 ( .IN1(n414), .IN2(n413), .IN3(n412), .IN4(n411), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N21 ) );
  NAND4X0 U511 ( .IN1(n418), .IN2(n417), .IN3(n416), .IN4(n415), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N22 ) );
  NAND4X0 U512 ( .IN1(n422), .IN2(n421), .IN3(n420), .IN4(n419), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N31 ) );
  NAND4X0 U513 ( .IN1(n426), .IN2(n425), .IN3(n424), .IN4(n423), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N32 ) );
  NAND4X0 U514 ( .IN1(n430), .IN2(n429), .IN3(n428), .IN4(n427), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N33 ) );
  AOI22X1 U515 ( .IN1(n390), .IN2(add_frac_out[40]), .IN3(n394), .IN4(
        div_frac_out[29]), .QN(n434) );
  AOI22X1 U516 ( .IN1(n392), .IN2(add_frac_out[43]), .IN3(n395), .IN4(
        add_frac_out[32]), .QN(n433) );
  AOI22X1 U517 ( .IN1(n391), .IN2(div_frac_out[32]), .IN3(n397), .IN4(
        mul_frac_out[29]), .QN(n432) );
  NAND4X0 U518 ( .IN1(n434), .IN2(n433), .IN3(n432), .IN4(n431), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N35 ) );
  AOI22X1 U519 ( .IN1(n390), .IN2(add_frac_out[41]), .IN3(n394), .IN4(
        div_frac_out[30]), .QN(n438) );
  AOI22X1 U520 ( .IN1(n392), .IN2(add_frac_out[44]), .IN3(n395), .IN4(
        add_frac_out[33]), .QN(n437) );
  AOI22X1 U521 ( .IN1(n391), .IN2(div_frac_out[33]), .IN3(n397), .IN4(
        mul_frac_out[30]), .QN(n436) );
  NAND4X0 U522 ( .IN1(n438), .IN2(n437), .IN3(n436), .IN4(n435), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N36 ) );
  AOI22X1 U523 ( .IN1(n390), .IN2(add_frac_out[42]), .IN3(n394), .IN4(
        div_frac_out[31]), .QN(n442) );
  AOI22X1 U524 ( .IN1(n392), .IN2(add_frac_out[45]), .IN3(n395), .IN4(
        add_frac_out[34]), .QN(n441) );
  AOI22X1 U525 ( .IN1(n391), .IN2(div_frac_out[34]), .IN3(n397), .IN4(
        mul_frac_out[31]), .QN(n440) );
  NAND4X0 U526 ( .IN1(n442), .IN2(n441), .IN3(n440), .IN4(n439), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N37 ) );
  AOI22X1 U527 ( .IN1(n390), .IN2(add_frac_out[43]), .IN3(n394), .IN4(
        div_frac_out[32]), .QN(n446) );
  AOI22X1 U528 ( .IN1(n392), .IN2(add_frac_out[46]), .IN3(n395), .IN4(
        add_frac_out[35]), .QN(n445) );
  AOI22X1 U529 ( .IN1(mul_frac_out[32]), .IN2(n397), .IN3(n391), .IN4(
        div_frac_out[35]), .QN(n444) );
  NAND4X0 U530 ( .IN1(n446), .IN2(n445), .IN3(n444), .IN4(n443), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N38 ) );
  AOI22X1 U531 ( .IN1(n390), .IN2(add_frac_out[44]), .IN3(n394), .IN4(
        div_frac_out[33]), .QN(n450) );
  AOI22X1 U532 ( .IN1(n392), .IN2(add_frac_out[47]), .IN3(n395), .IN4(
        add_frac_out[36]), .QN(n449) );
  AOI22X1 U533 ( .IN1(n391), .IN2(div_frac_out[36]), .IN3(n397), .IN4(
        mul_frac_out[33]), .QN(n448) );
  NAND4X0 U534 ( .IN1(n450), .IN2(n449), .IN3(n448), .IN4(n447), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N39 ) );
  AOI22X1 U535 ( .IN1(n390), .IN2(add_frac_out[45]), .IN3(n394), .IN4(
        div_frac_out[34]), .QN(n454) );
  AOI22X1 U536 ( .IN1(n392), .IN2(add_frac_out[48]), .IN3(n395), .IN4(
        add_frac_out[37]), .QN(n453) );
  AOI22X1 U537 ( .IN1(n391), .IN2(div_frac_out[37]), .IN3(n397), .IN4(
        mul_frac_out[34]), .QN(n452) );
  NAND4X0 U538 ( .IN1(n454), .IN2(n453), .IN3(n452), .IN4(n451), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N40 ) );
  AOI22X1 U539 ( .IN1(n390), .IN2(add_frac_out[46]), .IN3(n394), .IN4(
        div_frac_out[35]), .QN(n458) );
  AOI22X1 U540 ( .IN1(n392), .IN2(add_frac_out[49]), .IN3(n395), .IN4(
        add_frac_out[38]), .QN(n457) );
  AOI22X1 U541 ( .IN1(n391), .IN2(div_frac_out[38]), .IN3(n397), .IN4(
        mul_frac_out[35]), .QN(n456) );
  NAND4X0 U542 ( .IN1(n458), .IN2(n457), .IN3(n456), .IN4(n455), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N41 ) );
  AOI22X1 U543 ( .IN1(n390), .IN2(add_frac_out[47]), .IN3(n394), .IN4(
        div_frac_out[36]), .QN(n462) );
  AOI22X1 U544 ( .IN1(n392), .IN2(add_frac_out[50]), .IN3(n395), .IN4(
        add_frac_out[39]), .QN(n461) );
  AOI22X1 U545 ( .IN1(n391), .IN2(div_frac_out[39]), .IN3(n397), .IN4(
        mul_frac_out[36]), .QN(n460) );
  NAND4X0 U546 ( .IN1(n462), .IN2(n461), .IN3(n460), .IN4(n459), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N42 ) );
  AOI22X1 U547 ( .IN1(n390), .IN2(add_frac_out[48]), .IN3(n394), .IN4(
        div_frac_out[37]), .QN(n466) );
  AOI22X1 U548 ( .IN1(add_frac_out[40]), .IN2(n395), .IN3(n392), .IN4(
        add_frac_out[51]), .QN(n465) );
  AOI22X1 U549 ( .IN1(n391), .IN2(div_frac_out[40]), .IN3(n397), .IN4(
        mul_frac_out[37]), .QN(n464) );
  NAND4X0 U550 ( .IN1(n466), .IN2(n465), .IN3(n464), .IN4(n463), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N43 ) );
  AOI22X1 U551 ( .IN1(n390), .IN2(add_frac_out[49]), .IN3(n394), .IN4(
        div_frac_out[38]), .QN(n470) );
  AOI22X1 U552 ( .IN1(n392), .IN2(add_frac_out[52]), .IN3(n395), .IN4(
        add_frac_out[41]), .QN(n469) );
  AOI22X1 U553 ( .IN1(n391), .IN2(div_frac_out[41]), .IN3(n397), .IN4(
        mul_frac_out[38]), .QN(n468) );
  NAND4X0 U554 ( .IN1(n470), .IN2(n469), .IN3(n468), .IN4(n467), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N44 ) );
  AOI22X1 U555 ( .IN1(n390), .IN2(add_frac_out[50]), .IN3(n394), .IN4(
        div_frac_out[39]), .QN(n474) );
  AOI22X1 U556 ( .IN1(n392), .IN2(add_frac_out[53]), .IN3(n395), .IN4(
        add_frac_out[42]), .QN(n473) );
  AOI22X1 U557 ( .IN1(n391), .IN2(div_frac_out[42]), .IN3(n397), .IN4(
        mul_frac_out[39]), .QN(n472) );
  NAND4X0 U558 ( .IN1(n474), .IN2(n473), .IN3(n472), .IN4(n471), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N45 ) );
  AOI22X1 U559 ( .IN1(n390), .IN2(add_frac_out[51]), .IN3(n394), .IN4(
        div_frac_out[40]), .QN(n478) );
  AOI22X1 U560 ( .IN1(n392), .IN2(add_frac_out[54]), .IN3(add_frac_out[43]), 
        .IN4(n395), .QN(n477) );
  AOI22X1 U561 ( .IN1(n391), .IN2(div_frac_out[43]), .IN3(n397), .IN4(
        mul_frac_out[40]), .QN(n476) );
  NAND4X0 U562 ( .IN1(n478), .IN2(n477), .IN3(n476), .IN4(n475), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N46 ) );
  AOI22X1 U563 ( .IN1(n390), .IN2(add_frac_out[52]), .IN3(n394), .IN4(
        div_frac_out[41]), .QN(n482) );
  AOI22X1 U564 ( .IN1(n392), .IN2(add_frac_out[55]), .IN3(n395), .IN4(
        add_frac_out[44]), .QN(n481) );
  AOI22X1 U565 ( .IN1(n391), .IN2(div_frac_out[44]), .IN3(n397), .IN4(
        mul_frac_out[41]), .QN(n480) );
  NAND4X0 U566 ( .IN1(n482), .IN2(n481), .IN3(n480), .IN4(n479), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N47 ) );
  AOI22X1 U567 ( .IN1(n390), .IN2(add_frac_out[53]), .IN3(n394), .IN4(
        div_frac_out[42]), .QN(n486) );
  AOI22X1 U568 ( .IN1(n392), .IN2(add_frac_out[56]), .IN3(n395), .IN4(
        add_frac_out[45]), .QN(n485) );
  AOI22X1 U569 ( .IN1(n391), .IN2(div_frac_out[45]), .IN3(n397), .IN4(
        mul_frac_out[42]), .QN(n484) );
  NAND4X0 U570 ( .IN1(n486), .IN2(n485), .IN3(n484), .IN4(n483), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N48 ) );
  AOI22X1 U571 ( .IN1(n390), .IN2(add_frac_out[54]), .IN3(n394), .IN4(
        div_frac_out[43]), .QN(n490) );
  AOI22X1 U572 ( .IN1(n392), .IN2(add_frac_out[57]), .IN3(n395), .IN4(
        add_frac_out[46]), .QN(n489) );
  AOI22X1 U573 ( .IN1(n391), .IN2(div_frac_out[46]), .IN3(n397), .IN4(
        mul_frac_out[43]), .QN(n488) );
  NAND4X0 U574 ( .IN1(n490), .IN2(n489), .IN3(n488), .IN4(n487), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N49 ) );
  AOI22X1 U575 ( .IN1(n390), .IN2(add_frac_out[55]), .IN3(n394), .IN4(
        div_frac_out[44]), .QN(n494) );
  AOI22X1 U576 ( .IN1(n392), .IN2(add_frac_out[58]), .IN3(n395), .IN4(
        add_frac_out[47]), .QN(n493) );
  AOI22X1 U577 ( .IN1(n391), .IN2(div_frac_out[47]), .IN3(n397), .IN4(
        mul_frac_out[44]), .QN(n492) );
  NAND4X0 U578 ( .IN1(n494), .IN2(n493), .IN3(n492), .IN4(n491), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N50 ) );
  AOI22X1 U579 ( .IN1(n390), .IN2(add_frac_out[56]), .IN3(n394), .IN4(
        div_frac_out[45]), .QN(n498) );
  AOI22X1 U580 ( .IN1(n392), .IN2(add_frac_out[59]), .IN3(n395), .IN4(
        add_frac_out[48]), .QN(n497) );
  AOI22X1 U581 ( .IN1(n391), .IN2(div_frac_out[48]), .IN3(n397), .IN4(
        mul_frac_out[45]), .QN(n496) );
  NAND4X0 U582 ( .IN1(n498), .IN2(n497), .IN3(n496), .IN4(n495), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N51 ) );
  AOI22X1 U583 ( .IN1(n390), .IN2(add_frac_out[57]), .IN3(n394), .IN4(
        div_frac_out[46]), .QN(n502) );
  AOI22X1 U584 ( .IN1(n392), .IN2(add_frac_out[60]), .IN3(n395), .IN4(
        add_frac_out[49]), .QN(n501) );
  AOI22X1 U585 ( .IN1(n391), .IN2(div_frac_out[49]), .IN3(n397), .IN4(
        mul_frac_out[46]), .QN(n500) );
  NAND4X0 U586 ( .IN1(n502), .IN2(n501), .IN3(n500), .IN4(n499), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N52 ) );
  AOI22X1 U587 ( .IN1(n390), .IN2(add_frac_out[58]), .IN3(n394), .IN4(
        div_frac_out[47]), .QN(n506) );
  AOI22X1 U588 ( .IN1(n392), .IN2(add_frac_out[61]), .IN3(n395), .IN4(
        add_frac_out[50]), .QN(n505) );
  AOI22X1 U589 ( .IN1(n391), .IN2(div_frac_out[50]), .IN3(n397), .IN4(
        mul_frac_out[47]), .QN(n504) );
  NAND4X0 U590 ( .IN1(n506), .IN2(n505), .IN3(n504), .IN4(n503), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N53 ) );
  AOI22X1 U591 ( .IN1(n390), .IN2(add_frac_out[59]), .IN3(n394), .IN4(
        div_frac_out[48]), .QN(n510) );
  AOI22X1 U592 ( .IN1(n392), .IN2(add_frac_out[62]), .IN3(n395), .IN4(
        add_frac_out[51]), .QN(n509) );
  AOI22X1 U593 ( .IN1(n391), .IN2(div_frac_out[51]), .IN3(n397), .IN4(
        mul_frac_out[48]), .QN(n508) );
  NAND4X0 U594 ( .IN1(n510), .IN2(n509), .IN3(n508), .IN4(n507), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N54 ) );
  AOI22X1 U595 ( .IN1(n390), .IN2(add_frac_out[60]), .IN3(n394), .IN4(
        div_frac_out[49]), .QN(n514) );
  AOI22X1 U596 ( .IN1(n392), .IN2(add_exp_out[0]), .IN3(n395), .IN4(
        add_frac_out[52]), .QN(n513) );
  AOI22X1 U597 ( .IN1(n391), .IN2(div_exp_out[0]), .IN3(n397), .IN4(
        mul_frac_out[49]), .QN(n512) );
  NAND4X0 U598 ( .IN1(n514), .IN2(n513), .IN3(n512), .IN4(n511), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N55 ) );
  AOI22X1 U599 ( .IN1(n390), .IN2(add_frac_out[61]), .IN3(n394), .IN4(
        div_frac_out[50]), .QN(n518) );
  AOI22X1 U600 ( .IN1(n392), .IN2(add_exp_out[1]), .IN3(n395), .IN4(
        add_frac_out[53]), .QN(n517) );
  AOI22X1 U601 ( .IN1(n391), .IN2(div_exp_out[1]), .IN3(n397), .IN4(
        mul_frac_out[50]), .QN(n516) );
  NAND4X0 U602 ( .IN1(n518), .IN2(n517), .IN3(n516), .IN4(n515), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N56 ) );
  AOI22X1 U603 ( .IN1(n390), .IN2(add_frac_out[62]), .IN3(n394), .IN4(
        div_frac_out[51]), .QN(n522) );
  AOI22X1 U604 ( .IN1(n392), .IN2(add_exp_out[2]), .IN3(n395), .IN4(
        add_frac_out[54]), .QN(n521) );
  AOI22X1 U605 ( .IN1(n391), .IN2(div_exp_out[2]), .IN3(n397), .IN4(
        mul_frac_out[51]), .QN(n520) );
  NAND4X0 U606 ( .IN1(n522), .IN2(n521), .IN3(n520), .IN4(n519), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N57 ) );
  AOI22X1 U607 ( .IN1(n390), .IN2(add_exp_out[0]), .IN3(n394), .IN4(
        div_exp_out[0]), .QN(n526) );
  AOI22X1 U608 ( .IN1(n392), .IN2(add_exp_out[3]), .IN3(n395), .IN4(
        add_frac_out[55]), .QN(n525) );
  AOI22X1 U609 ( .IN1(n391), .IN2(div_exp_out[3]), .IN3(n397), .IN4(
        mul_exp_out[0]), .QN(n524) );
  NAND4X0 U610 ( .IN1(n526), .IN2(n525), .IN3(n524), .IN4(n523), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N58 ) );
  AOI22X1 U611 ( .IN1(n390), .IN2(add_exp_out[1]), .IN3(n394), .IN4(
        div_exp_out[1]), .QN(n530) );
  AOI22X1 U612 ( .IN1(n392), .IN2(add_exp_out[4]), .IN3(n395), .IN4(
        add_frac_out[56]), .QN(n529) );
  AOI22X1 U613 ( .IN1(n391), .IN2(div_exp_out[4]), .IN3(n397), .IN4(
        mul_exp_out[1]), .QN(n528) );
  NAND4X0 U614 ( .IN1(n530), .IN2(n529), .IN3(n528), .IN4(n527), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N59 ) );
  AOI22X1 U615 ( .IN1(n390), .IN2(add_exp_out[2]), .IN3(n394), .IN4(
        div_exp_out[2]), .QN(n534) );
  AOI22X1 U616 ( .IN1(n392), .IN2(add_exp_out[5]), .IN3(n395), .IN4(
        add_frac_out[57]), .QN(n533) );
  AOI22X1 U617 ( .IN1(n391), .IN2(div_exp_out[5]), .IN3(n397), .IN4(
        mul_exp_out[2]), .QN(n532) );
  NAND4X0 U618 ( .IN1(n534), .IN2(n533), .IN3(n532), .IN4(n531), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N60 ) );
  AOI22X1 U619 ( .IN1(n390), .IN2(add_exp_out[3]), .IN3(n394), .IN4(
        div_exp_out[3]), .QN(n538) );
  AOI22X1 U620 ( .IN1(n392), .IN2(add_exp_out[6]), .IN3(n395), .IN4(
        add_frac_out[58]), .QN(n537) );
  AOI22X1 U621 ( .IN1(n391), .IN2(div_exp_out[6]), .IN3(n397), .IN4(
        mul_exp_out[3]), .QN(n536) );
  NAND4X0 U622 ( .IN1(n538), .IN2(n537), .IN3(n536), .IN4(n535), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N61 ) );
  AOI22X1 U623 ( .IN1(n390), .IN2(add_exp_out[4]), .IN3(n394), .IN4(
        div_exp_out[4]), .QN(n542) );
  AOI22X1 U624 ( .IN1(n392), .IN2(add_exp_out[7]), .IN3(n395), .IN4(
        add_frac_out[59]), .QN(n541) );
  AOI22X1 U625 ( .IN1(n391), .IN2(div_exp_out[7]), .IN3(n397), .IN4(
        mul_exp_out[4]), .QN(n540) );
  NAND4X0 U626 ( .IN1(n542), .IN2(n541), .IN3(n540), .IN4(n539), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N62 ) );
  AOI22X1 U627 ( .IN1(n390), .IN2(add_exp_out[5]), .IN3(n394), .IN4(
        div_exp_out[5]), .QN(n546) );
  AOI22X1 U628 ( .IN1(n392), .IN2(add_exp_out[8]), .IN3(n395), .IN4(
        add_frac_out[60]), .QN(n545) );
  AOI22X1 U629 ( .IN1(n391), .IN2(div_exp_out[8]), .IN3(n397), .IN4(
        mul_exp_out[5]), .QN(n544) );
  NAND4X0 U630 ( .IN1(n546), .IN2(n545), .IN3(n544), .IN4(n543), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N63 ) );
  AOI22X1 U631 ( .IN1(n390), .IN2(add_exp_out[6]), .IN3(n394), .IN4(
        div_exp_out[6]), .QN(n550) );
  AOI22X1 U632 ( .IN1(n392), .IN2(add_exp_out[9]), .IN3(n395), .IN4(
        add_frac_out[61]), .QN(n549) );
  AOI22X1 U633 ( .IN1(n391), .IN2(div_exp_out[9]), .IN3(n397), .IN4(
        mul_exp_out[6]), .QN(n548) );
  NAND4X0 U634 ( .IN1(n550), .IN2(n549), .IN3(n548), .IN4(n547), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N64 ) );
  AOI22X1 U635 ( .IN1(n390), .IN2(add_exp_out[7]), .IN3(n394), .IN4(
        div_exp_out[7]), .QN(n554) );
  AOI22X1 U636 ( .IN1(n392), .IN2(add_exp_out[10]), .IN3(n395), .IN4(
        add_frac_out[62]), .QN(n553) );
  AOI22X1 U637 ( .IN1(n391), .IN2(div_exp_out[10]), .IN3(n397), .IN4(
        mul_exp_out[7]), .QN(n552) );
  NAND4X0 U638 ( .IN1(n554), .IN2(n553), .IN3(n552), .IN4(n551), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N65 ) );
  AND2X1 U639 ( .IN1(n557), .IN2(add_fcc_out[0]), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N68 ) );
  AND2X1 U640 ( .IN1(n557), .IN2(add_fcc_out[1]), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N69 ) );
  AND2X1 U641 ( .IN1(n557), .IN2(add_cc_out[0]), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N70 ) );
  AND2X1 U642 ( .IN1(n557), .IN2(add_cc_out[1]), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N71 ) );
  AND2X1 U643 ( .IN1(n557), .IN2(a6stg_fcmpop), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N72 ) );
  AO222X1 U644 ( .IN1(n559), .IN2(mul_exc_out[0]), .IN3(n558), .IN4(
        div_exc_out[0]), .IN5(add_exc_out[0]), .IN6(n557), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N75 ) );
  AO222X1 U645 ( .IN1(n559), .IN2(mul_exc_out[1]), .IN3(n558), .IN4(
        div_exc_out[1]), .IN5(add_exc_out[1]), .IN6(n557), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N76 ) );
  AO222X1 U646 ( .IN1(n559), .IN2(mul_exc_out[2]), .IN3(n558), .IN4(
        div_exc_out[2]), .IN5(add_exc_out[2]), .IN6(n557), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N77 ) );
  AO222X1 U647 ( .IN1(n559), .IN2(mul_exc_out[3]), .IN3(n558), .IN4(
        div_exc_out[3]), .IN5(add_exc_out[3]), .IN6(n557), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N78 ) );
  AO222X1 U648 ( .IN1(n559), .IN2(mul_exc_out[4]), .IN3(n558), .IN4(
        div_exc_out[4]), .IN5(add_exc_out[4]), .IN6(n557), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_76_0/N79 ) );
  NAND3X0 U649 ( .IN1(n562), .IN2(n561), .IN3(n560), .QN(
        \fpu_out_dp/i_fp_cpx_data_ca_84_77/N9 ) );
  AND2X1 U650 ( .IN1(req_thread[0]), .IN2(
        \fpu_out_dp/i_fp_cpx_data_ca_84_77/N9 ), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_84_77/N3 ) );
  AND2X1 U651 ( .IN1(req_thread[1]), .IN2(
        \fpu_out_dp/i_fp_cpx_data_ca_84_77/N9 ), .Q(
        \fpu_out_dp/i_fp_cpx_data_ca_84_77/N4 ) );
endmodule

