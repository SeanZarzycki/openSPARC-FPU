
module fpu_in ( pcx_fpio_data_rdy_px2, pcx_fpio_data_px2, a1stg_step, 
        m1stg_step, d1stg_step, add_pipe_active, mul_pipe_active, 
        div_pipe_active, inq_dout, sehold, arst_l, grst_l, rclk, fadd_clken_l, 
        fmul_clken_l, fdiv_clken_l, inq_add, inq_mul, inq_div, inq_id, 
        inq_rnd_mode, inq_fcc, inq_op, inq_in1_exp_neq_ffs, inq_in1_exp_eq_0, 
        inq_in1_53_0_neq_0, inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in1, 
        inq_in2_exp_neq_ffs, inq_in2_exp_eq_0, inq_in2_53_0_neq_0, 
        inq_in2_50_0_neq_0, inq_in2_53_32_neq_0, inq_in2, fp_id_in, 
        fp_rnd_mode_in, fp_fcc_in, fp_op_in, fp_src1_in, fp_src2_in, 
        inq_rdaddr, inq_wraddr, inq_read_en, inq_we, se, si, so );
  input [123:0] pcx_fpio_data_px2;
  input [154:0] inq_dout;
  output [4:0] inq_id;
  output [1:0] inq_rnd_mode;
  output [1:0] inq_fcc;
  output [7:0] inq_op;
  output [63:0] inq_in1;
  output [63:0] inq_in2;
  output [4:0] fp_id_in;
  output [1:0] fp_rnd_mode_in;
  output [1:0] fp_fcc_in;
  output [7:0] fp_op_in;
  output [68:0] fp_src1_in;
  output [68:0] fp_src2_in;
  output [3:0] inq_rdaddr;
  output [3:0] inq_wraddr;
  input pcx_fpio_data_rdy_px2, a1stg_step, m1stg_step, d1stg_step,
         add_pipe_active, mul_pipe_active, div_pipe_active, sehold, arst_l,
         grst_l, rclk, se, si;
  output fadd_clken_l, fmul_clken_l, fdiv_clken_l, inq_add, inq_mul, inq_div,
         inq_in1_exp_neq_ffs, inq_in1_exp_eq_0, inq_in1_53_0_neq_0,
         inq_in1_50_0_neq_0, inq_in1_53_32_neq_0, inq_in2_exp_neq_ffs,
         inq_in2_exp_eq_0, inq_in2_53_0_neq_0, inq_in2_50_0_neq_0,
         inq_in2_53_32_neq_0, inq_read_en, inq_we, so;
  wire   fp_op_in_7in, \fpu_in_ctl/in_ctl_rst_l , \fpu_in_ctl/dffrl_in_ctl/N4 ,
         \fpu_in_ctl/i_inq_rdptr/N6 , \fpu_in_ctl/i_inq_div_rdptr/N6 ,
         \fpu_in_ctl/i_inq_div_rdptr/N5 , \fpu_in_ctl/i_inq_div_rdptr/N4 ,
         \fpu_in_ctl/i_inq_div_rdptr/N3 , \fpu_in_ctl/i_inq_rdaddr_del/N6 ,
         \fpu_in_ctl/i_valid_packet_dly/N7 , \fpu_in_ctl/i_inq_rdptr_dec/N10 ,
         \fpu_in_ctl/i_inq_rdptr_dec/N9 , \fpu_in_ctl/i_inq_rdptr_dec/N8 ,
         \fpu_in_ctl/i_inq_rdptr_dec/N7 , \fpu_in_ctl/i_inq_rdptr_dec/N6 ,
         \fpu_in_ctl/i_inq_rdptr_dec/N5 , \fpu_in_ctl/i_inq_rdptr_dec/N4 ,
         \fpu_in_ctl/i_inq_rdptr_dec/N3 , \fpu_in_ctl/i_inq_div_rdptr_dec/N10 ,
         \fpu_in_ctl/i_inq_div_rdptr_dec/N9 ,
         \fpu_in_ctl/i_inq_div_rdptr_dec/N8 ,
         \fpu_in_ctl/i_inq_div_rdptr_dec/N7 ,
         \fpu_in_ctl/i_inq_div_rdptr_dec/N6 ,
         \fpu_in_ctl/i_inq_div_rdptr_dec/N5 ,
         \fpu_in_ctl/i_inq_div_rdptr_dec/N4 ,
         \fpu_in_ctl/i_inq_rdaddr_del_dec/N18 ,
         \fpu_in_ctl/i_inq_rdaddr_del_dec/N17 ,
         \fpu_in_ctl/i_inq_rdaddr_del_dec/N16 ,
         \fpu_in_ctl/i_inq_rdaddr_del_dec/N15 ,
         \fpu_in_ctl/i_inq_rdaddr_del_dec/N14 ,
         \fpu_in_ctl/i_inq_rdaddr_del_dec/N13 ,
         \fpu_in_ctl/i_inq_rdaddr_del_dec/N12 , n4, n6, n8, n41, n111, n114,
         n121, n255, n256, n257, n322, n323, n325, n326, n328, n329, n331,
         n332, n334, n335, n337, n338, n340, n341, n343, n344, n346, n347,
         n348, n349, n350, n353, n356, n359, n362, n365, n368, n371, n374,
         n375, n376, n377, n418, \fpu_in_dp/n105 , \fpu_in_dp/n714 ,
         \fpu_in_dp/n713 , \fpu_in_dp/n712 , \fpu_in_dp/n711 ,
         \fpu_in_dp/n710 , \fpu_in_dp/n709 , \fpu_in_dp/n708 ,
         \fpu_in_dp/n707 , \fpu_in_dp/n706 , \fpu_in_dp/n705 ,
         \fpu_in_dp/n704 , \fpu_in_dp/n703 , \fpu_in_dp/n702 ,
         \fpu_in_dp/n701 , \fpu_in_dp/n700 , \fpu_in_dp/n699 ,
         \fpu_in_dp/n698 , \fpu_in_dp/n697 , \fpu_in_dp/n696 ,
         \fpu_in_dp/n695 , \fpu_in_dp/n694 , \fpu_in_dp/n693 ,
         \fpu_in_dp/n692 , \fpu_in_dp/n691 , \fpu_in_dp/n690 ,
         \fpu_in_dp/n689 , \fpu_in_dp/n688 , \fpu_in_dp/n687 ,
         \fpu_in_dp/n686 , \fpu_in_dp/n685 , \fpu_in_dp/n684 ,
         \fpu_in_dp/n683 , \fpu_in_dp/n682 , \fpu_in_dp/n681 ,
         \fpu_in_dp/n680 , \fpu_in_dp/n679 , \fpu_in_dp/n678 ,
         \fpu_in_dp/n677 , \fpu_in_dp/n676 , \fpu_in_dp/n675 ,
         \fpu_in_dp/n674 , \fpu_in_dp/n673 , \fpu_in_dp/n672 ,
         \fpu_in_dp/n671 , \fpu_in_dp/n670 , \fpu_in_dp/n669 ,
         \fpu_in_dp/n668 , \fpu_in_dp/n667 , \fpu_in_dp/n666 ,
         \fpu_in_dp/n665 , \fpu_in_dp/n664 , \fpu_in_dp/n663 ,
         \fpu_in_dp/n662 , \fpu_in_dp/n661 , \fpu_in_dp/n660 ,
         \fpu_in_dp/n659 , \fpu_in_dp/n658 , \fpu_in_dp/n657 ,
         \fpu_in_dp/n656 , \fpu_in_dp/n655 , \fpu_in_dp/n654 ,
         \fpu_in_dp/n653 , \fpu_in_dp/n652 , \fpu_in_dp/n651 ,
         \fpu_in_dp/n650 , \fpu_in_dp/n649 , \fpu_in_dp/n648 ,
         \fpu_in_dp/n647 , \fpu_in_dp/n646 , \fpu_in_dp/n473 ,
         \fpu_in_dp/n469 , \fpu_in_dp/n467 , \fpu_in_dp/n465 ,
         \fpu_in_dp/n463 , \fpu_in_dp/n461 , \fpu_in_dp/n458 ,
         \fpu_in_dp/n456 , \fpu_in_dp/n454 , \fpu_in_dp/n452 ,
         \fpu_in_dp/n450 , \fpu_in_dp/n448 , \fpu_in_dp/n445 ,
         \fpu_in_dp/n443 , \fpu_in_dp/n441 , \fpu_in_dp/n439 , \fpu_in_dp/n32 ,
         \fpu_in_dp/n31 , \fpu_in_dp/n29 , \fpu_in_dp/n27 , \fpu_in_dp/n25 ,
         \fpu_in_dp/n23 , \fpu_in_dp/n21 , \fpu_in_dp/n18 , \fpu_in_dp/n16 ,
         \fpu_in_dp/n14 , \fpu_in_dp/n12 , \fpu_in_dp/n10 , \fpu_in_dp/n8 ,
         \fpu_in_dp/n6 , \fpu_in_dp/n4 , \fpu_in_dp/n2 ,
         \fpu_in_dp/i_inq_din_d1/N72 , \fpu_in_dp/i_inq_din_d1/N73 ,
         \fpu_in_dp/i_inq_din_d1/N74 , \fpu_in_dp/i_inq_din_d1/N75 ,
         \fpu_in_dp/i_inq_din_d1/N76 , \fpu_in_dp/i_inq_din_d1/N77 ,
         \fpu_in_dp/i_inq_din_d1/N78 , \fpu_in_dp/i_inq_din_d1/N79 ,
         \fpu_in_dp/i_inq_din_d1/N80 , \fpu_in_dp/i_inq_din_d1/N81 ,
         \fpu_in_dp/i_inq_din_d1/N82 , \fpu_in_dp/i_inq_din_d1/N83 ,
         \fpu_in_dp/i_inq_din_d1/N84 , \fpu_in_dp/i_inq_din_d1/N85 ,
         \fpu_in_dp/i_inq_din_d1/N86 , \fpu_in_dp/i_inq_din_d1/N87 ,
         \fpu_in_dp/i_inq_din_d1/N88 , \fpu_in_dp/i_inq_din_d1/N89 ,
         \fpu_in_dp/i_inq_din_d1/N90 , \fpu_in_dp/i_inq_din_d1/N91 ,
         \fpu_in_dp/i_inq_din_d1/N92 , \fpu_in_dp/i_inq_din_d1/N93 ,
         \fpu_in_dp/i_inq_din_d1/N94 , \fpu_in_dp/i_inq_din_d1/N95 ,
         \fpu_in_dp/i_inq_din_d1/N96 , \fpu_in_dp/i_inq_din_d1/N97 ,
         \fpu_in_dp/i_inq_din_d1/N98 , \fpu_in_dp/i_inq_din_d1/N99 ,
         \fpu_in_dp/i_inq_din_d1/N100 , \fpu_in_dp/i_inq_din_d1/N101 ,
         \fpu_in_dp/i_inq_din_d1/N102 , \fpu_in_dp/i_inq_din_d1/N103 ,
         \fpu_in_dp/i_inq_din_d1/N104 , \fpu_in_dp/i_inq_din_d1/N105 ,
         \fpu_in_dp/i_inq_din_d1/N106 , \fpu_in_dp/i_inq_din_d1/N107 ,
         \fpu_in_dp/i_inq_din_d1/N108 , \fpu_in_dp/i_inq_din_d1/N109 ,
         \fpu_in_dp/i_inq_din_d1/N110 , \fpu_in_dp/i_inq_din_d1/N111 ,
         \fpu_in_dp/i_inq_din_d1/N112 , \fpu_in_dp/i_inq_din_d1/N113 ,
         \fpu_in_dp/i_inq_din_d1/N114 , \fpu_in_dp/i_inq_din_d1/N115 ,
         \fpu_in_dp/i_inq_din_d1/N116 , \fpu_in_dp/i_inq_din_d1/N117 ,
         \fpu_in_dp/i_inq_din_d1/N118 , \fpu_in_dp/i_inq_din_d1/N119 ,
         \fpu_in_dp/i_inq_din_d1/N120 , \fpu_in_dp/i_inq_din_d1/N121 ,
         \fpu_in_dp/i_inq_din_d1/N122 , \fpu_in_dp/i_inq_din_d1/N123 ,
         \fpu_in_dp/i_inq_din_d1/N124 , \fpu_in_dp/i_inq_din_d1/N125 ,
         \fpu_in_dp/i_inq_din_d1/N126 , \fpu_in_dp/i_inq_din_d1/N127 ,
         \fpu_in_dp/i_inq_din_d1/N128 , \fpu_in_dp/i_inq_din_d1/N129 ,
         \fpu_in_dp/i_inq_din_d1/N130 , \fpu_in_dp/i_inq_din_d1/N131 ,
         \fpu_in_dp/i_inq_din_d1/N132 , \fpu_in_dp/i_inq_din_d1/N133 ,
         \fpu_in_dp/i_inq_din_d1/N134 , \fpu_in_dp/i_inq_din_d1/N135 ,
         \fpu_in_dp/i_inq_din_d1/N136 , \fpu_in_dp/i_inq_din_d1/N138 ,
         \fpu_in_dp/i_inq_din_d1/N139 , \fpu_in_dp/i_inq_din_d1/N140 ,
         \fpu_in_dp/i_inq_din_d1/N141 , \fpu_in_dp/i_inq_din_d1/N148 , n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n911, n912, n913, n914,
         n916, n917, n1155, n1159, n1161, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1619,
         n1620, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988;
  assign fp_op_in[7] = fp_op_in_7in;
  assign so = 1'b0;

  DFFARX1 \fpu_in_ctl/dffrl_in_ctl/q_reg[0]  ( .D(\fpu_in_ctl/dffrl_in_ctl/N4 ), .CLK(rclk), .RSTB(arst_l), .Q(\fpu_in_ctl/in_ctl_rst_l ), .QN(n418) );
  DFFSSRX1 \fpu_in_ctl/i_fp_data_rdy/q_reg[0]  ( .D(n1848), .RSTB(
        pcx_fpio_data_rdy_px2), .SETB(1'b1), .CLK(rclk), .Q(n1571), .QN(n1679)
         );
  DFFSSRX1 \fpu_in_ctl/i_fp_vld_in/q_reg[0]  ( .D(pcx_fpio_data_px2[123]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n1570) );
  DFFSSRX1 \fpu_in_ctl/i_fp_type_in/q_reg[0]  ( .D(pcx_fpio_data_px2[118]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n1567) );
  DFFSSRX1 \fpu_in_ctl/i_fp_type_in/q_reg[1]  ( .D(pcx_fpio_data_px2[119]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n1572) );
  DFFSSRX1 \fpu_in_ctl/i_fp_type_in/q_reg[2]  ( .D(pcx_fpio_data_px2[120]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n1568) );
  DFFSSRX1 \fpu_in_ctl/i_fp_type_in/q_reg[3]  ( .D(pcx_fpio_data_px2[121]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .QN(n121) );
  DFFSSRX1 \fpu_in_ctl/i_fp_type_in/q_reg[4]  ( .D(pcx_fpio_data_px2[122]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n1569) );
  DFFX1 \fpu_in_ctl/i_valid_packet_dly/q_reg[0]  ( .D(
        \fpu_in_ctl/i_valid_packet_dly/N7 ), .CLK(rclk), .Q(n1544) );
  DFFSSRX1 \fpu_in_ctl/i_d1stg_step_dly/q_reg[0]  ( .D(d1stg_step), .RSTB(
        n1848), .SETB(1'b1), .CLK(rclk), .Q(n1549) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr_dec/q_reg[7]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N10 ), .CLK(rclk), .Q(n891) );
  DFFSSRX1 \fpu_in_ctl/i_inq_div_rdptr_dec/q_reg[0]  ( .D(
        \fpu_in_ctl/in_ctl_rst_l ), .RSTB(n1161), .SETB(n1850), .CLK(rclk), 
        .Q(n114), .QN(n917) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr_dec/q_reg[1]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N4 ), .CLK(rclk), .Q(n805) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr_dec/q_reg[2]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N5 ), .CLK(rclk), .Q(n885) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr_dec/q_reg[3]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N6 ), .CLK(rclk), .Q(n804) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr_dec/q_reg[4]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N7 ), .CLK(rclk), .Q(n884) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr_dec/q_reg[5]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N8 ), .CLK(rclk), .Q(n752) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr_dec/q_reg[6]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N9 ), .CLK(rclk), .Q(n806) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr/q_reg[0]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr/N3 ), .CLK(rclk), .Q(n813) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr/q_reg[2]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr/N5 ), .CLK(rclk), .Q(n1671), .QN(n1560) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr/q_reg[3]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr/N6 ), .CLK(rclk), .Q(n1677), .QN(n1562) );
  DFFX1 \fpu_in_ctl/i_inq_div_rdptr/q_reg[1]  ( .D(
        \fpu_in_ctl/i_inq_div_rdptr/N4 ), .CLK(rclk), .Q(n755) );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del/q_reg[1]  ( .D(n1850), .RSTB(
        inq_rdaddr[1]), .SETB(1'b1), .CLK(rclk), .QN(n111) );
  DFFX1 \fpu_in_ctl/i_inq_div_wrptr/q_reg[0]  ( .D(n377), .CLK(rclk), .Q(n1649), .QN(n889) );
  DFFX1 \fpu_in_ctl/i_inq_div_wrptr/q_reg[1]  ( .D(n376), .CLK(rclk), .Q(n754), 
        .QN(n1675) );
  DFFSSRX1 \fpu_in_ctl/i_inq_wraddr_del/q_reg[3]  ( .D(n1849), .RSTB(
        inq_wraddr[3]), .SETB(1'b1), .CLK(rclk), .Q(n1545) );
  DFFX1 \fpu_in_ctl/i_inq_div_wrptr/q_reg[2]  ( .D(n375), .CLK(rclk), .Q(n1651), .QN(n1561) );
  DFFX1 \fpu_in_ctl/i_inq_pipe12/q_reg[2]  ( .D(n362), .CLK(rclk), .Q(n1695)
         );
  DFFX1 \fpu_in_ctl/i_inq_pipe13/q_reg[2]  ( .D(n365), .CLK(rclk), .Q(n1669)
         );
  DFFX1 \fpu_in_ctl/i_inq_pipe14/q_reg[2]  ( .D(n368), .CLK(rclk), .Q(n1696)
         );
  DFFX1 \fpu_in_ctl/i_inq_pipe15/q_reg[2]  ( .D(n371), .CLK(rclk), .Q(n1557)
         );
  DFFX1 \fpu_in_ctl/i_inq_div_wrptr/q_reg[3]  ( .D(n374), .CLK(rclk), .Q(n1652), .QN(n1563) );
  DFFX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[15]  ( .D(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N18 ), .CLK(rclk), .Q(n1556) );
  DFFX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[14]  ( .D(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N17 ), .CLK(rclk), .Q(n1558) );
  DFFX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[13]  ( .D(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N16 ), .CLK(rclk), .Q(n1554) );
  DFFX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[12]  ( .D(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N15 ), .CLK(rclk), .Q(n1555) );
  DFFX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[11]  ( .D(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N14 ), .CLK(rclk), .Q(n1551) );
  DFFX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[10]  ( .D(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N13 ), .CLK(rclk), .Q(n1550) );
  DFFX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[9]  ( .D(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N12 ), .CLK(rclk), .Q(n1553) );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[8]  ( .D(n114), .RSTB(
        \fpu_in_ctl/in_ctl_rst_l ), .SETB(\fpu_in_ctl/i_inq_rdaddr_del/N6 ), 
        .CLK(rclk), .QN(n1552) );
  DFFSSRX1 \fpu_in_ctl/i_inq_div_rd/q_reg[0]  ( .D(n1849), .RSTB(inq_rdaddr[3]), .SETB(1'b1), .CLK(rclk), .QN(n1682) );
  DFFX1 \fpu_in_ctl/i_inq_pipe8/q_reg[2]  ( .D(n350), .CLK(rclk), .Q(n914) );
  DFFX1 \fpu_in_ctl/i_inq_pipe9/q_reg[2]  ( .D(n353), .CLK(rclk), .Q(n912) );
  DFFX1 \fpu_in_ctl/i_inq_pipe10/q_reg[2]  ( .D(n356), .CLK(rclk), .Q(n913) );
  DFFX1 \fpu_in_ctl/i_inq_pipe11/q_reg[2]  ( .D(n359), .CLK(rclk), .Q(n911) );
  DFFX1 \fpu_in_ctl/i_inq_wrptr/q_reg[0]  ( .D(n349), .CLK(rclk), .Q(n1670), 
        .QN(n807) );
  DFFSSRX1 \fpu_in_ctl/i_inq_wraddr_del/q_reg[0]  ( .D(n1849), .RSTB(
        inq_wraddr[0]), .SETB(1'b1), .CLK(rclk), .Q(n1546) );
  DFFX1 \fpu_in_ctl/i_inq_wrptr/q_reg[1]  ( .D(n348), .CLK(rclk), .Q(n1650), 
        .QN(n886) );
  DFFSSRX1 \fpu_in_ctl/i_inq_wraddr_del/q_reg[1]  ( .D(n1849), .RSTB(
        inq_wraddr[1]), .SETB(1'b1), .CLK(rclk), .Q(n1548) );
  DFFX1 \fpu_in_ctl/i_inq_wrptr/q_reg[2]  ( .D(n347), .CLK(rclk), .Q(n1673), 
        .QN(n812) );
  DFFSSRX1 \fpu_in_ctl/i_inq_wraddr_del/q_reg[2]  ( .D(n1850), .RSTB(
        inq_wraddr[2]), .SETB(1'b1), .CLK(rclk), .Q(n1547) );
  DFFX1 \fpu_in_ctl/i_inq_wrptr/q_reg[3]  ( .D(n346), .CLK(rclk), .Q(n1566) );
  DFFX1 \fpu_in_ctl/i_inq_pipe3/q_reg[1]  ( .D(n335), .CLK(rclk), .Q(n894) );
  DFFX1 \fpu_in_ctl/i_inq_pipe2/q_reg[1]  ( .D(n338), .CLK(rclk), .Q(n902) );
  DFFX1 \fpu_in_ctl/i_inq_pipe1/q_reg[1]  ( .D(n341), .CLK(rclk), .Q(n892) );
  DFFX1 \fpu_in_ctl/i_inq_pipe0/q_reg[1]  ( .D(n344), .CLK(rclk), .Q(n900) );
  DFFX1 \fpu_in_ctl/i_inq_pipe7/q_reg[1]  ( .D(n323), .CLK(rclk), .Q(n898) );
  DFFX1 \fpu_in_ctl/i_inq_pipe6/q_reg[1]  ( .D(n326), .CLK(rclk), .Q(n906) );
  DFFX1 \fpu_in_ctl/i_inq_pipe5/q_reg[1]  ( .D(n329), .CLK(rclk), .Q(n896) );
  DFFX1 \fpu_in_ctl/i_inq_pipe4/q_reg[1]  ( .D(n332), .CLK(rclk), .Q(n904) );
  DFFX1 \fpu_in_ctl/i_inq_pipe7/q_reg[0]  ( .D(n322), .CLK(rclk), .Q(n899) );
  DFFX1 \fpu_in_ctl/i_inq_pipe6/q_reg[0]  ( .D(n325), .CLK(rclk), .Q(n907) );
  DFFX1 \fpu_in_ctl/i_inq_pipe5/q_reg[0]  ( .D(n328), .CLK(rclk), .Q(n897) );
  DFFX1 \fpu_in_ctl/i_inq_pipe4/q_reg[0]  ( .D(n331), .CLK(rclk), .Q(n905) );
  DFFX1 \fpu_in_ctl/i_inq_pipe3/q_reg[0]  ( .D(n334), .CLK(rclk), .Q(n895) );
  DFFX1 \fpu_in_ctl/i_inq_pipe2/q_reg[0]  ( .D(n337), .CLK(rclk), .Q(n903) );
  DFFX1 \fpu_in_ctl/i_inq_pipe1/q_reg[0]  ( .D(n340), .CLK(rclk), .Q(n893) );
  DFFX1 \fpu_in_ctl/i_inq_pipe0/q_reg[0]  ( .D(n343), .CLK(rclk), .Q(n901) );
  DFFSSRX1 \fpu_in_ctl/i_inq_adda_dly/q_reg[0]  ( .D(inq_add), .RSTB(n1848), 
        .SETB(1'b1), .CLK(rclk), .QN(n41) );
  DFFX1 \fpu_in_ctl/i_inq_rdptr_dec/q_reg[7]  ( .D(
        \fpu_in_ctl/i_inq_rdptr_dec/N10 ), .CLK(rclk), .Q(n908) );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdptr_dec/q_reg[0]  ( .D(
        \fpu_in_ctl/in_ctl_rst_l ), .RSTB(n1155), .SETB(n1850), .CLK(rclk), 
        .QN(n916) );
  DFFX1 \fpu_in_ctl/i_inq_rdptr_dec/q_reg[1]  ( .D(
        \fpu_in_ctl/i_inq_rdptr_dec/N4 ), .CLK(rclk), .Q(n809) );
  DFFX1 \fpu_in_ctl/i_inq_rdptr_dec/q_reg[2]  ( .D(
        \fpu_in_ctl/i_inq_rdptr_dec/N5 ), .CLK(rclk), .Q(n888) );
  DFFX1 \fpu_in_ctl/i_inq_rdptr_dec/q_reg[3]  ( .D(
        \fpu_in_ctl/i_inq_rdptr_dec/N6 ), .CLK(rclk), .Q(n808) );
  DFFX1 \fpu_in_ctl/i_inq_rdptr_dec/q_reg[4]  ( .D(
        \fpu_in_ctl/i_inq_rdptr_dec/N7 ), .CLK(rclk), .Q(n887) );
  DFFX1 \fpu_in_ctl/i_inq_rdptr_dec/q_reg[5]  ( .D(
        \fpu_in_ctl/i_inq_rdptr_dec/N8 ), .CLK(rclk), .Q(n753) );
  DFFX1 \fpu_in_ctl/i_inq_rdptr_dec/q_reg[6]  ( .D(
        \fpu_in_ctl/i_inq_rdptr_dec/N9 ), .CLK(rclk), .Q(n810) );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[6]  ( .D(n1159), .RSTB(
        \fpu_in_ctl/i_inq_rdptr_dec/N9 ), .SETB(1'b1), .CLK(rclk), .Q(n1579)
         );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[5]  ( .D(n1159), .RSTB(
        \fpu_in_ctl/i_inq_rdptr_dec/N8 ), .SETB(1'b1), .CLK(rclk), .Q(n1580)
         );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[4]  ( .D(n1159), .RSTB(
        \fpu_in_ctl/i_inq_rdptr_dec/N7 ), .SETB(1'b1), .CLK(rclk), .Q(n1577)
         );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[3]  ( .D(n1159), .RSTB(
        \fpu_in_ctl/i_inq_rdptr_dec/N6 ), .SETB(1'b1), .CLK(rclk), .Q(n1578)
         );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[2]  ( .D(n1159), .RSTB(
        \fpu_in_ctl/i_inq_rdptr_dec/N5 ), .SETB(1'b1), .CLK(rclk), .Q(n1575)
         );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[1]  ( .D(n1159), .RSTB(
        \fpu_in_ctl/i_inq_rdptr_dec/N4 ), .SETB(1'b1), .CLK(rclk), .Q(n1576)
         );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[0]  ( .D(
        \fpu_in_ctl/i_inq_rdptr_dec/N3 ), .RSTB(n1159), .SETB(1'b1), .CLK(rclk), .Q(n1573) );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del_dec/q_reg[7]  ( .D(n1159), .RSTB(
        \fpu_in_ctl/i_inq_rdptr_dec/N10 ), .SETB(1'b1), .CLK(rclk), .Q(n1574)
         );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdptr/q_reg[0]  ( .D(n1850), .RSTB(n257), .SETB(
        1'b1), .CLK(rclk), .Q(n756) );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdptr/q_reg[1]  ( .D(n256), .RSTB(n1849), .SETB(
        1'b1), .CLK(rclk), .Q(n814), .QN(n1672) );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdptr/q_reg[2]  ( .D(n255), .RSTB(n1849), .SETB(
        1'b1), .CLK(rclk), .Q(n1564) );
  DFFX1 \fpu_in_ctl/i_inq_rdptr/q_reg[3]  ( .D(\fpu_in_ctl/i_inq_rdptr/N6 ), 
        .CLK(rclk), .Q(n1698), .QN(n1565) );
  DFFSSRX1 \fpu_in_ctl/i_inq_mula_dly/q_reg[0]  ( .D(inq_mul), .RSTB(n1848), 
        .SETB(1'b1), .CLK(rclk), .QN(n8) );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del/q_reg[2]  ( .D(n1849), .RSTB(
        inq_rdaddr[2]), .SETB(1'b1), .CLK(rclk), .QN(n6) );
  DFFSSRX1 \fpu_in_ctl/i_inq_rdaddr_del/q_reg[0]  ( .D(n1849), .RSTB(
        inq_rdaddr[0]), .SETB(1'b1), .CLK(rclk), .QN(n4) );
  DFFSSRX1 \fpu_in_ctl/i_inq_diva_dly/q_reg[0]  ( .D(inq_div), .RSTB(n1848), 
        .SETB(1'b1), .CLK(rclk), .Q(n890) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[154]  ( .D(fp_id_in[4]), .RSTB(n1849), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n2 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[153]  ( .D(fp_id_in[3]), .RSTB(n1850), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n4 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[152]  ( .D(fp_id_in[2]), .RSTB(n1849), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n6 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[151]  ( .D(fp_id_in[1]), .RSTB(n1849), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n8 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[150]  ( .D(fp_id_in[0]), .RSTB(n1850), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n10 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[149]  ( .D(fp_rnd_mode_in[1]), .RSTB(
        n1849), .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n12 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[148]  ( .D(fp_rnd_mode_in[0]), .RSTB(
        n1849), .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n14 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[147]  ( .D(fp_fcc_in[1]), .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n16 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[146]  ( .D(fp_fcc_in[0]), .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n18 ) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[145]  ( .D(\fpu_in_dp/i_inq_din_d1/N148 ), .CLK(rclk), .Q(n1837) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[144]  ( .D(fp_op_in[6]), .RSTB(n1849), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n21 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[143]  ( .D(fp_op_in[5]), .RSTB(n1849), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n23 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[142]  ( .D(fp_op_in[4]), .RSTB(n1850), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n25 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[141]  ( .D(fp_op_in[3]), .RSTB(n1849), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n27 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[140]  ( .D(fp_op_in[2]), .RSTB(n1849), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n29 ) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[139]  ( .D(n1849), .RSTB(fp_op_in[1]), 
        .SETB(1'b1), .CLK(rclk), .QN(\fpu_in_dp/n31 ) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[138]  ( .D(\fpu_in_dp/i_inq_din_d1/N141 ), .CLK(rclk), .QN(\fpu_in_dp/n32 ) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[137]  ( .D(\fpu_in_dp/i_inq_din_d1/N140 ), .CLK(rclk), .Q(n1836) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[136]  ( .D(\fpu_in_dp/i_inq_din_d1/N139 ), .CLK(rclk), .Q(n1835) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[135]  ( .D(\fpu_in_dp/i_inq_din_d1/N138 ), .CLK(rclk), .Q(n1833) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[134]  ( .D(n1850), .RSTB(
        fp_src1_in[65]), .SETB(1'b1), .CLK(rclk), .Q(n1699) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[133]  ( .D(\fpu_in_dp/i_inq_din_d1/N136 ), .CLK(rclk), .Q(n1834) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[132]  ( .D(\fpu_in_dp/i_inq_din_d1/N135 ), .CLK(rclk), .Q(n1828) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[131]  ( .D(\fpu_in_dp/i_inq_din_d1/N134 ), .CLK(rclk), .Q(n1827) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[130]  ( .D(\fpu_in_dp/i_inq_din_d1/N133 ), .CLK(rclk), .Q(n1826) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[129]  ( .D(\fpu_in_dp/i_inq_din_d1/N132 ), .CLK(rclk), .Q(n1825) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[128]  ( .D(\fpu_in_dp/i_inq_din_d1/N131 ), .CLK(rclk), .Q(n1823) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[127]  ( .D(\fpu_in_dp/i_inq_din_d1/N130 ), .CLK(rclk), .Q(n1822) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[126]  ( .D(\fpu_in_dp/i_inq_din_d1/N129 ), .CLK(rclk), .Q(n1821) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[125]  ( .D(\fpu_in_dp/i_inq_din_d1/N128 ), .CLK(rclk), .Q(n1820) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[124]  ( .D(\fpu_in_dp/i_inq_din_d1/N127 ), .CLK(rclk), .Q(n1819) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[123]  ( .D(\fpu_in_dp/i_inq_din_d1/N126 ), .CLK(rclk), .Q(n1818) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[122]  ( .D(\fpu_in_dp/i_inq_din_d1/N125 ), .CLK(rclk), .Q(n1817) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[121]  ( .D(\fpu_in_dp/i_inq_din_d1/N124 ), .CLK(rclk), .Q(n1816) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[120]  ( .D(\fpu_in_dp/i_inq_din_d1/N123 ), .CLK(rclk), .Q(n1815) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[119]  ( .D(\fpu_in_dp/i_inq_din_d1/N122 ), .CLK(rclk), .Q(n1814) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[118]  ( .D(\fpu_in_dp/i_inq_din_d1/N121 ), .CLK(rclk), .Q(n1812) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[117]  ( .D(\fpu_in_dp/i_inq_din_d1/N120 ), .CLK(rclk), .Q(n1811) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[116]  ( .D(\fpu_in_dp/i_inq_din_d1/N119 ), .CLK(rclk), .Q(n1810) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[115]  ( .D(\fpu_in_dp/i_inq_din_d1/N118 ), .CLK(rclk), .Q(n1809) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[114]  ( .D(\fpu_in_dp/i_inq_din_d1/N117 ), .CLK(rclk), .Q(n1808) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[113]  ( .D(\fpu_in_dp/i_inq_din_d1/N116 ), .CLK(rclk), .Q(n1807) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[112]  ( .D(\fpu_in_dp/i_inq_din_d1/N115 ), .CLK(rclk), .Q(n1806) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[111]  ( .D(\fpu_in_dp/i_inq_din_d1/N114 ), .CLK(rclk), .Q(n1805) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[110]  ( .D(\fpu_in_dp/i_inq_din_d1/N113 ), .CLK(rclk), .Q(n1804) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[109]  ( .D(\fpu_in_dp/i_inq_din_d1/N112 ), .CLK(rclk), .Q(n1803) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[108]  ( .D(\fpu_in_dp/i_inq_din_d1/N111 ), .CLK(rclk), .Q(n1801) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[107]  ( .D(\fpu_in_dp/i_inq_din_d1/N110 ), .CLK(rclk), .Q(n1800) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[106]  ( .D(\fpu_in_dp/i_inq_din_d1/N109 ), .CLK(rclk), .Q(n1799) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[105]  ( .D(\fpu_in_dp/i_inq_din_d1/N108 ), .CLK(rclk), .Q(n1798) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[104]  ( .D(\fpu_in_dp/i_inq_din_d1/N107 ), .CLK(rclk), .Q(n1797) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[103]  ( .D(\fpu_in_dp/i_inq_din_d1/N106 ), .CLK(rclk), .Q(n1796) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[102]  ( .D(\fpu_in_dp/i_inq_din_d1/N105 ), .CLK(rclk), .Q(n1795) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[101]  ( .D(\fpu_in_dp/i_inq_din_d1/N104 ), .CLK(rclk), .Q(n1794) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[100]  ( .D(\fpu_in_dp/i_inq_din_d1/N103 ), .CLK(rclk), .Q(n1793) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[99]  ( .D(\fpu_in_dp/i_inq_din_d1/N102 ), 
        .CLK(rclk), .Q(n1792) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[98]  ( .D(\fpu_in_dp/i_inq_din_d1/N101 ), 
        .CLK(rclk), .Q(n1790) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[97]  ( .D(\fpu_in_dp/i_inq_din_d1/N100 ), 
        .CLK(rclk), .Q(n1789) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[96]  ( .D(\fpu_in_dp/i_inq_din_d1/N99 ), 
        .CLK(rclk), .Q(n1788) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[95]  ( .D(\fpu_in_dp/i_inq_din_d1/N98 ), 
        .CLK(rclk), .Q(n1787) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[94]  ( .D(\fpu_in_dp/i_inq_din_d1/N97 ), 
        .CLK(rclk), .Q(n1786) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[93]  ( .D(\fpu_in_dp/i_inq_din_d1/N96 ), 
        .CLK(rclk), .Q(n1785) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[92]  ( .D(\fpu_in_dp/i_inq_din_d1/N95 ), 
        .CLK(rclk), .Q(n1784) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[91]  ( .D(\fpu_in_dp/i_inq_din_d1/N94 ), 
        .CLK(rclk), .Q(n1783) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[90]  ( .D(\fpu_in_dp/i_inq_din_d1/N93 ), 
        .CLK(rclk), .Q(n1782) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[89]  ( .D(\fpu_in_dp/i_inq_din_d1/N92 ), 
        .CLK(rclk), .Q(n1781) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[88]  ( .D(\fpu_in_dp/i_inq_din_d1/N91 ), 
        .CLK(rclk), .Q(n1779) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[87]  ( .D(\fpu_in_dp/i_inq_din_d1/N90 ), 
        .CLK(rclk), .Q(n1778) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[86]  ( .D(\fpu_in_dp/i_inq_din_d1/N89 ), 
        .CLK(rclk), .Q(n1777) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[85]  ( .D(\fpu_in_dp/i_inq_din_d1/N88 ), 
        .CLK(rclk), .Q(n1776) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[84]  ( .D(\fpu_in_dp/i_inq_din_d1/N87 ), 
        .CLK(rclk), .Q(n1775) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[83]  ( .D(\fpu_in_dp/i_inq_din_d1/N86 ), 
        .CLK(rclk), .Q(n1774) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[82]  ( .D(\fpu_in_dp/i_inq_din_d1/N85 ), 
        .CLK(rclk), .Q(n1773) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[81]  ( .D(\fpu_in_dp/i_inq_din_d1/N84 ), 
        .CLK(rclk), .Q(n1772) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[80]  ( .D(\fpu_in_dp/i_inq_din_d1/N83 ), 
        .CLK(rclk), .Q(n1771) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[79]  ( .D(\fpu_in_dp/i_inq_din_d1/N82 ), 
        .CLK(rclk), .Q(n1770) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[78]  ( .D(\fpu_in_dp/i_inq_din_d1/N81 ), 
        .CLK(rclk), .Q(n1832) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[77]  ( .D(\fpu_in_dp/i_inq_din_d1/N80 ), 
        .CLK(rclk), .Q(n1831) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[76]  ( .D(\fpu_in_dp/i_inq_din_d1/N79 ), 
        .CLK(rclk), .Q(n1830) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[75]  ( .D(\fpu_in_dp/i_inq_din_d1/N78 ), 
        .CLK(rclk), .Q(n1829) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[74]  ( .D(\fpu_in_dp/i_inq_din_d1/N77 ), 
        .CLK(rclk), .Q(n1824) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[73]  ( .D(\fpu_in_dp/i_inq_din_d1/N76 ), 
        .CLK(rclk), .Q(n1813) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[72]  ( .D(\fpu_in_dp/i_inq_din_d1/N75 ), 
        .CLK(rclk), .Q(n1802) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[71]  ( .D(\fpu_in_dp/i_inq_din_d1/N74 ), 
        .CLK(rclk), .Q(n1791) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[70]  ( .D(\fpu_in_dp/i_inq_din_d1/N73 ), 
        .CLK(rclk), .Q(n1780) );
  DFFX1 \fpu_in_dp/i_inq_din_d1/q_reg[69]  ( .D(\fpu_in_dp/i_inq_din_d1/N72 ), 
        .CLK(rclk), .Q(n1769) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[68]  ( .D(n1849), .RSTB(
        fp_src2_in[68]), .SETB(1'b1), .CLK(rclk), .Q(n1768) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[67]  ( .D(n1849), .RSTB(
        fp_src2_in[67]), .SETB(1'b1), .CLK(rclk), .Q(n1767) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[66]  ( .D(fp_src2_in[66]), .RSTB(
        n1849), .SETB(1'b1), .CLK(rclk), .Q(n1765) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[65]  ( .D(n1849), .RSTB(
        fp_src2_in[65]), .SETB(1'b1), .CLK(rclk), .Q(n1764) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[64]  ( .D(n1849), .RSTB(
        fp_src2_in[64]), .SETB(1'b1), .CLK(rclk), .Q(n1766) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[63]  ( .D(n1849), .RSTB(
        fp_src2_in[63]), .SETB(1'b1), .CLK(rclk), .Q(n1759) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[62]  ( .D(n1850), .RSTB(
        fp_src2_in[62]), .SETB(1'b1), .CLK(rclk), .Q(n1758) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[61]  ( .D(n1849), .RSTB(
        fp_src2_in[61]), .SETB(1'b1), .CLK(rclk), .Q(n1757) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[60]  ( .D(n1850), .RSTB(
        fp_src2_in[60]), .SETB(1'b1), .CLK(rclk), .Q(n1756) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[59]  ( .D(n1849), .RSTB(
        fp_src2_in[59]), .SETB(1'b1), .CLK(rclk), .Q(n1754) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[58]  ( .D(n1849), .RSTB(
        fp_src2_in[58]), .SETB(1'b1), .CLK(rclk), .Q(n1753) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[57]  ( .D(n1849), .RSTB(
        fp_src2_in[57]), .SETB(1'b1), .CLK(rclk), .Q(n1752) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[56]  ( .D(n1849), .RSTB(
        fp_src2_in[56]), .SETB(1'b1), .CLK(rclk), .Q(n1751) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[55]  ( .D(n1849), .RSTB(
        fp_src2_in[55]), .SETB(1'b1), .CLK(rclk), .Q(n1750) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[54]  ( .D(n1850), .RSTB(
        fp_src2_in[54]), .SETB(1'b1), .CLK(rclk), .Q(n1749) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[53]  ( .D(n1849), .RSTB(
        fp_src2_in[53]), .SETB(1'b1), .CLK(rclk), .Q(n1748) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[52]  ( .D(n1850), .RSTB(
        fp_src2_in[52]), .SETB(1'b1), .CLK(rclk), .Q(n1747) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[51]  ( .D(n1849), .RSTB(
        fp_src2_in[51]), .SETB(1'b1), .CLK(rclk), .Q(n1746) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[50]  ( .D(n1849), .RSTB(
        fp_src2_in[50]), .SETB(1'b1), .CLK(rclk), .Q(n1745) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[49]  ( .D(n1849), .RSTB(
        fp_src2_in[49]), .SETB(1'b1), .CLK(rclk), .Q(n1743) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[48]  ( .D(n1849), .RSTB(
        fp_src2_in[48]), .SETB(1'b1), .CLK(rclk), .Q(n1742) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[47]  ( .D(n1849), .RSTB(
        fp_src2_in[47]), .SETB(1'b1), .CLK(rclk), .Q(n1741) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[46]  ( .D(n1849), .RSTB(
        fp_src2_in[46]), .SETB(1'b1), .CLK(rclk), .Q(n1740) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[45]  ( .D(n1850), .RSTB(
        fp_src2_in[45]), .SETB(1'b1), .CLK(rclk), .Q(n1739) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[44]  ( .D(n1849), .RSTB(
        fp_src2_in[44]), .SETB(1'b1), .CLK(rclk), .Q(n1738) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[43]  ( .D(n1849), .RSTB(
        fp_src2_in[43]), .SETB(1'b1), .CLK(rclk), .Q(n1737) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[42]  ( .D(n1849), .RSTB(
        fp_src2_in[42]), .SETB(1'b1), .CLK(rclk), .Q(n1736) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[41]  ( .D(n1850), .RSTB(
        fp_src2_in[41]), .SETB(1'b1), .CLK(rclk), .Q(n1735) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[40]  ( .D(n1849), .RSTB(
        fp_src2_in[40]), .SETB(1'b1), .CLK(rclk), .Q(n1734) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[39]  ( .D(n1849), .RSTB(
        fp_src2_in[39]), .SETB(1'b1), .CLK(rclk), .Q(n1732) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[38]  ( .D(n1849), .RSTB(
        fp_src2_in[38]), .SETB(1'b1), .CLK(rclk), .Q(n1731) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[37]  ( .D(n1849), .RSTB(
        fp_src2_in[37]), .SETB(1'b1), .CLK(rclk), .Q(n1730) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[36]  ( .D(n1849), .RSTB(
        fp_src2_in[36]), .SETB(1'b1), .CLK(rclk), .Q(n1729) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[35]  ( .D(n1850), .RSTB(
        fp_src2_in[35]), .SETB(1'b1), .CLK(rclk), .Q(n1728) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[34]  ( .D(n1850), .RSTB(
        fp_src2_in[34]), .SETB(1'b1), .CLK(rclk), .Q(n1727) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[33]  ( .D(n1850), .RSTB(
        fp_src2_in[33]), .SETB(1'b1), .CLK(rclk), .Q(n1726) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[32]  ( .D(n1849), .RSTB(
        fp_src2_in[32]), .SETB(1'b1), .CLK(rclk), .Q(n1725) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[31]  ( .D(n1850), .RSTB(
        fp_src2_in[31]), .SETB(1'b1), .CLK(rclk), .Q(n1724) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[30]  ( .D(n1849), .RSTB(
        fp_src2_in[30]), .SETB(1'b1), .CLK(rclk), .Q(n1723) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[29]  ( .D(n1849), .RSTB(
        fp_src2_in[29]), .SETB(1'b1), .CLK(rclk), .Q(n1721) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[28]  ( .D(n1850), .RSTB(
        fp_src2_in[28]), .SETB(1'b1), .CLK(rclk), .Q(n1720) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[27]  ( .D(n1850), .RSTB(
        fp_src2_in[27]), .SETB(1'b1), .CLK(rclk), .Q(n1719) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[26]  ( .D(n1849), .RSTB(
        fp_src2_in[26]), .SETB(1'b1), .CLK(rclk), .Q(n1718) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[25]  ( .D(n1849), .RSTB(
        fp_src2_in[25]), .SETB(1'b1), .CLK(rclk), .Q(n1717) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[24]  ( .D(n1849), .RSTB(
        fp_src2_in[24]), .SETB(1'b1), .CLK(rclk), .Q(n1716) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[23]  ( .D(n1849), .RSTB(
        fp_src2_in[23]), .SETB(1'b1), .CLK(rclk), .Q(n1715) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[22]  ( .D(n1850), .RSTB(
        fp_src2_in[22]), .SETB(1'b1), .CLK(rclk), .Q(n1714) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[21]  ( .D(n1849), .RSTB(
        fp_src2_in[21]), .SETB(1'b1), .CLK(rclk), .Q(n1713) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[20]  ( .D(n1849), .RSTB(
        fp_src2_in[20]), .SETB(1'b1), .CLK(rclk), .Q(n1712) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[19]  ( .D(n1849), .RSTB(
        fp_src2_in[19]), .SETB(1'b1), .CLK(rclk), .Q(n1710) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[18]  ( .D(n1849), .RSTB(
        fp_src2_in[18]), .SETB(1'b1), .CLK(rclk), .Q(n1709) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[17]  ( .D(n1850), .RSTB(
        fp_src2_in[17]), .SETB(1'b1), .CLK(rclk), .Q(n1708) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[16]  ( .D(n1849), .RSTB(
        fp_src2_in[16]), .SETB(1'b1), .CLK(rclk), .Q(n1707) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[15]  ( .D(n1849), .RSTB(
        fp_src2_in[15]), .SETB(1'b1), .CLK(rclk), .Q(n1706) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[14]  ( .D(n1849), .RSTB(
        fp_src2_in[14]), .SETB(1'b1), .CLK(rclk), .Q(n1705) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[13]  ( .D(n1850), .RSTB(
        fp_src2_in[13]), .SETB(1'b1), .CLK(rclk), .Q(n1704) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[12]  ( .D(n1849), .RSTB(
        fp_src2_in[12]), .SETB(1'b1), .CLK(rclk), .Q(n1703) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[11]  ( .D(n1850), .RSTB(
        fp_src2_in[11]), .SETB(1'b1), .CLK(rclk), .Q(n1702) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[10]  ( .D(n1849), .RSTB(
        fp_src2_in[10]), .SETB(1'b1), .CLK(rclk), .Q(n1701) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[9]  ( .D(n1849), .RSTB(fp_src2_in[9]), 
        .SETB(1'b1), .CLK(rclk), .Q(n1763) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[8]  ( .D(n1849), .RSTB(fp_src2_in[8]), 
        .SETB(1'b1), .CLK(rclk), .Q(n1762) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[7]  ( .D(n1850), .RSTB(fp_src2_in[7]), 
        .SETB(1'b1), .CLK(rclk), .Q(n1761) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[6]  ( .D(n1849), .RSTB(fp_src2_in[6]), 
        .SETB(1'b1), .CLK(rclk), .Q(n1760) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[5]  ( .D(n1849), .RSTB(fp_src2_in[5]), 
        .SETB(1'b1), .CLK(rclk), .Q(n1755) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[4]  ( .D(n1850), .RSTB(fp_src2_in[4]), 
        .SETB(1'b1), .CLK(rclk), .Q(n1744) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[3]  ( .D(n1850), .RSTB(fp_src2_in[3]), 
        .SETB(1'b1), .CLK(rclk), .Q(n1733) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[2]  ( .D(n1850), .RSTB(fp_src2_in[2]), 
        .SETB(1'b1), .CLK(rclk), .Q(n1722) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[1]  ( .D(n1850), .RSTB(fp_src2_in[1]), 
        .SETB(1'b1), .CLK(rclk), .Q(n1711) );
  DFFSSRX1 \fpu_in_dp/i_inq_din_d1/q_reg[0]  ( .D(n1849), .RSTB(fp_src2_in[0]), 
        .SETB(1'b1), .CLK(rclk), .Q(n1700) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[68]  ( .D(\fpu_in_dp/n646 ), .CLK(rclk), 
        .Q(n819) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[67]  ( .D(\fpu_in_dp/n647 ), .CLK(rclk), 
        .Q(n820) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[66]  ( .D(\fpu_in_dp/n648 ), .CLK(rclk), 
        .Q(n821) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[65]  ( .D(\fpu_in_dp/n649 ), .CLK(rclk), 
        .Q(n822) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[64]  ( .D(\fpu_in_dp/n650 ), .CLK(rclk), 
        .Q(n823) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[63]  ( .D(\fpu_in_dp/n651 ), .CLK(rclk), 
        .Q(n824) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[62]  ( .D(\fpu_in_dp/n652 ), .CLK(rclk), 
        .Q(n825) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[61]  ( .D(\fpu_in_dp/n653 ), .CLK(rclk), 
        .Q(n826) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[60]  ( .D(\fpu_in_dp/n654 ), .CLK(rclk), 
        .Q(n827) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[59]  ( .D(\fpu_in_dp/n655 ), .CLK(rclk), 
        .Q(n829) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[58]  ( .D(\fpu_in_dp/n656 ), .CLK(rclk), 
        .Q(n830) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[57]  ( .D(\fpu_in_dp/n657 ), .CLK(rclk), 
        .Q(n831) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[56]  ( .D(\fpu_in_dp/n658 ), .CLK(rclk), 
        .Q(n832) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[55]  ( .D(\fpu_in_dp/n659 ), .CLK(rclk), 
        .Q(n833) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[54]  ( .D(\fpu_in_dp/n660 ), .CLK(rclk), 
        .Q(n834) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[53]  ( .D(\fpu_in_dp/n661 ), .CLK(rclk), 
        .Q(n835) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[52]  ( .D(\fpu_in_dp/n662 ), .CLK(rclk), 
        .Q(n836) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[51]  ( .D(\fpu_in_dp/n663 ), .CLK(rclk), 
        .Q(n837) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[50]  ( .D(\fpu_in_dp/n664 ), .CLK(rclk), 
        .Q(n838) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[49]  ( .D(\fpu_in_dp/n665 ), .CLK(rclk), 
        .Q(n840) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[48]  ( .D(\fpu_in_dp/n666 ), .CLK(rclk), 
        .Q(n841) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[47]  ( .D(\fpu_in_dp/n667 ), .CLK(rclk), 
        .Q(n842) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[46]  ( .D(\fpu_in_dp/n668 ), .CLK(rclk), 
        .Q(n843) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[45]  ( .D(\fpu_in_dp/n669 ), .CLK(rclk), 
        .Q(n844) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[44]  ( .D(\fpu_in_dp/n670 ), .CLK(rclk), 
        .Q(n845) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[43]  ( .D(\fpu_in_dp/n671 ), .CLK(rclk), 
        .Q(n846) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[42]  ( .D(\fpu_in_dp/n672 ), .CLK(rclk), 
        .Q(n847) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[41]  ( .D(\fpu_in_dp/n673 ), .CLK(rclk), 
        .Q(n848) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[40]  ( .D(\fpu_in_dp/n674 ), .CLK(rclk), 
        .Q(n849) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[39]  ( .D(\fpu_in_dp/n675 ), .CLK(rclk), 
        .Q(n851) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[38]  ( .D(\fpu_in_dp/n676 ), .CLK(rclk), 
        .Q(n852) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[37]  ( .D(\fpu_in_dp/n677 ), .CLK(rclk), 
        .Q(n853) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[36]  ( .D(\fpu_in_dp/n678 ), .CLK(rclk), 
        .Q(n854) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[35]  ( .D(\fpu_in_dp/n679 ), .CLK(rclk), 
        .Q(n855) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[34]  ( .D(\fpu_in_dp/n680 ), .CLK(rclk), 
        .Q(n856) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[33]  ( .D(\fpu_in_dp/n681 ), .CLK(rclk), 
        .Q(n857) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[32]  ( .D(\fpu_in_dp/n682 ), .CLK(rclk), 
        .Q(n858) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[31]  ( .D(\fpu_in_dp/n683 ), .CLK(rclk), 
        .Q(n859) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[30]  ( .D(\fpu_in_dp/n684 ), .CLK(rclk), 
        .Q(n860) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[29]  ( .D(\fpu_in_dp/n685 ), .CLK(rclk), 
        .Q(n862) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[28]  ( .D(\fpu_in_dp/n686 ), .CLK(rclk), 
        .Q(n863) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[27]  ( .D(\fpu_in_dp/n687 ), .CLK(rclk), 
        .Q(n864) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[26]  ( .D(\fpu_in_dp/n688 ), .CLK(rclk), 
        .Q(n865) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[25]  ( .D(\fpu_in_dp/n689 ), .CLK(rclk), 
        .Q(n866) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[24]  ( .D(\fpu_in_dp/n690 ), .CLK(rclk), 
        .Q(n867) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[23]  ( .D(\fpu_in_dp/n691 ), .CLK(rclk), 
        .Q(n868) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[22]  ( .D(\fpu_in_dp/n692 ), .CLK(rclk), 
        .Q(n869) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[21]  ( .D(\fpu_in_dp/n693 ), .CLK(rclk), 
        .Q(n870) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[20]  ( .D(\fpu_in_dp/n694 ), .CLK(rclk), 
        .Q(n871) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[19]  ( .D(\fpu_in_dp/n695 ), .CLK(rclk), 
        .Q(n873) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[18]  ( .D(\fpu_in_dp/n696 ), .CLK(rclk), 
        .Q(n874) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[17]  ( .D(\fpu_in_dp/n697 ), .CLK(rclk), 
        .Q(n875) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[16]  ( .D(\fpu_in_dp/n698 ), .CLK(rclk), 
        .Q(n876) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[15]  ( .D(\fpu_in_dp/n699 ), .CLK(rclk), 
        .Q(n877) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[14]  ( .D(\fpu_in_dp/n700 ), .CLK(rclk), 
        .Q(n878) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[13]  ( .D(\fpu_in_dp/n701 ), .CLK(rclk), 
        .Q(n879) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[12]  ( .D(\fpu_in_dp/n702 ), .CLK(rclk), 
        .Q(n880) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[11]  ( .D(\fpu_in_dp/n703 ), .CLK(rclk), 
        .Q(n881) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[10]  ( .D(\fpu_in_dp/n704 ), .CLK(rclk), 
        .Q(n882) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[9]  ( .D(\fpu_in_dp/n705 ), .CLK(rclk), 
        .Q(n815) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[8]  ( .D(\fpu_in_dp/n706 ), .CLK(rclk), 
        .Q(n816) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[7]  ( .D(\fpu_in_dp/n707 ), .CLK(rclk), 
        .Q(n817) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[6]  ( .D(\fpu_in_dp/n708 ), .CLK(rclk), 
        .Q(n818) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[5]  ( .D(\fpu_in_dp/n709 ), .CLK(rclk), 
        .Q(n828) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[4]  ( .D(\fpu_in_dp/n710 ), .CLK(rclk), 
        .Q(n839) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[3]  ( .D(\fpu_in_dp/n711 ), .CLK(rclk), 
        .Q(n850) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[2]  ( .D(\fpu_in_dp/n712 ), .CLK(rclk), 
        .Q(n861) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[1]  ( .D(\fpu_in_dp/n713 ), .CLK(rclk), 
        .Q(n872) );
  DFFX1 \fpu_in_dp/i_fp_srcb_in/q_reg[0]  ( .D(\fpu_in_dp/n714 ), .CLK(rclk), 
        .Q(n883) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[63]  ( .D(pcx_fpio_data_px2[63]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n803) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[62]  ( .D(pcx_fpio_data_px2[62]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n763), .QN(n1656) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[61]  ( .D(pcx_fpio_data_px2[61]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n767), .QN(n1623) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[60]  ( .D(pcx_fpio_data_px2[60]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n757), .QN(n1636) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[59]  ( .D(pcx_fpio_data_px2[59]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n735), .QN(n1680) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[58]  ( .D(pcx_fpio_data_px2[58]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n744), .QN(n1676) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[57]  ( .D(pcx_fpio_data_px2[57]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n739), .QN(n1654) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[56]  ( .D(pcx_fpio_data_px2[56]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n748), .QN(n1678) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[55]  ( .D(pcx_fpio_data_px2[55]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n742), .QN(n1655) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[54]  ( .D(pcx_fpio_data_px2[54]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n759), .QN(n1694) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[53]  ( .D(pcx_fpio_data_px2[53]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n743), .QN(n1653) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[52]  ( .D(pcx_fpio_data_px2[52]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n738), .QN(n1635) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[51]  ( .D(pcx_fpio_data_px2[51]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n758), .QN(n1674) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[50]  ( .D(pcx_fpio_data_px2[50]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n773) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[49]  ( .D(pcx_fpio_data_px2[49]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n786), .QN(n1660) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[48]  ( .D(pcx_fpio_data_px2[48]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n796), .QN(n1626) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[47]  ( .D(pcx_fpio_data_px2[47]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n765) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[46]  ( .D(pcx_fpio_data_px2[46]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n751) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[45]  ( .D(pcx_fpio_data_px2[45]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n764) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[44]  ( .D(pcx_fpio_data_px2[44]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n749), .QN(n1681) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[43]  ( .D(pcx_fpio_data_px2[43]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n750), .QN(n1658) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[42]  ( .D(pcx_fpio_data_px2[42]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n787), .QN(n1624) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[41]  ( .D(pcx_fpio_data_px2[41]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n774), .QN(n1637) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[40]  ( .D(pcx_fpio_data_px2[40]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n797), .QN(n1638) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[39]  ( .D(pcx_fpio_data_px2[39]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n766), .QN(n1683) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[38]  ( .D(pcx_fpio_data_px2[38]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n789), .QN(n1659) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[37]  ( .D(pcx_fpio_data_px2[37]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n775), .QN(n1625) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[36]  ( .D(pcx_fpio_data_px2[36]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n798), .QN(n1640) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[35]  ( .D(pcx_fpio_data_px2[35]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n790), .QN(n1657) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[34]  ( .D(pcx_fpio_data_px2[34]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n776), .QN(n1639) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[33]  ( .D(pcx_fpio_data_px2[33]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n777), .QN(n1684) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[32]  ( .D(pcx_fpio_data_px2[32]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n799), .QN(n1685) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[31]  ( .D(pcx_fpio_data_px2[31]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n769), .QN(n1686) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[30]  ( .D(pcx_fpio_data_px2[30]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n768), .QN(n1662) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[29]  ( .D(pcx_fpio_data_px2[29]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n745), .QN(n1642) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[28]  ( .D(pcx_fpio_data_px2[28]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n760), .QN(n1687) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[27]  ( .D(pcx_fpio_data_px2[27]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n791), .QN(n1663) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[26]  ( .D(pcx_fpio_data_px2[26]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n779), .QN(n1629) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[25]  ( .D(pcx_fpio_data_px2[25]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n780), .QN(n1643) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[24]  ( .D(pcx_fpio_data_px2[24]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n800), .QN(n1688) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[23]  ( .D(pcx_fpio_data_px2[23]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n736), .QN(n1665) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[22]  ( .D(pcx_fpio_data_px2[22]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n740), .QN(n1631) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[21]  ( .D(pcx_fpio_data_px2[21]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n746), .QN(n1645) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[20]  ( .D(pcx_fpio_data_px2[20]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n761), .QN(n1690) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[19]  ( .D(pcx_fpio_data_px2[19]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n737), .QN(n1630) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[18]  ( .D(pcx_fpio_data_px2[18]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n741), .QN(n1644) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[17]  ( .D(pcx_fpio_data_px2[17]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n747), .QN(n1689) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[16]  ( .D(pcx_fpio_data_px2[16]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n762), .QN(n1667) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[15]  ( .D(pcx_fpio_data_px2[15]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n792), .QN(n1633) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[14]  ( .D(pcx_fpio_data_px2[14]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n782), .QN(n1647) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[13]  ( .D(pcx_fpio_data_px2[13]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n783), .QN(n1692) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[12]  ( .D(pcx_fpio_data_px2[12]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n801), .QN(n1666) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[11]  ( .D(pcx_fpio_data_px2[11]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n793), .QN(n1632) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[10]  ( .D(pcx_fpio_data_px2[10]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n784), .QN(n1646) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[9]  ( .D(pcx_fpio_data_px2[9]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n770), .QN(n1668) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[8]  ( .D(pcx_fpio_data_px2[8]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n794), .QN(n1634) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[7]  ( .D(pcx_fpio_data_px2[7]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n785), .QN(n1648) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[6]  ( .D(pcx_fpio_data_px2[6]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n771), .QN(n1693) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[5]  ( .D(pcx_fpio_data_px2[5]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n772), .QN(n1661) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[4]  ( .D(pcx_fpio_data_px2[4]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n795), .QN(n1627) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[3]  ( .D(pcx_fpio_data_px2[3]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n788), .QN(n1641) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[2]  ( .D(pcx_fpio_data_px2[2]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n778), .QN(n1628) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[1]  ( .D(pcx_fpio_data_px2[1]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(n781), .QN(n1664) );
  DFFSSRX1 \fpu_in_dp/i_fp_srca_in/q_reg[0]  ( .D(pcx_fpio_data_px2[0]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(n802), .QN(n1691) );
  DFFSSRX1 \fpu_in_dp/i_fp_rnd_mode_in/q_reg[1]  ( .D(pcx_fpio_data_px2[65]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(fp_rnd_mode_in[1]), .QN(
        \fpu_in_dp/n439 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_rnd_mode_in/q_reg[0]  ( .D(pcx_fpio_data_px2[64]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_rnd_mode_in[0]), .QN(
        \fpu_in_dp/n441 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_fcc_in/q_reg[1]  ( .D(pcx_fpio_data_px2[67]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_fcc_in[1]), .QN(
        \fpu_in_dp/n443 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_fcc_in/q_reg[0]  ( .D(pcx_fpio_data_px2[66]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(fp_fcc_in[0]), .QN(
        \fpu_in_dp/n445 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_op_in/q_reg[7]  ( .D(pcx_fpio_data_px2[79]), .RSTB(
        n1850), .SETB(1'b1), .CLK(rclk), .Q(fp_op_in_7in), .QN(
        \fpu_in_dp/n105 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_op_in/q_reg[6]  ( .D(pcx_fpio_data_px2[78]), .RSTB(
        n1850), .SETB(1'b1), .CLK(rclk), .Q(fp_op_in[6]), .QN(\fpu_in_dp/n448 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_op_in/q_reg[5]  ( .D(pcx_fpio_data_px2[77]), .RSTB(
        n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_op_in[5]), .QN(\fpu_in_dp/n450 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_op_in/q_reg[4]  ( .D(pcx_fpio_data_px2[76]), .RSTB(
        n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_op_in[4]), .QN(\fpu_in_dp/n452 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_op_in/q_reg[3]  ( .D(pcx_fpio_data_px2[75]), .RSTB(
        n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_op_in[3]), .QN(\fpu_in_dp/n454 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_op_in/q_reg[2]  ( .D(pcx_fpio_data_px2[74]), .RSTB(
        n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_op_in[2]), .QN(\fpu_in_dp/n456 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_op_in/q_reg[1]  ( .D(pcx_fpio_data_px2[73]), .RSTB(
        n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_op_in[1]), .QN(\fpu_in_dp/n458 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_op_in/q_reg[0]  ( .D(pcx_fpio_data_px2[72]), .RSTB(
        n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_op_in[0]), .QN(\fpu_in_dp/n473 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_id_in/q_reg[4]  ( .D(pcx_fpio_data_px2[116]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_id_in[4]), .QN(
        \fpu_in_dp/n461 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_id_in/q_reg[3]  ( .D(pcx_fpio_data_px2[115]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_id_in[3]), .QN(
        \fpu_in_dp/n463 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_id_in/q_reg[2]  ( .D(pcx_fpio_data_px2[114]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_id_in[2]), .QN(
        \fpu_in_dp/n465 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_id_in/q_reg[1]  ( .D(pcx_fpio_data_px2[113]), 
        .RSTB(n1849), .SETB(1'b1), .CLK(rclk), .Q(fp_id_in[1]), .QN(
        \fpu_in_dp/n467 ) );
  DFFSSRX1 \fpu_in_dp/i_fp_id_in/q_reg[0]  ( .D(pcx_fpio_data_px2[112]), 
        .RSTB(n1850), .SETB(1'b1), .CLK(rclk), .Q(fp_id_in[0]), .QN(
        \fpu_in_dp/n469 ) );
  OA221X1 U1482 ( .IN1(1'b0), .IN2(n1848), .IN3(n1888), .IN4(n1671), .IN5(
        n1889), .Q(\fpu_in_ctl/i_inq_div_rdptr/N5 ) );
  OA221X1 U1483 ( .IN1(1'b0), .IN2(\fpu_in_ctl/in_ctl_rst_l ), .IN3(n756), 
        .IN4(n1926), .IN5(n1927), .Q(n257) );
  OA221X1 U1484 ( .IN1(1'b0), .IN2(\fpu_in_ctl/in_ctl_rst_l ), .IN3(n1564), 
        .IN4(n1929), .IN5(n1928), .Q(n255) );
  INVX0 U1485 ( .INP(n1895), .ZN(n1904) );
  NOR2X0 U1486 ( .IN1(n1970), .IN2(n1948), .QN(n1943) );
  NOR2X0 U1487 ( .IN1(n1966), .IN2(n1970), .QN(n1956) );
  NOR2X0 U1488 ( .IN1(n1673), .IN2(n1942), .QN(n1948) );
  INVX0 U1489 ( .INP(n1986), .ZN(n1887) );
  INVX0 U1490 ( .INP(n1856), .ZN(n1938) );
  INVX0 U1491 ( .INP(n1896), .ZN(n1899) );
  INVX0 U1492 ( .INP(n1897), .ZN(n1898) );
  INVX0 U1493 ( .INP(n1901), .ZN(n1886) );
  NAND2X1 U1494 ( .IN1(n1682), .IN2(n1931), .QN(n1868) );
  NOR2X0 U1495 ( .IN1(n1672), .IN2(n1927), .QN(n1929) );
  NAND2X1 U1496 ( .IN1(n1564), .IN2(n1929), .QN(n1928) );
  NAND2X1 U1497 ( .IN1(n756), .IN2(n1926), .QN(n1927) );
  NOR2X0 U1498 ( .IN1(n1926), .IN2(n1942), .QN(n1894) );
  NAND2X1 U1499 ( .IN1(n1867), .IN2(n1868), .QN(n1905) );
  NAND2X1 U1500 ( .IN1(n1943), .IN2(n1955), .QN(n1946) );
  NAND2X1 U1501 ( .IN1(n1943), .IN2(n1953), .QN(n1941) );
  NAND2X1 U1502 ( .IN1(n1943), .IN2(n1951), .QN(n1940) );
  NAND2X1 U1503 ( .IN1(n1943), .IN2(n1963), .QN(n1939) );
  NOR2X0 U1504 ( .IN1(n1670), .IN2(n1650), .QN(n1959) );
  NAND2X1 U1505 ( .IN1(n1956), .IN2(n1955), .QN(n1960) );
  NAND2X1 U1506 ( .IN1(n1956), .IN2(n1953), .QN(n1954) );
  NAND2X1 U1507 ( .IN1(n1956), .IN2(n1951), .QN(n1952) );
  NOR2X0 U1508 ( .IN1(n1949), .IN2(n1964), .QN(n1958) );
  NAND2X1 U1509 ( .IN1(n1973), .IN2(n1848), .QN(n1962) );
  INVX0 U1510 ( .INP(n1961), .ZN(n1966) );
  NOR2X0 U1511 ( .IN1(n807), .IN2(n886), .QN(n1967) );
  NAND2X1 U1512 ( .IN1(n1967), .IN2(n1972), .QN(n1965) );
  NAND2X1 U1513 ( .IN1(n1972), .IN2(n1948), .QN(n1964) );
  NOR2X0 U1514 ( .IN1(n1650), .IN2(n807), .QN(n1969) );
  NOR2X0 U1515 ( .IN1(n1670), .IN2(n886), .QN(n1968) );
  INVX0 U1516 ( .INP(n1962), .ZN(n1970) );
  NAND2X1 U1517 ( .IN1(n1985), .IN2(inq_we), .QN(n1973) );
  INVX0 U1518 ( .INP(n1973), .ZN(n1972) );
  NOR2X0 U1519 ( .IN1(n1159), .IN2(n1942), .QN(n1892) );
  INVX0 U1520 ( .INP(n1974), .ZN(n1982) );
  NOR2X0 U1521 ( .IN1(n1980), .IN2(n1979), .QN(n1981) );
  NOR2X0 U1522 ( .IN1(n1649), .IN2(n1675), .QN(n1978) );
  NOR2X0 U1523 ( .IN1(n889), .IN2(n754), .QN(n1976) );
  NOR2X0 U1524 ( .IN1(n754), .IN2(n1649), .QN(n1975) );
  INVX0 U1525 ( .INP(n1979), .ZN(n1977) );
  NOR2X0 U1526 ( .IN1(n1980), .IN2(n1974), .QN(n1983) );
  INVX0 U1527 ( .INP(inq_wraddr[3]), .ZN(n1985) );
  NOR2X0 U1528 ( .IN1(n418), .IN2(n1159), .QN(n1930) );
  NAND2X1 U1529 ( .IN1(n1888), .IN2(n1671), .QN(n1889) );
  NAND2X1 U1530 ( .IN1(inq_div), .IN2(d1stg_step), .QN(n1986) );
  NOR2X0 U1531 ( .IN1(n1887), .IN2(n1942), .QN(n1890) );
  NOR2X0 U1532 ( .IN1(n1942), .IN2(n1986), .QN(n1891) );
  NAND2X1 U1533 ( .IN1(n1932), .IN2(n1931), .QN(inq_read_en) );
  NOR2X0 U1534 ( .IN1(n1844), .IN2(n1628), .QN(fp_src1_in[2]) );
  NOR2X0 U1535 ( .IN1(n1844), .IN2(n1641), .QN(fp_src1_in[3]) );
  NOR2X0 U1536 ( .IN1(n1844), .IN2(n1627), .QN(fp_src1_in[4]) );
  NOR2X0 U1537 ( .IN1(n1844), .IN2(n1661), .QN(fp_src1_in[5]) );
  NOR2X0 U1538 ( .IN1(n1844), .IN2(n1634), .QN(fp_src1_in[8]) );
  NOR2X0 U1539 ( .IN1(n1844), .IN2(n1668), .QN(fp_src1_in[9]) );
  NOR2X0 U1540 ( .IN1(fp_op_in_7in), .IN2(n1689), .QN(fp_src1_in[17]) );
  NOR2X0 U1541 ( .IN1(fp_op_in_7in), .IN2(n1645), .QN(fp_src1_in[21]) );
  NOR2X0 U1542 ( .IN1(fp_op_in_7in), .IN2(n1643), .QN(fp_src1_in[25]) );
  NOR2X0 U1543 ( .IN1(n1844), .IN2(n1629), .QN(fp_src1_in[26]) );
  NOR2X0 U1544 ( .IN1(fp_op_in_7in), .IN2(n1663), .QN(fp_src1_in[27]) );
  NOR2X0 U1545 ( .IN1(n1844), .IN2(n1687), .QN(fp_src1_in[28]) );
  NOR2X0 U1546 ( .IN1(n1844), .IN2(n1642), .QN(fp_src1_in[29]) );
  NOR2X0 U1547 ( .IN1(n1844), .IN2(n1684), .QN(fp_src1_in[33]) );
  NOR2X0 U1548 ( .IN1(n1844), .IN2(n1639), .QN(fp_src1_in[34]) );
  NOR2X0 U1549 ( .IN1(n1844), .IN2(n1640), .QN(fp_src1_in[36]) );
  NOR2X0 U1550 ( .IN1(n1844), .IN2(n1659), .QN(fp_src1_in[38]) );
  NOR2X0 U1551 ( .IN1(fp_op_in_7in), .IN2(n1683), .QN(fp_src1_in[39]) );
  NOR2X0 U1552 ( .IN1(n1844), .IN2(n1637), .QN(fp_src1_in[41]) );
  NOR2X0 U1553 ( .IN1(n1844), .IN2(n1624), .QN(fp_src1_in[42]) );
  NOR2X0 U1554 ( .IN1(n1844), .IN2(n1658), .QN(fp_src1_in[43]) );
  NOR2X0 U1555 ( .IN1(n1844), .IN2(n1660), .QN(fp_src1_in[49]) );
  NOR2X0 U1556 ( .IN1(n1844), .IN2(n1694), .QN(fp_src1_in[54]) );
  NOR2X0 U1557 ( .IN1(n1844), .IN2(n1655), .QN(fp_src1_in[55]) );
  NOR2X0 U1558 ( .IN1(n1844), .IN2(n1676), .QN(fp_src1_in[58]) );
  NOR2X0 U1559 ( .IN1(n1844), .IN2(n1623), .QN(fp_src1_in[61]) );
  NOR2X0 U1560 ( .IN1(n1844), .IN2(n1656), .QN(fp_src1_in[62]) );
  NOR2X0 U1561 ( .IN1(n1886), .IN2(n1844), .QN(fp_src1_in[65]) );
  NOR2X0 U1562 ( .IN1(se), .IN2(\fpu_in_dp/n473 ), .QN(
        \fpu_in_dp/i_inq_din_d1/N141 ) );
  NOR2X0 U1563 ( .IN1(\fpu_in_dp/n105 ), .IN2(se), .QN(
        \fpu_in_dp/i_inq_din_d1/N148 ) );
  INVX0 U1564 ( .INP(inq_rdaddr[3]), .ZN(n1159) );
  INVX0 U1565 ( .INP(n1988), .ZN(n1155) );
  NOR2X0 U1566 ( .IN1(se), .IN2(n1159), .QN(\fpu_in_ctl/i_inq_rdaddr_del/N6 )
         );
  NOR2X0 U1567 ( .IN1(\fpu_in_dp/n456 ), .IN2(n1949), .QN(inq_wraddr[3]) );
  NOR2X0 U1568 ( .IN1(n1895), .IN2(n1942), .QN(
        \fpu_in_ctl/i_valid_packet_dly/N7 ) );
  INVX0 U1569 ( .INP(n1942), .ZN(n1848) );
  AO22X1 U1570 ( .IN1(n1669), .IN2(n1554), .IN3(n1696), .IN4(n1558), .Q(n1589)
         );
  AO22X1 U1571 ( .IN1(n1695), .IN2(n1555), .IN3(n1556), .IN4(n1557), .Q(n1590)
         );
  AO22X1 U1572 ( .IN1(n1553), .IN2(n912), .IN3(n1551), .IN4(n911), .Q(n1591)
         );
  AO22X1 U1573 ( .IN1(n1550), .IN2(n913), .IN3(n1552), .IN4(n914), .Q(n1592)
         );
  NOR4X0 U1574 ( .IN1(n1589), .IN2(n1590), .IN3(n1591), .IN4(n1592), .QN(n1593) );
  NOR2X0 U1575 ( .IN1(n1905), .IN2(n1593), .QN(n1594) );
  NOR2X0 U1576 ( .IN1(n1867), .IN2(n890), .QN(n1595) );
  AO21X1 U1577 ( .IN1(n1595), .IN2(n1549), .IN3(n1594), .Q(inq_div) );
  AO22X1 U1578 ( .IN1(n904), .IN2(n1577), .IN3(n906), .IN4(n1579), .Q(n1596)
         );
  AO22X1 U1579 ( .IN1(n902), .IN2(n1575), .IN3(n900), .IN4(n1573), .Q(n1597)
         );
  AO22X1 U1580 ( .IN1(n896), .IN2(n1580), .IN3(n898), .IN4(n1574), .Q(n1598)
         );
  AO22X1 U1581 ( .IN1(n892), .IN2(n1576), .IN3(n894), .IN4(n1578), .Q(n1599)
         );
  NOR4X0 U1582 ( .IN1(n1596), .IN2(n1597), .IN3(n1598), .IN4(n1599), .QN(n1600) );
  NOR2X0 U1583 ( .IN1(n1905), .IN2(n1600), .QN(n1601) );
  NOR2X0 U1584 ( .IN1(n1868), .IN2(n1949), .QN(n1602) );
  AO21X1 U1585 ( .IN1(n1602), .IN2(\fpu_in_dp/n456 ), .IN3(n1601), .Q(inq_mul)
         );
  AOI22X1 U1587 ( .IN1(n1848), .IN2(n755), .IN3(n1891), .IN4(n813), .QN(n1604)
         );
  NOR2X0 U1588 ( .IN1(n1888), .IN2(n1604), .QN(\fpu_in_ctl/i_inq_div_rdptr/N4 ) );
  NAND4X0 U1589 ( .IN1(n1656), .IN2(n1623), .IN3(n1636), .IN4(n1680), .QN(
        n1605) );
  NOR3X0 U1590 ( .IN1(n739), .IN2(n744), .IN3(n1605), .QN(n1606) );
  NOR2X0 U1591 ( .IN1(n738), .IN2(n743), .QN(n1607) );
  AO21X1 U1592 ( .IN1(n1607), .IN2(n1694), .IN3(\fpu_in_dp/n458 ), .Q(n1608)
         );
  NAND4X0 U1593 ( .IN1(n1655), .IN2(n1678), .IN3(n1606), .IN4(n1608), .QN(
        n1896) );
  INVX0 U1594 ( .INP(n1927), .ZN(n1609) );
  OA221X1 U1595 ( .IN1(n1927), .IN2(n1672), .IN3(n1609), .IN4(n814), .IN5(
        \fpu_in_ctl/in_ctl_rst_l ), .Q(n256) );
  NAND3X0 U1596 ( .IN1(n1963), .IN2(n1964), .IN3(n1962), .QN(n1610) );
  NOR2X0 U1597 ( .IN1(n1961), .IN2(n1965), .QN(n1611) );
  MUX21X1 U1598 ( .IN1(n1611), .IN2(n1610), .S(n1566), .Q(n346) );
  INVX0 U1599 ( .INP(n1889), .ZN(n1612) );
  OA221X1 U1600 ( .IN1(n1889), .IN2(n1562), .IN3(n1612), .IN4(n1677), .IN5(
        n1848), .Q(\fpu_in_ctl/i_inq_div_rdptr/N6 ) );
  NAND3X0 U1601 ( .IN1(n743), .IN2(n759), .IN3(n738), .QN(n1613) );
  NAND2X0 U1602 ( .IN1(n1613), .IN2(\fpu_in_dp/n473 ), .QN(n1614) );
  NAND3X0 U1603 ( .IN1(n748), .IN2(n742), .IN3(n1614), .QN(n1615) );
  NAND4X0 U1604 ( .IN1(n763), .IN2(n767), .IN3(n757), .IN4(n735), .QN(n1616)
         );
  NOR4X0 U1605 ( .IN1(n1676), .IN2(n1654), .IN3(n1615), .IN4(n1616), .QN(n1897) );
  INVX0 U1606 ( .INP(n1928), .ZN(n1617) );
  OA221X1 U1607 ( .IN1(n1928), .IN2(n1565), .IN3(n1617), .IN4(n1698), .IN5(
        n1848), .Q(\fpu_in_ctl/i_inq_rdptr/N6 ) );
  INVX0 U1609 ( .INP(n1964), .ZN(n1619) );
  AO22X1 U1610 ( .IN1(n1967), .IN2(n1619), .IN3(n1966), .IN4(n1965), .Q(n347)
         );
  INVX0 U1611 ( .INP(d1stg_step), .ZN(n1620) );
  NOR3X0 U1612 ( .IN1(inq_div), .IN2(n1932), .IN3(n1620), .QN(inq_rdaddr[3])
         );
  NOR2X1 U1614 ( .IN1(n1571), .IN2(se), .QN(n1622) );
  INVX0 U1615 ( .INP(n1934), .ZN(n1842) );
  INVX0 U1616 ( .INP(n1934), .ZN(n1843) );
  INVX0 U1617 ( .INP(n1934), .ZN(n1841) );
  INVX0 U1618 ( .INP(n1935), .ZN(n1840) );
  INVX0 U1619 ( .INP(n1935), .ZN(n1839) );
  INVX0 U1620 ( .INP(n1935), .ZN(n1838) );
  NOR2X1 U1621 ( .IN1(se), .IN2(n1679), .QN(n1903) );
  INVX0 U1622 ( .INP(n1697), .ZN(n1846) );
  INVX0 U1623 ( .INP(n1697), .ZN(n1847) );
  INVX0 U1624 ( .INP(n1697), .ZN(n1845) );
  NAND2X1 U1625 ( .IN1(n1934), .IN2(n1911), .QN(n1935) );
  INVX0 U1626 ( .INP(se), .ZN(n1850) );
  NAND2X1 U1627 ( .IN1(\fpu_in_dp/n105 ), .IN2(n1897), .QN(fp_src1_in[68]) );
  NAND2X1 U1628 ( .IN1(\fpu_in_dp/n105 ), .IN2(n1896), .QN(fp_src1_in[67]) );
  NAND2X1 U1629 ( .IN1(n1673), .IN2(n1848), .QN(n1961) );
  NAND2X1 U1630 ( .IN1(\fpu_in_ctl/in_ctl_rst_l ), .IN2(n41), .QN(n1866) );
  INVX2 U1631 ( .INP(\fpu_in_dp/n105 ), .ZN(n1844) );
  NAND2X1 U1632 ( .IN1(\fpu_in_ctl/in_ctl_rst_l ), .IN2(n8), .QN(n1869) );
  NAND2X1 U1633 ( .IN1(n754), .IN2(n1649), .QN(n1980) );
  NAND2X1 U1634 ( .IN1(\fpu_in_ctl/in_ctl_rst_l ), .IN2(n1850), .QN(n1942) );
  INVX2 U1635 ( .INP(se), .ZN(n1849) );
  NAND3X0 U1636 ( .IN1(n1904), .IN2(n1567), .IN3(\fpu_in_dp/n105 ), .QN(n1856)
         );
  OR2X1 U1637 ( .IN1(n1911), .IN2(n1841), .Q(n1697) );
  NAND3X0 U1638 ( .IN1(n1905), .IN2(n1908), .IN3(n1904), .QN(n1934) );
  INVX0 U1639 ( .INP(sehold), .ZN(n1908) );
  AND2X1 U1640 ( .IN1(\fpu_in_dp/n105 ), .IN2(n764), .Q(fp_src1_in[45]) );
  AND2X1 U1641 ( .IN1(\fpu_in_dp/n105 ), .IN2(n751), .Q(fp_src1_in[46]) );
  AND2X1 U1642 ( .IN1(\fpu_in_dp/n105 ), .IN2(n765), .Q(fp_src1_in[47]) );
  AND2X1 U1643 ( .IN1(\fpu_in_dp/n105 ), .IN2(n773), .Q(fp_src1_in[50]) );
  AND2X1 U1644 ( .IN1(\fpu_in_dp/n105 ), .IN2(n803), .Q(fp_src1_in[63]) );
  AND3X1 U1645 ( .IN1(n1864), .IN2(n1863), .IN3(n1862), .Q(n1931) );
  OR2X1 U1646 ( .IN1(\fpu_in_dp/n454 ), .IN2(n1856), .Q(n1949) );
  NOR4X0 U1647 ( .IN1(n121), .IN2(n1569), .IN3(n1568), .IN4(n1679), .QN(n1851)
         );
  AND2X1 U1648 ( .IN1(n1926), .IN2(n1848), .Q(n1893) );
  NAND3X0 U1649 ( .IN1(n1572), .IN2(n1570), .IN3(n1851), .QN(n1895) );
  AO22X1 U1650 ( .IN1(n1574), .IN2(n899), .IN3(n1580), .IN4(n897), .Q(n1855)
         );
  AO22X1 U1651 ( .IN1(n1578), .IN2(n895), .IN3(n1576), .IN4(n893), .Q(n1854)
         );
  AO22X1 U1652 ( .IN1(n1573), .IN2(n901), .IN3(n1575), .IN4(n903), .Q(n1853)
         );
  AO22X1 U1653 ( .IN1(n1579), .IN2(n907), .IN3(n1577), .IN4(n905), .Q(n1852)
         );
  OR4X1 U1654 ( .IN1(n1855), .IN2(n1854), .IN3(n1853), .IN4(n1852), .Q(n1865)
         );
  NOR3X0 U1655 ( .IN1(n1567), .IN2(\fpu_in_dp/n105 ), .IN3(n1895), .QN(n1937)
         );
  AO21X1 U1656 ( .IN1(\fpu_in_dp/n454 ), .IN2(n1938), .IN3(n1937), .Q(n1947)
         );
  MUX21X1 U1657 ( .IN1(n1671), .IN2(n1560), .S(n1651), .Q(n1860) );
  MUX21X1 U1658 ( .IN1(n1677), .IN2(n1562), .S(n1652), .Q(n1859) );
  MUX21X1 U1659 ( .IN1(n754), .IN2(n1675), .S(n755), .Q(n1858) );
  MUX21X1 U1660 ( .IN1(n1649), .IN2(n889), .S(n813), .Q(n1857) );
  NOR4X0 U1661 ( .IN1(n1860), .IN2(n1859), .IN3(n1858), .IN4(n1857), .QN(n1932) );
  NAND3X0 U1662 ( .IN1(n1932), .IN2(d1stg_step), .IN3(inq_wraddr[3]), .QN(
        n1867) );
  MUX21X1 U1663 ( .IN1(n807), .IN2(n1670), .S(n756), .Q(n1864) );
  MUX21X1 U1664 ( .IN1(n1650), .IN2(n886), .S(n1672), .Q(n1863) );
  AOI22X1 U1665 ( .IN1(n1565), .IN2(n1566), .IN3(n812), .IN4(n1564), .QN(n1861) );
  OA221X1 U1666 ( .IN1(n1565), .IN2(n1566), .IN3(n812), .IN4(n1564), .IN5(
        n1861), .Q(n1862) );
  MUX21X1 U1667 ( .IN1(n1865), .IN2(n1947), .S(n1905), .Q(inq_add) );
  NOR3X0 U1668 ( .IN1(n1866), .IN2(inq_add), .IN3(add_pipe_active), .QN(
        fadd_clken_l) );
  NOR4X0 U1669 ( .IN1(n418), .IN2(n890), .IN3(div_pipe_active), .IN4(inq_div), 
        .QN(fdiv_clken_l) );
  NOR3X0 U1670 ( .IN1(n1869), .IN2(inq_mul), .IN3(mul_pipe_active), .QN(
        fmul_clken_l) );
  NOR2X0 U1671 ( .IN1(fp_op_in_7in), .IN2(n1691), .QN(fp_src1_in[0]) );
  NOR2X0 U1672 ( .IN1(fp_op_in_7in), .IN2(n1646), .QN(fp_src1_in[10]) );
  NOR2X0 U1673 ( .IN1(fp_op_in_7in), .IN2(n1632), .QN(fp_src1_in[11]) );
  NOR2X0 U1674 ( .IN1(fp_op_in_7in), .IN2(n1666), .QN(fp_src1_in[12]) );
  NOR2X0 U1675 ( .IN1(fp_op_in_7in), .IN2(n1692), .QN(fp_src1_in[13]) );
  NOR2X0 U1676 ( .IN1(fp_op_in_7in), .IN2(n1647), .QN(fp_src1_in[14]) );
  NOR2X0 U1677 ( .IN1(fp_op_in_7in), .IN2(n1633), .QN(fp_src1_in[15]) );
  NOR2X0 U1678 ( .IN1(fp_op_in_7in), .IN2(n1667), .QN(fp_src1_in[16]) );
  NOR2X0 U1679 ( .IN1(fp_op_in_7in), .IN2(n1644), .QN(fp_src1_in[18]) );
  NOR2X0 U1680 ( .IN1(fp_op_in_7in), .IN2(n1630), .QN(fp_src1_in[19]) );
  NOR2X0 U1681 ( .IN1(fp_op_in_7in), .IN2(n1664), .QN(fp_src1_in[1]) );
  NOR2X0 U1682 ( .IN1(fp_op_in_7in), .IN2(n1690), .QN(fp_src1_in[20]) );
  NOR2X0 U1683 ( .IN1(fp_op_in_7in), .IN2(n1631), .QN(fp_src1_in[22]) );
  NOR2X0 U1684 ( .IN1(fp_op_in_7in), .IN2(n1665), .QN(fp_src1_in[23]) );
  NOR2X0 U1685 ( .IN1(fp_op_in_7in), .IN2(n1688), .QN(fp_src1_in[24]) );
  NOR2X0 U1686 ( .IN1(fp_op_in_7in), .IN2(n1662), .QN(fp_src1_in[30]) );
  NOR2X0 U1687 ( .IN1(fp_op_in_7in), .IN2(n1686), .QN(fp_src1_in[31]) );
  NOR2X0 U1688 ( .IN1(fp_op_in_7in), .IN2(n1685), .QN(fp_src1_in[32]) );
  NOR2X0 U1689 ( .IN1(fp_op_in_7in), .IN2(n1657), .QN(fp_src1_in[35]) );
  NOR2X0 U1690 ( .IN1(fp_op_in_7in), .IN2(n1625), .QN(fp_src1_in[37]) );
  NOR2X0 U1691 ( .IN1(fp_op_in_7in), .IN2(n1638), .QN(fp_src1_in[40]) );
  NOR2X0 U1692 ( .IN1(fp_op_in_7in), .IN2(n1681), .QN(fp_src1_in[44]) );
  NOR2X0 U1693 ( .IN1(fp_op_in_7in), .IN2(n1626), .QN(fp_src1_in[48]) );
  NOR2X0 U1694 ( .IN1(fp_op_in_7in), .IN2(n1674), .QN(fp_src1_in[51]) );
  NOR2X0 U1695 ( .IN1(fp_op_in_7in), .IN2(n1635), .QN(fp_src1_in[52]) );
  NOR2X0 U1696 ( .IN1(fp_op_in_7in), .IN2(n1653), .QN(fp_src1_in[53]) );
  NOR2X0 U1697 ( .IN1(fp_op_in_7in), .IN2(n1678), .QN(fp_src1_in[56]) );
  NOR2X0 U1698 ( .IN1(fp_op_in_7in), .IN2(n1654), .QN(fp_src1_in[57]) );
  NOR2X0 U1699 ( .IN1(fp_op_in_7in), .IN2(n1680), .QN(fp_src1_in[59]) );
  NOR2X0 U1700 ( .IN1(fp_op_in_7in), .IN2(n1636), .QN(fp_src1_in[60]) );
  NAND4X0 U1701 ( .IN1(n1683), .IN2(n1638), .IN3(n1624), .IN4(n1658), .QN(
        n1874) );
  NAND4X0 U1702 ( .IN1(n1684), .IN2(n1639), .IN3(n1625), .IN4(n1659), .QN(
        n1873) );
  NAND4X0 U1703 ( .IN1(n1685), .IN2(n1640), .IN3(n1626), .IN4(n1660), .QN(
        n1872) );
  NOR4X0 U1704 ( .IN1(n764), .IN2(n751), .IN3(n765), .IN4(n773), .QN(n1870) );
  NAND4X0 U1705 ( .IN1(n1870), .IN2(n1657), .IN3(n1637), .IN4(n1681), .QN(
        n1871) );
  NOR4X0 U1706 ( .IN1(n1874), .IN2(n1873), .IN3(n1872), .IN4(n1871), .QN(n1885) );
  NAND4X0 U1707 ( .IN1(n1693), .IN2(n1648), .IN3(n1634), .IN4(n1668), .QN(
        n1878) );
  NAND4X0 U1708 ( .IN1(n1686), .IN2(n1641), .IN3(n1627), .IN4(n1661), .QN(
        n1877) );
  NAND4X0 U1709 ( .IN1(n1687), .IN2(n1642), .IN3(n1628), .IN4(n1662), .QN(
        n1876) );
  NAND4X0 U1710 ( .IN1(n1688), .IN2(n1643), .IN3(n1629), .IN4(n1663), .QN(
        n1875) );
  NOR4X0 U1711 ( .IN1(n1878), .IN2(n1877), .IN3(n1876), .IN4(n1875), .QN(n1884) );
  NAND4X0 U1712 ( .IN1(n1689), .IN2(n1644), .IN3(n1630), .IN4(n1664), .QN(
        n1882) );
  NAND4X0 U1713 ( .IN1(n1690), .IN2(n1645), .IN3(n1631), .IN4(n1665), .QN(
        n1881) );
  NAND4X0 U1714 ( .IN1(n1691), .IN2(n1646), .IN3(n1632), .IN4(n1666), .QN(
        n1880) );
  NAND4X0 U1715 ( .IN1(n1692), .IN2(n1647), .IN3(n1633), .IN4(n1667), .QN(
        n1879) );
  NOR4X0 U1716 ( .IN1(n1882), .IN2(n1881), .IN3(n1880), .IN4(n1879), .QN(n1883) );
  NAND3X0 U1717 ( .IN1(n1885), .IN2(n1884), .IN3(n1883), .QN(n1901) );
  NOR2X0 U1718 ( .IN1(fp_op_in_7in), .IN2(n1693), .QN(fp_src1_in[6]) );
  NOR2X0 U1719 ( .IN1(fp_op_in_7in), .IN2(n1648), .QN(fp_src1_in[7]) );
  MUX21X1 U1720 ( .IN1(n883), .IN2(n802), .S(fp_op_in_7in), .Q(fp_src2_in[0])
         );
  MUX21X1 U1721 ( .IN1(n882), .IN2(n784), .S(n1844), .Q(fp_src2_in[10]) );
  MUX21X1 U1722 ( .IN1(n881), .IN2(n793), .S(fp_op_in_7in), .Q(fp_src2_in[11])
         );
  MUX21X1 U1723 ( .IN1(n880), .IN2(n801), .S(n1844), .Q(fp_src2_in[12]) );
  MUX21X1 U1724 ( .IN1(n879), .IN2(n783), .S(fp_op_in_7in), .Q(fp_src2_in[13])
         );
  MUX21X1 U1725 ( .IN1(n878), .IN2(n782), .S(n1844), .Q(fp_src2_in[14]) );
  MUX21X1 U1726 ( .IN1(n877), .IN2(n792), .S(n1844), .Q(fp_src2_in[15]) );
  MUX21X1 U1727 ( .IN1(n876), .IN2(n762), .S(n1844), .Q(fp_src2_in[16]) );
  MUX21X1 U1728 ( .IN1(n875), .IN2(n747), .S(fp_op_in_7in), .Q(fp_src2_in[17])
         );
  MUX21X1 U1729 ( .IN1(n874), .IN2(n741), .S(n1844), .Q(fp_src2_in[18]) );
  MUX21X1 U1730 ( .IN1(n873), .IN2(n737), .S(fp_op_in_7in), .Q(fp_src2_in[19])
         );
  MUX21X1 U1731 ( .IN1(n872), .IN2(n781), .S(n1844), .Q(fp_src2_in[1]) );
  MUX21X1 U1732 ( .IN1(n871), .IN2(n761), .S(n1844), .Q(fp_src2_in[20]) );
  MUX21X1 U1733 ( .IN1(n870), .IN2(n746), .S(fp_op_in_7in), .Q(fp_src2_in[21])
         );
  MUX21X1 U1734 ( .IN1(n869), .IN2(n740), .S(n1844), .Q(fp_src2_in[22]) );
  MUX21X1 U1735 ( .IN1(n868), .IN2(n736), .S(fp_op_in_7in), .Q(fp_src2_in[23])
         );
  MUX21X1 U1736 ( .IN1(n867), .IN2(n800), .S(fp_op_in_7in), .Q(fp_src2_in[24])
         );
  MUX21X1 U1737 ( .IN1(n866), .IN2(n780), .S(n1844), .Q(fp_src2_in[25]) );
  MUX21X1 U1738 ( .IN1(n865), .IN2(n779), .S(fp_op_in_7in), .Q(fp_src2_in[26])
         );
  MUX21X1 U1739 ( .IN1(n864), .IN2(n791), .S(n1844), .Q(fp_src2_in[27]) );
  MUX21X1 U1740 ( .IN1(n863), .IN2(n760), .S(fp_op_in_7in), .Q(fp_src2_in[28])
         );
  MUX21X1 U1741 ( .IN1(n862), .IN2(n745), .S(n1844), .Q(fp_src2_in[29]) );
  MUX21X1 U1742 ( .IN1(n861), .IN2(n778), .S(fp_op_in_7in), .Q(fp_src2_in[2])
         );
  MUX21X1 U1743 ( .IN1(n860), .IN2(n768), .S(n1844), .Q(fp_src2_in[30]) );
  MUX21X1 U1744 ( .IN1(n859), .IN2(n769), .S(fp_op_in_7in), .Q(fp_src2_in[31])
         );
  MUX21X1 U1745 ( .IN1(n858), .IN2(n799), .S(n1844), .Q(fp_src2_in[32]) );
  MUX21X1 U1746 ( .IN1(n857), .IN2(n777), .S(fp_op_in_7in), .Q(fp_src2_in[33])
         );
  MUX21X1 U1747 ( .IN1(n856), .IN2(n776), .S(n1844), .Q(fp_src2_in[34]) );
  MUX21X1 U1748 ( .IN1(n855), .IN2(n790), .S(fp_op_in_7in), .Q(fp_src2_in[35])
         );
  MUX21X1 U1749 ( .IN1(n854), .IN2(n798), .S(n1844), .Q(fp_src2_in[36]) );
  MUX21X1 U1750 ( .IN1(n853), .IN2(n775), .S(fp_op_in_7in), .Q(fp_src2_in[37])
         );
  MUX21X1 U1751 ( .IN1(n852), .IN2(n789), .S(n1844), .Q(fp_src2_in[38]) );
  MUX21X1 U1752 ( .IN1(n851), .IN2(n766), .S(fp_op_in_7in), .Q(fp_src2_in[39])
         );
  MUX21X1 U1753 ( .IN1(n850), .IN2(n788), .S(fp_op_in_7in), .Q(fp_src2_in[3])
         );
  MUX21X1 U1754 ( .IN1(n849), .IN2(n797), .S(fp_op_in_7in), .Q(fp_src2_in[40])
         );
  MUX21X1 U1755 ( .IN1(n848), .IN2(n774), .S(fp_op_in_7in), .Q(fp_src2_in[41])
         );
  MUX21X1 U1756 ( .IN1(n847), .IN2(n787), .S(fp_op_in_7in), .Q(fp_src2_in[42])
         );
  MUX21X1 U1757 ( .IN1(n846), .IN2(n750), .S(fp_op_in_7in), .Q(fp_src2_in[43])
         );
  MUX21X1 U1758 ( .IN1(n845), .IN2(n749), .S(fp_op_in_7in), .Q(fp_src2_in[44])
         );
  MUX21X1 U1759 ( .IN1(n844), .IN2(n764), .S(fp_op_in_7in), .Q(fp_src2_in[45])
         );
  MUX21X1 U1760 ( .IN1(n843), .IN2(n751), .S(fp_op_in_7in), .Q(fp_src2_in[46])
         );
  MUX21X1 U1761 ( .IN1(n842), .IN2(n765), .S(fp_op_in_7in), .Q(fp_src2_in[47])
         );
  MUX21X1 U1762 ( .IN1(n841), .IN2(n796), .S(fp_op_in_7in), .Q(fp_src2_in[48])
         );
  MUX21X1 U1763 ( .IN1(n840), .IN2(n786), .S(fp_op_in_7in), .Q(fp_src2_in[49])
         );
  MUX21X1 U1764 ( .IN1(n839), .IN2(n795), .S(fp_op_in_7in), .Q(fp_src2_in[4])
         );
  MUX21X1 U1765 ( .IN1(n838), .IN2(n773), .S(n1844), .Q(fp_src2_in[50]) );
  MUX21X1 U1766 ( .IN1(n837), .IN2(n758), .S(n1844), .Q(fp_src2_in[51]) );
  MUX21X1 U1767 ( .IN1(n836), .IN2(n738), .S(n1844), .Q(fp_src2_in[52]) );
  MUX21X1 U1768 ( .IN1(n835), .IN2(n743), .S(n1844), .Q(fp_src2_in[53]) );
  MUX21X1 U1769 ( .IN1(n834), .IN2(n759), .S(n1844), .Q(fp_src2_in[54]) );
  MUX21X1 U1770 ( .IN1(n833), .IN2(n742), .S(n1844), .Q(fp_src2_in[55]) );
  MUX21X1 U1771 ( .IN1(n832), .IN2(n748), .S(n1844), .Q(fp_src2_in[56]) );
  MUX21X1 U1772 ( .IN1(n831), .IN2(n739), .S(n1844), .Q(fp_src2_in[57]) );
  MUX21X1 U1773 ( .IN1(n830), .IN2(n744), .S(n1844), .Q(fp_src2_in[58]) );
  MUX21X1 U1774 ( .IN1(n829), .IN2(n735), .S(n1844), .Q(fp_src2_in[59]) );
  MUX21X1 U1775 ( .IN1(n828), .IN2(n772), .S(n1844), .Q(fp_src2_in[5]) );
  MUX21X1 U1776 ( .IN1(n827), .IN2(n757), .S(n1844), .Q(fp_src2_in[60]) );
  MUX21X1 U1777 ( .IN1(n826), .IN2(n767), .S(n1844), .Q(fp_src2_in[61]) );
  MUX21X1 U1778 ( .IN1(n825), .IN2(n763), .S(n1844), .Q(fp_src2_in[62]) );
  MUX21X1 U1779 ( .IN1(n824), .IN2(n803), .S(n1844), .Q(fp_src2_in[63]) );
  NAND4X0 U1780 ( .IN1(n1885), .IN2(n1674), .IN3(n1635), .IN4(n1653), .QN(
        n1902) );
  MUX21X1 U1781 ( .IN1(n823), .IN2(n1902), .S(n1844), .Q(fp_src2_in[64]) );
  MUX21X1 U1782 ( .IN1(n822), .IN2(n1901), .S(n1844), .Q(fp_src2_in[65]) );
  NAND4X0 U1783 ( .IN1(n1886), .IN2(n1674), .IN3(n1635), .IN4(n1653), .QN(
        n1900) );
  MUX21X1 U1784 ( .IN1(n821), .IN2(n1900), .S(n1844), .Q(fp_src2_in[66]) );
  MUX21X1 U1785 ( .IN1(n820), .IN2(n1899), .S(n1844), .Q(fp_src2_in[67]) );
  MUX21X1 U1786 ( .IN1(n819), .IN2(n1898), .S(n1844), .Q(fp_src2_in[68]) );
  MUX21X1 U1787 ( .IN1(n818), .IN2(n771), .S(n1844), .Q(fp_src2_in[6]) );
  MUX21X1 U1788 ( .IN1(n817), .IN2(n785), .S(n1844), .Q(fp_src2_in[7]) );
  MUX21X1 U1789 ( .IN1(n816), .IN2(n794), .S(n1844), .Q(fp_src2_in[8]) );
  MUX21X1 U1790 ( .IN1(n815), .IN2(n770), .S(n1844), .Q(fp_src2_in[9]) );
  AND2X1 U1791 ( .IN1(grst_l), .IN2(n1849), .Q(\fpu_in_ctl/dffrl_in_ctl/N4 )
         );
  MUX21X1 U1792 ( .IN1(n1891), .IN2(n1890), .S(n813), .Q(
        \fpu_in_ctl/i_inq_div_rdptr/N3 ) );
  AND3X1 U1793 ( .IN1(n813), .IN2(n755), .IN3(n1887), .Q(n1888) );
  AO22X1 U1795 ( .IN1(n1891), .IN2(n806), .IN3(n1890), .IN4(n891), .Q(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N10 ) );
  AO22X1 U1796 ( .IN1(n1891), .IN2(n917), .IN3(n1890), .IN4(n805), .Q(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N4 ) );
  AO22X1 U1797 ( .IN1(n1891), .IN2(n805), .IN3(n1890), .IN4(n885), .Q(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N5 ) );
  AO22X1 U1798 ( .IN1(n1891), .IN2(n885), .IN3(n1890), .IN4(n804), .Q(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N6 ) );
  AO22X1 U1799 ( .IN1(n1891), .IN2(n804), .IN3(n1890), .IN4(n884), .Q(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N7 ) );
  AO22X1 U1800 ( .IN1(n1891), .IN2(n884), .IN3(n1890), .IN4(n752), .Q(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N8 ) );
  AO22X1 U1801 ( .IN1(n1891), .IN2(n752), .IN3(n1890), .IN4(n806), .Q(
        \fpu_in_ctl/i_inq_div_rdptr_dec/N9 ) );
  AND2X1 U1802 ( .IN1(n805), .IN2(n1892), .Q(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N12 ) );
  AND2X1 U1803 ( .IN1(n885), .IN2(n1892), .Q(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N13 ) );
  AND2X1 U1804 ( .IN1(n804), .IN2(n1892), .Q(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N14 ) );
  AND2X1 U1805 ( .IN1(n884), .IN2(n1892), .Q(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N15 ) );
  AND2X1 U1806 ( .IN1(n752), .IN2(n1892), .Q(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N16 ) );
  AND2X1 U1807 ( .IN1(n806), .IN2(n1892), .Q(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N17 ) );
  AND2X1 U1808 ( .IN1(n891), .IN2(n1892), .Q(
        \fpu_in_ctl/i_inq_rdaddr_del_dec/N18 ) );
  AO22X1 U1809 ( .IN1(inq_add), .IN2(a1stg_step), .IN3(m1stg_step), .IN4(
        inq_mul), .Q(n1926) );
  AO22X1 U1810 ( .IN1(n908), .IN2(n1894), .IN3(n810), .IN4(n1893), .Q(
        \fpu_in_ctl/i_inq_rdptr_dec/N10 ) );
  MUX21X1 U1811 ( .IN1(n916), .IN2(n908), .S(n1926), .Q(n1988) );
  OA21X1 U1812 ( .IN1(n418), .IN2(n1988), .IN3(n1850), .Q(
        \fpu_in_ctl/i_inq_rdptr_dec/N3 ) );
  AO22X1 U1813 ( .IN1(n916), .IN2(n1893), .IN3(n1894), .IN4(n809), .Q(
        \fpu_in_ctl/i_inq_rdptr_dec/N4 ) );
  AO22X1 U1814 ( .IN1(n1894), .IN2(n888), .IN3(n1893), .IN4(n809), .Q(
        \fpu_in_ctl/i_inq_rdptr_dec/N5 ) );
  AO22X1 U1815 ( .IN1(n1894), .IN2(n808), .IN3(n1893), .IN4(n888), .Q(
        \fpu_in_ctl/i_inq_rdptr_dec/N6 ) );
  AO22X1 U1816 ( .IN1(n1894), .IN2(n887), .IN3(n1893), .IN4(n808), .Q(
        \fpu_in_ctl/i_inq_rdptr_dec/N7 ) );
  AO22X1 U1817 ( .IN1(n1894), .IN2(n753), .IN3(n1893), .IN4(n887), .Q(
        \fpu_in_ctl/i_inq_rdptr_dec/N8 ) );
  AO22X1 U1818 ( .IN1(n1894), .IN2(n810), .IN3(n1893), .IN4(n753), .Q(
        \fpu_in_ctl/i_inq_rdptr_dec/N9 ) );
  AND2X1 U1819 ( .IN1(fp_src1_in[28]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N100 ) );
  AND2X1 U1820 ( .IN1(fp_src1_in[29]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N101 ) );
  AND2X1 U1821 ( .IN1(fp_src1_in[30]), .IN2(n1850), .Q(
        \fpu_in_dp/i_inq_din_d1/N102 ) );
  AND2X1 U1822 ( .IN1(fp_src1_in[31]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N103 ) );
  AND2X1 U1823 ( .IN1(fp_src1_in[32]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N104 ) );
  AND2X1 U1824 ( .IN1(fp_src1_in[33]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N105 ) );
  AND2X1 U1825 ( .IN1(fp_src1_in[34]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N106 ) );
  AND2X1 U1826 ( .IN1(fp_src1_in[35]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N107 ) );
  AND2X1 U1827 ( .IN1(fp_src1_in[36]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N108 ) );
  AND2X1 U1828 ( .IN1(fp_src1_in[37]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N109 ) );
  AND2X1 U1829 ( .IN1(fp_src1_in[38]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N110 ) );
  AND2X1 U1830 ( .IN1(fp_src1_in[39]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N111 ) );
  AND2X1 U1831 ( .IN1(fp_src1_in[40]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N112 ) );
  AND2X1 U1832 ( .IN1(fp_src1_in[41]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N113 ) );
  AND2X1 U1833 ( .IN1(fp_src1_in[42]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N114 ) );
  AND2X1 U1834 ( .IN1(fp_src1_in[43]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N115 ) );
  AND2X1 U1835 ( .IN1(fp_src1_in[44]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N116 ) );
  AND2X1 U1836 ( .IN1(fp_src1_in[45]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N117 ) );
  AND2X1 U1837 ( .IN1(fp_src1_in[46]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N118 ) );
  AND2X1 U1838 ( .IN1(fp_src1_in[47]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N119 ) );
  AND2X1 U1839 ( .IN1(fp_src1_in[48]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N120 ) );
  AND2X1 U1840 ( .IN1(fp_src1_in[49]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N121 ) );
  AND2X1 U1841 ( .IN1(fp_src1_in[50]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N122 ) );
  AND2X1 U1842 ( .IN1(fp_src1_in[51]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N123 ) );
  AND2X1 U1843 ( .IN1(fp_src1_in[52]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N124 ) );
  AND2X1 U1844 ( .IN1(fp_src1_in[53]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N125 ) );
  AND2X1 U1845 ( .IN1(fp_src1_in[54]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N126 ) );
  AND2X1 U1846 ( .IN1(fp_src1_in[55]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N127 ) );
  AND2X1 U1847 ( .IN1(fp_src1_in[56]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N128 ) );
  AND2X1 U1848 ( .IN1(fp_src1_in[57]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N129 ) );
  AND2X1 U1849 ( .IN1(fp_src1_in[58]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N130 ) );
  AND2X1 U1850 ( .IN1(fp_src1_in[59]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N131 ) );
  AND2X1 U1851 ( .IN1(fp_src1_in[60]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N132 ) );
  AND2X1 U1852 ( .IN1(fp_src1_in[61]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N133 ) );
  AND2X1 U1853 ( .IN1(fp_src1_in[62]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N134 ) );
  AND2X1 U1854 ( .IN1(fp_src1_in[63]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N135 ) );
  AND2X1 U1855 ( .IN1(n1902), .IN2(\fpu_in_dp/n105 ), .Q(fp_src1_in[64]) );
  AND2X1 U1856 ( .IN1(fp_src1_in[64]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N136 ) );
  AND2X1 U1857 ( .IN1(n1900), .IN2(\fpu_in_dp/n105 ), .Q(fp_src1_in[66]) );
  AND2X1 U1858 ( .IN1(fp_src1_in[66]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N138 ) );
  AND2X1 U1859 ( .IN1(n1850), .IN2(fp_src1_in[67]), .Q(
        \fpu_in_dp/i_inq_din_d1/N139 ) );
  AND2X1 U1860 ( .IN1(n1850), .IN2(fp_src1_in[68]), .Q(
        \fpu_in_dp/i_inq_din_d1/N140 ) );
  AND2X1 U1861 ( .IN1(fp_src1_in[0]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N72 ) );
  AND2X1 U1862 ( .IN1(fp_src1_in[1]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N73 ) );
  AND2X1 U1863 ( .IN1(fp_src1_in[2]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N74 ) );
  AND2X1 U1864 ( .IN1(fp_src1_in[3]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N75 ) );
  AND2X1 U1865 ( .IN1(fp_src1_in[4]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N76 ) );
  AND2X1 U1866 ( .IN1(fp_src1_in[5]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N77 ) );
  AND2X1 U1867 ( .IN1(fp_src1_in[6]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N78 ) );
  AND2X1 U1868 ( .IN1(fp_src1_in[7]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N79 ) );
  AND2X1 U1869 ( .IN1(fp_src1_in[8]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N80 ) );
  AND2X1 U1870 ( .IN1(fp_src1_in[9]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N81 ) );
  AND2X1 U1871 ( .IN1(fp_src1_in[10]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N82 ) );
  AND2X1 U1872 ( .IN1(fp_src1_in[11]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N83 ) );
  AND2X1 U1873 ( .IN1(fp_src1_in[12]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N84 ) );
  AND2X1 U1874 ( .IN1(fp_src1_in[13]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N85 ) );
  AND2X1 U1875 ( .IN1(fp_src1_in[14]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N86 ) );
  AND2X1 U1876 ( .IN1(fp_src1_in[15]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N87 ) );
  AND2X1 U1877 ( .IN1(fp_src1_in[16]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N88 ) );
  AND2X1 U1878 ( .IN1(fp_src1_in[17]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N89 ) );
  AND2X1 U1879 ( .IN1(fp_src1_in[18]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N90 ) );
  AND2X1 U1880 ( .IN1(fp_src1_in[19]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N91 ) );
  AND2X1 U1881 ( .IN1(fp_src1_in[20]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N92 ) );
  AND2X1 U1882 ( .IN1(fp_src1_in[21]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N93 ) );
  AND2X1 U1883 ( .IN1(fp_src1_in[22]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N94 ) );
  AND2X1 U1884 ( .IN1(fp_src1_in[23]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N95 ) );
  AND2X1 U1885 ( .IN1(fp_src1_in[24]), .IN2(n1850), .Q(
        \fpu_in_dp/i_inq_din_d1/N96 ) );
  AND2X1 U1886 ( .IN1(fp_src1_in[25]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N97 ) );
  AND2X1 U1887 ( .IN1(fp_src1_in[26]), .IN2(n1849), .Q(
        \fpu_in_dp/i_inq_din_d1/N98 ) );
  AND2X1 U1888 ( .IN1(fp_src1_in[27]), .IN2(n1850), .Q(
        \fpu_in_dp/i_inq_din_d1/N99 ) );
  AO22X1 U1889 ( .IN1(n1622), .IN2(n819), .IN3(n1903), .IN4(n1898), .Q(
        \fpu_in_dp/n646 ) );
  AO22X1 U1890 ( .IN1(n1899), .IN2(n1903), .IN3(n820), .IN4(n1622), .Q(
        \fpu_in_dp/n647 ) );
  AO22X1 U1891 ( .IN1(n1622), .IN2(n821), .IN3(n1903), .IN4(n1900), .Q(
        \fpu_in_dp/n648 ) );
  AO22X1 U1892 ( .IN1(n1622), .IN2(n822), .IN3(n1903), .IN4(n1901), .Q(
        \fpu_in_dp/n649 ) );
  AO22X1 U1893 ( .IN1(n1622), .IN2(n823), .IN3(n1903), .IN4(n1902), .Q(
        \fpu_in_dp/n650 ) );
  AO22X1 U1894 ( .IN1(n803), .IN2(n1903), .IN3(n824), .IN4(n1622), .Q(
        \fpu_in_dp/n651 ) );
  AO22X1 U1895 ( .IN1(n763), .IN2(n1903), .IN3(n825), .IN4(n1622), .Q(
        \fpu_in_dp/n652 ) );
  AO22X1 U1896 ( .IN1(n767), .IN2(n1903), .IN3(n826), .IN4(n1622), .Q(
        \fpu_in_dp/n653 ) );
  AO22X1 U1897 ( .IN1(n757), .IN2(n1903), .IN3(n827), .IN4(n1622), .Q(
        \fpu_in_dp/n654 ) );
  AO22X1 U1898 ( .IN1(n735), .IN2(n1903), .IN3(n829), .IN4(n1622), .Q(
        \fpu_in_dp/n655 ) );
  AO22X1 U1899 ( .IN1(n744), .IN2(n1903), .IN3(n830), .IN4(n1622), .Q(
        \fpu_in_dp/n656 ) );
  AO22X1 U1900 ( .IN1(n739), .IN2(n1903), .IN3(n831), .IN4(n1622), .Q(
        \fpu_in_dp/n657 ) );
  AO22X1 U1901 ( .IN1(n748), .IN2(n1903), .IN3(n832), .IN4(n1622), .Q(
        \fpu_in_dp/n658 ) );
  AO22X1 U1902 ( .IN1(n742), .IN2(n1903), .IN3(n833), .IN4(n1622), .Q(
        \fpu_in_dp/n659 ) );
  AO22X1 U1903 ( .IN1(n759), .IN2(n1903), .IN3(n834), .IN4(n1622), .Q(
        \fpu_in_dp/n660 ) );
  AO22X1 U1904 ( .IN1(n743), .IN2(n1903), .IN3(n835), .IN4(n1622), .Q(
        \fpu_in_dp/n661 ) );
  AO22X1 U1905 ( .IN1(n738), .IN2(n1903), .IN3(n836), .IN4(n1622), .Q(
        \fpu_in_dp/n662 ) );
  AO22X1 U1906 ( .IN1(n758), .IN2(n1903), .IN3(n837), .IN4(n1622), .Q(
        \fpu_in_dp/n663 ) );
  AO22X1 U1907 ( .IN1(n773), .IN2(n1903), .IN3(n838), .IN4(n1622), .Q(
        \fpu_in_dp/n664 ) );
  AO22X1 U1908 ( .IN1(n786), .IN2(n1903), .IN3(n840), .IN4(n1622), .Q(
        \fpu_in_dp/n665 ) );
  AO22X1 U1909 ( .IN1(n796), .IN2(n1903), .IN3(n841), .IN4(n1622), .Q(
        \fpu_in_dp/n666 ) );
  AO22X1 U1910 ( .IN1(n765), .IN2(n1903), .IN3(n842), .IN4(n1622), .Q(
        \fpu_in_dp/n667 ) );
  AO22X1 U1911 ( .IN1(n751), .IN2(n1903), .IN3(n843), .IN4(n1622), .Q(
        \fpu_in_dp/n668 ) );
  AO22X1 U1912 ( .IN1(n764), .IN2(n1903), .IN3(n844), .IN4(n1622), .Q(
        \fpu_in_dp/n669 ) );
  AO22X1 U1913 ( .IN1(n749), .IN2(n1903), .IN3(n845), .IN4(n1622), .Q(
        \fpu_in_dp/n670 ) );
  AO22X1 U1914 ( .IN1(n750), .IN2(n1903), .IN3(n846), .IN4(n1622), .Q(
        \fpu_in_dp/n671 ) );
  AO22X1 U1915 ( .IN1(n787), .IN2(n1903), .IN3(n847), .IN4(n1622), .Q(
        \fpu_in_dp/n672 ) );
  AO22X1 U1916 ( .IN1(n774), .IN2(n1903), .IN3(n848), .IN4(n1622), .Q(
        \fpu_in_dp/n673 ) );
  AO22X1 U1917 ( .IN1(n797), .IN2(n1903), .IN3(n849), .IN4(n1622), .Q(
        \fpu_in_dp/n674 ) );
  AO22X1 U1918 ( .IN1(n766), .IN2(n1903), .IN3(n851), .IN4(n1622), .Q(
        \fpu_in_dp/n675 ) );
  AO22X1 U1919 ( .IN1(n789), .IN2(n1903), .IN3(n852), .IN4(n1622), .Q(
        \fpu_in_dp/n676 ) );
  AO22X1 U1920 ( .IN1(n775), .IN2(n1903), .IN3(n853), .IN4(n1622), .Q(
        \fpu_in_dp/n677 ) );
  AO22X1 U1921 ( .IN1(n798), .IN2(n1903), .IN3(n854), .IN4(n1622), .Q(
        \fpu_in_dp/n678 ) );
  AO22X1 U1922 ( .IN1(n790), .IN2(n1903), .IN3(n855), .IN4(n1622), .Q(
        \fpu_in_dp/n679 ) );
  AO22X1 U1923 ( .IN1(n776), .IN2(n1903), .IN3(n856), .IN4(n1622), .Q(
        \fpu_in_dp/n680 ) );
  AO22X1 U1924 ( .IN1(n777), .IN2(n1903), .IN3(n857), .IN4(n1622), .Q(
        \fpu_in_dp/n681 ) );
  AO22X1 U1925 ( .IN1(n799), .IN2(n1903), .IN3(n858), .IN4(n1622), .Q(
        \fpu_in_dp/n682 ) );
  AO22X1 U1926 ( .IN1(n769), .IN2(n1903), .IN3(n859), .IN4(n1622), .Q(
        \fpu_in_dp/n683 ) );
  AO22X1 U1927 ( .IN1(n768), .IN2(n1903), .IN3(n860), .IN4(n1622), .Q(
        \fpu_in_dp/n684 ) );
  AO22X1 U1928 ( .IN1(n745), .IN2(n1903), .IN3(n862), .IN4(n1622), .Q(
        \fpu_in_dp/n685 ) );
  AO22X1 U1929 ( .IN1(n760), .IN2(n1903), .IN3(n863), .IN4(n1622), .Q(
        \fpu_in_dp/n686 ) );
  AO22X1 U1930 ( .IN1(n791), .IN2(n1903), .IN3(n864), .IN4(n1622), .Q(
        \fpu_in_dp/n687 ) );
  AO22X1 U1931 ( .IN1(n779), .IN2(n1903), .IN3(n865), .IN4(n1622), .Q(
        \fpu_in_dp/n688 ) );
  AO22X1 U1932 ( .IN1(n780), .IN2(n1903), .IN3(n866), .IN4(n1622), .Q(
        \fpu_in_dp/n689 ) );
  AO22X1 U1933 ( .IN1(n800), .IN2(n1903), .IN3(n867), .IN4(n1622), .Q(
        \fpu_in_dp/n690 ) );
  AO22X1 U1934 ( .IN1(n736), .IN2(n1903), .IN3(n868), .IN4(n1622), .Q(
        \fpu_in_dp/n691 ) );
  AO22X1 U1935 ( .IN1(n740), .IN2(n1903), .IN3(n869), .IN4(n1622), .Q(
        \fpu_in_dp/n692 ) );
  AO22X1 U1936 ( .IN1(n746), .IN2(n1903), .IN3(n870), .IN4(n1622), .Q(
        \fpu_in_dp/n693 ) );
  AO22X1 U1937 ( .IN1(n761), .IN2(n1903), .IN3(n871), .IN4(n1622), .Q(
        \fpu_in_dp/n694 ) );
  AO22X1 U1938 ( .IN1(n737), .IN2(n1903), .IN3(n873), .IN4(n1622), .Q(
        \fpu_in_dp/n695 ) );
  AO22X1 U1939 ( .IN1(n741), .IN2(n1903), .IN3(n874), .IN4(n1622), .Q(
        \fpu_in_dp/n696 ) );
  AO22X1 U1940 ( .IN1(n747), .IN2(n1903), .IN3(n875), .IN4(n1622), .Q(
        \fpu_in_dp/n697 ) );
  AO22X1 U1941 ( .IN1(n762), .IN2(n1903), .IN3(n876), .IN4(n1622), .Q(
        \fpu_in_dp/n698 ) );
  AO22X1 U1942 ( .IN1(n792), .IN2(n1903), .IN3(n877), .IN4(n1622), .Q(
        \fpu_in_dp/n699 ) );
  AO22X1 U1943 ( .IN1(n782), .IN2(n1903), .IN3(n878), .IN4(n1622), .Q(
        \fpu_in_dp/n700 ) );
  AO22X1 U1944 ( .IN1(n783), .IN2(n1903), .IN3(n879), .IN4(n1622), .Q(
        \fpu_in_dp/n701 ) );
  AO22X1 U1945 ( .IN1(n801), .IN2(n1903), .IN3(n880), .IN4(n1622), .Q(
        \fpu_in_dp/n702 ) );
  AO22X1 U1946 ( .IN1(n793), .IN2(n1903), .IN3(n881), .IN4(n1622), .Q(
        \fpu_in_dp/n703 ) );
  AO22X1 U1947 ( .IN1(n784), .IN2(n1903), .IN3(n882), .IN4(n1622), .Q(
        \fpu_in_dp/n704 ) );
  AO22X1 U1948 ( .IN1(n770), .IN2(n1903), .IN3(n815), .IN4(n1622), .Q(
        \fpu_in_dp/n705 ) );
  AO22X1 U1949 ( .IN1(n794), .IN2(n1903), .IN3(n816), .IN4(n1622), .Q(
        \fpu_in_dp/n706 ) );
  AO22X1 U1950 ( .IN1(n785), .IN2(n1903), .IN3(n817), .IN4(n1622), .Q(
        \fpu_in_dp/n707 ) );
  AO22X1 U1951 ( .IN1(n771), .IN2(n1903), .IN3(n818), .IN4(n1622), .Q(
        \fpu_in_dp/n708 ) );
  AO22X1 U1952 ( .IN1(n772), .IN2(n1903), .IN3(n828), .IN4(n1622), .Q(
        \fpu_in_dp/n709 ) );
  AO22X1 U1953 ( .IN1(n795), .IN2(n1903), .IN3(n839), .IN4(n1622), .Q(
        \fpu_in_dp/n710 ) );
  AO22X1 U1954 ( .IN1(n788), .IN2(n1903), .IN3(n850), .IN4(n1622), .Q(
        \fpu_in_dp/n711 ) );
  AO22X1 U1955 ( .IN1(n778), .IN2(n1903), .IN3(n861), .IN4(n1622), .Q(
        \fpu_in_dp/n712 ) );
  AO22X1 U1956 ( .IN1(n781), .IN2(n1903), .IN3(n872), .IN4(n1622), .Q(
        \fpu_in_dp/n713 ) );
  AO22X1 U1957 ( .IN1(n802), .IN2(n1903), .IN3(n883), .IN4(n1622), .Q(
        \fpu_in_dp/n714 ) );
  AOI22X1 U1958 ( .IN1(n6), .IN2(n1547), .IN3(n111), .IN4(n1548), .QN(n1906)
         );
  OA221X1 U1959 ( .IN1(n6), .IN2(n1547), .IN3(n111), .IN4(n1548), .IN5(n1906), 
        .Q(n1910) );
  AOI22X1 U1960 ( .IN1(n1682), .IN2(n1545), .IN3(n4), .IN4(n1546), .QN(n1907)
         );
  OA221X1 U1961 ( .IN1(n1682), .IN2(n1545), .IN3(n4), .IN4(n1546), .IN5(n1907), 
        .Q(n1909) );
  NAND4X0 U1962 ( .IN1(n1544), .IN2(n1910), .IN3(n1909), .IN4(n1908), .QN(
        n1911) );
  INVX0 U1963 ( .INP(inq_dout[146]), .ZN(n1912) );
  OAI222X1 U1964 ( .IN1(n1935), .IN2(n1912), .IN3(n1697), .IN4(\fpu_in_dp/n18 ), .IN5(n1934), .IN6(\fpu_in_dp/n445 ), .QN(inq_fcc[0]) );
  INVX0 U1965 ( .INP(inq_dout[147]), .ZN(n1913) );
  OAI222X1 U1966 ( .IN1(n1913), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n443 ), .IN5(n1697), .IN6(\fpu_in_dp/n16 ), .QN(inq_fcc[1])
         );
  INVX0 U1967 ( .INP(inq_dout[150]), .ZN(n1914) );
  OAI222X1 U1968 ( .IN1(n1914), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n469 ), .IN5(n1697), .IN6(\fpu_in_dp/n10 ), .QN(inq_id[0])
         );
  INVX0 U1969 ( .INP(inq_dout[151]), .ZN(n1915) );
  OAI222X1 U1970 ( .IN1(n1915), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n467 ), .IN5(n1697), .IN6(\fpu_in_dp/n8 ), .QN(inq_id[1])
         );
  INVX0 U1971 ( .INP(inq_dout[152]), .ZN(n1916) );
  OAI222X1 U1972 ( .IN1(n1916), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n465 ), .IN5(n1697), .IN6(\fpu_in_dp/n6 ), .QN(inq_id[2])
         );
  INVX0 U1973 ( .INP(inq_dout[153]), .ZN(n1917) );
  OAI222X1 U1974 ( .IN1(n1917), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n463 ), .IN5(n1697), .IN6(\fpu_in_dp/n4 ), .QN(inq_id[3])
         );
  INVX0 U1975 ( .INP(inq_dout[154]), .ZN(n1918) );
  OAI222X1 U1976 ( .IN1(n1918), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n461 ), .IN5(n1697), .IN6(\fpu_in_dp/n2 ), .QN(inq_id[4])
         );
  AO222X1 U1977 ( .IN1(n1769), .IN2(n1845), .IN3(n1839), .IN4(inq_dout[69]), 
        .IN5(n1841), .IN6(fp_src1_in[0]), .Q(inq_in1[0]) );
  AO222X1 U1978 ( .IN1(n1770), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[79]), 
        .IN5(n1843), .IN6(fp_src1_in[10]), .Q(inq_in1[10]) );
  AO222X1 U1979 ( .IN1(n1771), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[80]), 
        .IN5(n1842), .IN6(fp_src1_in[11]), .Q(inq_in1[11]) );
  AO222X1 U1980 ( .IN1(n1772), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[81]), 
        .IN5(n1841), .IN6(fp_src1_in[12]), .Q(inq_in1[12]) );
  AO222X1 U1981 ( .IN1(n1773), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[82]), 
        .IN5(n1842), .IN6(fp_src1_in[13]), .Q(inq_in1[13]) );
  AO222X1 U1982 ( .IN1(n1774), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[83]), 
        .IN5(n1842), .IN6(fp_src1_in[14]), .Q(inq_in1[14]) );
  AO222X1 U1983 ( .IN1(n1775), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[84]), 
        .IN5(n1842), .IN6(fp_src1_in[15]), .Q(inq_in1[15]) );
  AO222X1 U1984 ( .IN1(n1776), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[85]), 
        .IN5(n1842), .IN6(fp_src1_in[16]), .Q(inq_in1[16]) );
  AO222X1 U1985 ( .IN1(n1777), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[86]), 
        .IN5(n1842), .IN6(fp_src1_in[17]), .Q(inq_in1[17]) );
  AO222X1 U1986 ( .IN1(n1778), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[87]), 
        .IN5(n1842), .IN6(fp_src1_in[18]), .Q(inq_in1[18]) );
  AO222X1 U1987 ( .IN1(n1779), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[88]), 
        .IN5(n1842), .IN6(fp_src1_in[19]), .Q(inq_in1[19]) );
  AO222X1 U1988 ( .IN1(n1780), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[70]), 
        .IN5(n1842), .IN6(fp_src1_in[1]), .Q(inq_in1[1]) );
  AO222X1 U1989 ( .IN1(n1781), .IN2(n1847), .IN3(n1838), .IN4(inq_dout[89]), 
        .IN5(n1842), .IN6(fp_src1_in[20]), .Q(inq_in1[20]) );
  AO222X1 U1990 ( .IN1(n1782), .IN2(n1845), .IN3(n1839), .IN4(inq_dout[90]), 
        .IN5(n1842), .IN6(fp_src1_in[21]), .Q(inq_in1[21]) );
  AO222X1 U1991 ( .IN1(n1783), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[91]), 
        .IN5(n1842), .IN6(fp_src1_in[22]), .Q(inq_in1[22]) );
  AO222X1 U1992 ( .IN1(n1784), .IN2(n1847), .IN3(n1838), .IN4(inq_dout[92]), 
        .IN5(n1843), .IN6(fp_src1_in[23]), .Q(inq_in1[23]) );
  AO222X1 U1993 ( .IN1(n1785), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[93]), 
        .IN5(n1842), .IN6(fp_src1_in[24]), .Q(inq_in1[24]) );
  AO222X1 U1994 ( .IN1(n1786), .IN2(n1846), .IN3(n1838), .IN4(inq_dout[94]), 
        .IN5(n1842), .IN6(fp_src1_in[25]), .Q(inq_in1[25]) );
  AO222X1 U1995 ( .IN1(n1787), .IN2(n1847), .IN3(n1839), .IN4(inq_dout[95]), 
        .IN5(n1842), .IN6(fp_src1_in[26]), .Q(inq_in1[26]) );
  AO222X1 U1996 ( .IN1(n1788), .IN2(n1845), .IN3(n1839), .IN4(inq_dout[96]), 
        .IN5(n1841), .IN6(fp_src1_in[27]), .Q(inq_in1[27]) );
  AO222X1 U1997 ( .IN1(n1789), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[97]), 
        .IN5(n1841), .IN6(fp_src1_in[28]), .Q(inq_in1[28]) );
  AO222X1 U1998 ( .IN1(n1790), .IN2(n1847), .IN3(n1839), .IN4(inq_dout[98]), 
        .IN5(n1842), .IN6(fp_src1_in[29]), .Q(inq_in1[29]) );
  AO222X1 U1999 ( .IN1(n1791), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[71]), 
        .IN5(n1841), .IN6(fp_src1_in[2]), .Q(inq_in1[2]) );
  AO222X1 U2000 ( .IN1(n1792), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[99]), 
        .IN5(n1843), .IN6(fp_src1_in[30]), .Q(inq_in1[30]) );
  AO222X1 U2001 ( .IN1(n1793), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[100]), 
        .IN5(n1842), .IN6(fp_src1_in[31]), .Q(inq_in1[31]) );
  AO222X1 U2002 ( .IN1(n1794), .IN2(n1846), .IN3(n1839), .IN4(inq_dout[101]), 
        .IN5(n1843), .IN6(fp_src1_in[32]), .Q(inq_in1[32]) );
  AO222X1 U2003 ( .IN1(n1795), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[102]), 
        .IN5(n1843), .IN6(fp_src1_in[33]), .Q(inq_in1[33]) );
  AO222X1 U2004 ( .IN1(n1796), .IN2(n1846), .IN3(n1838), .IN4(inq_dout[103]), 
        .IN5(n1842), .IN6(fp_src1_in[34]), .Q(inq_in1[34]) );
  AO222X1 U2005 ( .IN1(n1797), .IN2(n1846), .IN3(n1838), .IN4(inq_dout[104]), 
        .IN5(n1841), .IN6(fp_src1_in[35]), .Q(inq_in1[35]) );
  AO222X1 U2006 ( .IN1(n1798), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[105]), 
        .IN5(n1843), .IN6(fp_src1_in[36]), .Q(inq_in1[36]) );
  AO222X1 U2007 ( .IN1(n1799), .IN2(n1846), .IN3(n1839), .IN4(inq_dout[106]), 
        .IN5(n1842), .IN6(fp_src1_in[37]), .Q(inq_in1[37]) );
  AO222X1 U2008 ( .IN1(n1800), .IN2(n1846), .IN3(n1838), .IN4(inq_dout[107]), 
        .IN5(n1841), .IN6(fp_src1_in[38]), .Q(inq_in1[38]) );
  AO222X1 U2009 ( .IN1(n1801), .IN2(n1846), .IN3(n1839), .IN4(inq_dout[108]), 
        .IN5(n1843), .IN6(fp_src1_in[39]), .Q(inq_in1[39]) );
  AO222X1 U2010 ( .IN1(n1802), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[72]), 
        .IN5(n1842), .IN6(fp_src1_in[3]), .Q(inq_in1[3]) );
  AO222X1 U2011 ( .IN1(n1803), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[109]), 
        .IN5(n1842), .IN6(fp_src1_in[40]), .Q(inq_in1[40]) );
  AO222X1 U2012 ( .IN1(n1804), .IN2(n1846), .IN3(n1838), .IN4(inq_dout[110]), 
        .IN5(n1841), .IN6(fp_src1_in[41]), .Q(inq_in1[41]) );
  AO222X1 U2013 ( .IN1(n1805), .IN2(n1847), .IN3(n1838), .IN4(inq_dout[111]), 
        .IN5(n1842), .IN6(fp_src1_in[42]), .Q(inq_in1[42]) );
  AO222X1 U2014 ( .IN1(n1806), .IN2(n1847), .IN3(n1839), .IN4(inq_dout[112]), 
        .IN5(n1841), .IN6(fp_src1_in[43]), .Q(inq_in1[43]) );
  AO222X1 U2015 ( .IN1(n1807), .IN2(n1847), .IN3(n1839), .IN4(inq_dout[113]), 
        .IN5(n1841), .IN6(fp_src1_in[44]), .Q(inq_in1[44]) );
  AO222X1 U2016 ( .IN1(n1808), .IN2(n1847), .IN3(n1840), .IN4(inq_dout[114]), 
        .IN5(n1843), .IN6(fp_src1_in[45]), .Q(inq_in1[45]) );
  AO222X1 U2017 ( .IN1(n1809), .IN2(n1847), .IN3(n1839), .IN4(inq_dout[115]), 
        .IN5(n1842), .IN6(fp_src1_in[46]), .Q(inq_in1[46]) );
  AO222X1 U2018 ( .IN1(n1810), .IN2(n1847), .IN3(n1838), .IN4(inq_dout[116]), 
        .IN5(n1843), .IN6(fp_src1_in[47]), .Q(inq_in1[47]) );
  AO222X1 U2019 ( .IN1(n1811), .IN2(n1847), .IN3(n1838), .IN4(inq_dout[117]), 
        .IN5(n1841), .IN6(fp_src1_in[48]), .Q(inq_in1[48]) );
  AO222X1 U2020 ( .IN1(n1812), .IN2(n1847), .IN3(n1840), .IN4(inq_dout[118]), 
        .IN5(n1843), .IN6(fp_src1_in[49]), .Q(inq_in1[49]) );
  AO222X1 U2021 ( .IN1(n1813), .IN2(n1847), .IN3(n1840), .IN4(inq_dout[73]), 
        .IN5(n1842), .IN6(fp_src1_in[4]), .Q(inq_in1[4]) );
  AO222X1 U2022 ( .IN1(n1814), .IN2(n1847), .IN3(n1840), .IN4(inq_dout[119]), 
        .IN5(n1842), .IN6(fp_src1_in[50]), .Q(inq_in1[50]) );
  AO222X1 U2023 ( .IN1(n1815), .IN2(n1847), .IN3(n1839), .IN4(inq_dout[120]), 
        .IN5(n1842), .IN6(fp_src1_in[51]), .Q(inq_in1[51]) );
  AO222X1 U2024 ( .IN1(n1816), .IN2(n1847), .IN3(n1838), .IN4(inq_dout[121]), 
        .IN5(n1843), .IN6(fp_src1_in[52]), .Q(inq_in1[52]) );
  AO222X1 U2025 ( .IN1(n1817), .IN2(n1845), .IN3(n1839), .IN4(inq_dout[122]), 
        .IN5(n1841), .IN6(fp_src1_in[53]), .Q(inq_in1[53]) );
  AO222X1 U2026 ( .IN1(n1818), .IN2(n1845), .IN3(n1840), .IN4(inq_dout[123]), 
        .IN5(n1843), .IN6(fp_src1_in[54]), .Q(inq_in1[54]) );
  AO222X1 U2027 ( .IN1(n1819), .IN2(n1847), .IN3(n1840), .IN4(inq_dout[124]), 
        .IN5(n1842), .IN6(fp_src1_in[55]), .Q(inq_in1[55]) );
  AO222X1 U2028 ( .IN1(n1820), .IN2(n1846), .IN3(n1838), .IN4(inq_dout[125]), 
        .IN5(n1841), .IN6(fp_src1_in[56]), .Q(inq_in1[56]) );
  AO222X1 U2029 ( .IN1(n1821), .IN2(n1846), .IN3(n1838), .IN4(inq_dout[126]), 
        .IN5(n1842), .IN6(fp_src1_in[57]), .Q(inq_in1[57]) );
  AO222X1 U2030 ( .IN1(n1822), .IN2(n1845), .IN3(n1838), .IN4(inq_dout[127]), 
        .IN5(n1841), .IN6(fp_src1_in[58]), .Q(inq_in1[58]) );
  AO222X1 U2031 ( .IN1(n1823), .IN2(n1847), .IN3(n1840), .IN4(inq_dout[128]), 
        .IN5(n1843), .IN6(fp_src1_in[59]), .Q(inq_in1[59]) );
  AO222X1 U2032 ( .IN1(n1824), .IN2(n1846), .IN3(n1838), .IN4(inq_dout[74]), 
        .IN5(n1842), .IN6(fp_src1_in[5]), .Q(inq_in1[5]) );
  AO222X1 U2033 ( .IN1(n1825), .IN2(n1847), .IN3(n1839), .IN4(inq_dout[129]), 
        .IN5(n1843), .IN6(fp_src1_in[60]), .Q(inq_in1[60]) );
  AO222X1 U2034 ( .IN1(n1826), .IN2(n1845), .IN3(n1839), .IN4(inq_dout[130]), 
        .IN5(n1843), .IN6(fp_src1_in[61]), .Q(inq_in1[61]) );
  AO222X1 U2035 ( .IN1(n1827), .IN2(n1847), .IN3(n1840), .IN4(inq_dout[131]), 
        .IN5(n1841), .IN6(fp_src1_in[62]), .Q(inq_in1[62]) );
  AO222X1 U2036 ( .IN1(n1828), .IN2(n1846), .IN3(n1838), .IN4(inq_dout[132]), 
        .IN5(n1841), .IN6(fp_src1_in[63]), .Q(inq_in1[63]) );
  AO222X1 U2037 ( .IN1(n1829), .IN2(n1847), .IN3(n1838), .IN4(inq_dout[75]), 
        .IN5(n1841), .IN6(fp_src1_in[6]), .Q(inq_in1[6]) );
  AO222X1 U2038 ( .IN1(n1830), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[76]), 
        .IN5(n1841), .IN6(fp_src1_in[7]), .Q(inq_in1[7]) );
  AO222X1 U2039 ( .IN1(n1831), .IN2(n1846), .IN3(n1839), .IN4(inq_dout[77]), 
        .IN5(n1841), .IN6(fp_src1_in[8]), .Q(inq_in1[8]) );
  AO222X1 U2040 ( .IN1(n1832), .IN2(n1845), .IN3(n1840), .IN4(inq_dout[78]), 
        .IN5(n1841), .IN6(fp_src1_in[9]), .Q(inq_in1[9]) );
  AO222X1 U2041 ( .IN1(n1699), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[134]), 
        .IN5(n1841), .IN6(fp_src1_in[65]), .Q(inq_in1_50_0_neq_0) );
  AO222X1 U2042 ( .IN1(n1833), .IN2(n1847), .IN3(n1839), .IN4(inq_dout[135]), 
        .IN5(n1841), .IN6(fp_src1_in[66]), .Q(inq_in1_53_0_neq_0) );
  AO222X1 U2043 ( .IN1(n1834), .IN2(n1846), .IN3(n1840), .IN4(inq_dout[133]), 
        .IN5(n1841), .IN6(fp_src1_in[64]), .Q(inq_in1_53_32_neq_0) );
  AO222X1 U2044 ( .IN1(n1835), .IN2(n1847), .IN3(fp_src1_in[67]), .IN4(n1842), 
        .IN5(inq_dout[136]), .IN6(n1838), .Q(inq_in1_exp_eq_0) );
  AO222X1 U2045 ( .IN1(n1836), .IN2(n1845), .IN3(fp_src1_in[68]), .IN4(n1843), 
        .IN5(inq_dout[137]), .IN6(n1838), .Q(inq_in1_exp_neq_ffs) );
  AO222X1 U2046 ( .IN1(n1700), .IN2(n1846), .IN3(fp_src2_in[0]), .IN4(n1843), 
        .IN5(inq_dout[0]), .IN6(n1840), .Q(inq_in2[0]) );
  AO222X1 U2047 ( .IN1(n1701), .IN2(n1847), .IN3(fp_src2_in[10]), .IN4(n1842), 
        .IN5(inq_dout[10]), .IN6(n1840), .Q(inq_in2[10]) );
  AO222X1 U2048 ( .IN1(n1702), .IN2(n1845), .IN3(fp_src2_in[11]), .IN4(n1843), 
        .IN5(inq_dout[11]), .IN6(n1840), .Q(inq_in2[11]) );
  AO222X1 U2049 ( .IN1(n1703), .IN2(n1845), .IN3(fp_src2_in[12]), .IN4(n1842), 
        .IN5(inq_dout[12]), .IN6(n1840), .Q(inq_in2[12]) );
  AO222X1 U2050 ( .IN1(n1704), .IN2(n1846), .IN3(fp_src2_in[13]), .IN4(n1843), 
        .IN5(inq_dout[13]), .IN6(n1840), .Q(inq_in2[13]) );
  AO222X1 U2051 ( .IN1(n1705), .IN2(n1847), .IN3(fp_src2_in[14]), .IN4(n1841), 
        .IN5(inq_dout[14]), .IN6(n1840), .Q(inq_in2[14]) );
  AO222X1 U2052 ( .IN1(n1706), .IN2(n1847), .IN3(fp_src2_in[15]), .IN4(n1843), 
        .IN5(inq_dout[15]), .IN6(n1840), .Q(inq_in2[15]) );
  AO222X1 U2053 ( .IN1(n1707), .IN2(n1847), .IN3(fp_src2_in[16]), .IN4(n1842), 
        .IN5(inq_dout[16]), .IN6(n1840), .Q(inq_in2[16]) );
  AO222X1 U2054 ( .IN1(n1708), .IN2(n1846), .IN3(fp_src2_in[17]), .IN4(n1841), 
        .IN5(inq_dout[17]), .IN6(n1840), .Q(inq_in2[17]) );
  AO222X1 U2055 ( .IN1(n1709), .IN2(n1845), .IN3(fp_src2_in[18]), .IN4(n1842), 
        .IN5(inq_dout[18]), .IN6(n1840), .Q(inq_in2[18]) );
  AO222X1 U2056 ( .IN1(n1710), .IN2(n1846), .IN3(fp_src2_in[19]), .IN4(n1842), 
        .IN5(inq_dout[19]), .IN6(n1840), .Q(inq_in2[19]) );
  AO222X1 U2057 ( .IN1(n1711), .IN2(n1847), .IN3(fp_src2_in[1]), .IN4(n1842), 
        .IN5(inq_dout[1]), .IN6(n1840), .Q(inq_in2[1]) );
  AO222X1 U2058 ( .IN1(n1712), .IN2(n1845), .IN3(fp_src2_in[20]), .IN4(n1841), 
        .IN5(inq_dout[20]), .IN6(n1840), .Q(inq_in2[20]) );
  AO222X1 U2059 ( .IN1(n1713), .IN2(n1846), .IN3(fp_src2_in[21]), .IN4(n1841), 
        .IN5(inq_dout[21]), .IN6(n1839), .Q(inq_in2[21]) );
  AO222X1 U2060 ( .IN1(n1714), .IN2(n1847), .IN3(fp_src2_in[22]), .IN4(n1841), 
        .IN5(inq_dout[22]), .IN6(n1840), .Q(inq_in2[22]) );
  AO222X1 U2061 ( .IN1(n1715), .IN2(n1847), .IN3(fp_src2_in[23]), .IN4(n1843), 
        .IN5(inq_dout[23]), .IN6(n1838), .Q(inq_in2[23]) );
  AO222X1 U2062 ( .IN1(n1716), .IN2(n1845), .IN3(fp_src2_in[24]), .IN4(n1841), 
        .IN5(inq_dout[24]), .IN6(n1839), .Q(inq_in2[24]) );
  AO222X1 U2063 ( .IN1(n1717), .IN2(n1845), .IN3(fp_src2_in[25]), .IN4(n1841), 
        .IN5(inq_dout[25]), .IN6(n1840), .Q(inq_in2[25]) );
  AO222X1 U2064 ( .IN1(n1718), .IN2(n1845), .IN3(fp_src2_in[26]), .IN4(n1841), 
        .IN5(inq_dout[26]), .IN6(n1838), .Q(inq_in2[26]) );
  AO222X1 U2065 ( .IN1(n1719), .IN2(n1847), .IN3(fp_src2_in[27]), .IN4(n1842), 
        .IN5(inq_dout[27]), .IN6(n1839), .Q(inq_in2[27]) );
  AO222X1 U2066 ( .IN1(n1720), .IN2(n1845), .IN3(fp_src2_in[28]), .IN4(n1842), 
        .IN5(inq_dout[28]), .IN6(n1840), .Q(inq_in2[28]) );
  AO222X1 U2067 ( .IN1(n1721), .IN2(n1846), .IN3(fp_src2_in[29]), .IN4(n1843), 
        .IN5(inq_dout[29]), .IN6(n1838), .Q(inq_in2[29]) );
  AO222X1 U2068 ( .IN1(n1722), .IN2(n1847), .IN3(fp_src2_in[2]), .IN4(n1841), 
        .IN5(inq_dout[2]), .IN6(n1839), .Q(inq_in2[2]) );
  AO222X1 U2069 ( .IN1(n1723), .IN2(n1845), .IN3(fp_src2_in[30]), .IN4(n1843), 
        .IN5(inq_dout[30]), .IN6(n1840), .Q(inq_in2[30]) );
  AO222X1 U2070 ( .IN1(n1724), .IN2(n1847), .IN3(fp_src2_in[31]), .IN4(n1842), 
        .IN5(inq_dout[31]), .IN6(n1838), .Q(inq_in2[31]) );
  AO222X1 U2071 ( .IN1(n1725), .IN2(n1846), .IN3(fp_src2_in[32]), .IN4(n1841), 
        .IN5(inq_dout[32]), .IN6(n1839), .Q(inq_in2[32]) );
  AO222X1 U2072 ( .IN1(n1726), .IN2(n1845), .IN3(fp_src2_in[33]), .IN4(n1842), 
        .IN5(inq_dout[33]), .IN6(n1840), .Q(inq_in2[33]) );
  AO222X1 U2073 ( .IN1(n1727), .IN2(n1847), .IN3(fp_src2_in[34]), .IN4(n1843), 
        .IN5(inq_dout[34]), .IN6(n1839), .Q(inq_in2[34]) );
  AO222X1 U2074 ( .IN1(n1728), .IN2(n1845), .IN3(fp_src2_in[35]), .IN4(n1843), 
        .IN5(inq_dout[35]), .IN6(n1839), .Q(inq_in2[35]) );
  AO222X1 U2075 ( .IN1(n1729), .IN2(n1845), .IN3(fp_src2_in[36]), .IN4(n1841), 
        .IN5(inq_dout[36]), .IN6(n1838), .Q(inq_in2[36]) );
  AO222X1 U2076 ( .IN1(n1730), .IN2(n1846), .IN3(fp_src2_in[37]), .IN4(n1843), 
        .IN5(inq_dout[37]), .IN6(n1840), .Q(inq_in2[37]) );
  AO222X1 U2077 ( .IN1(n1731), .IN2(n1846), .IN3(fp_src2_in[38]), .IN4(n1841), 
        .IN5(inq_dout[38]), .IN6(n1840), .Q(inq_in2[38]) );
  AO222X1 U2078 ( .IN1(n1732), .IN2(n1847), .IN3(fp_src2_in[39]), .IN4(n1841), 
        .IN5(inq_dout[39]), .IN6(n1839), .Q(inq_in2[39]) );
  AO222X1 U2079 ( .IN1(n1733), .IN2(n1847), .IN3(fp_src2_in[3]), .IN4(n1842), 
        .IN5(inq_dout[3]), .IN6(n1838), .Q(inq_in2[3]) );
  AO222X1 U2080 ( .IN1(n1734), .IN2(n1846), .IN3(fp_src2_in[40]), .IN4(n1843), 
        .IN5(inq_dout[40]), .IN6(n1840), .Q(inq_in2[40]) );
  AO222X1 U2081 ( .IN1(n1735), .IN2(n1846), .IN3(fp_src2_in[41]), .IN4(n1843), 
        .IN5(inq_dout[41]), .IN6(n1838), .Q(inq_in2[41]) );
  AO222X1 U2082 ( .IN1(n1736), .IN2(n1846), .IN3(fp_src2_in[42]), .IN4(n1842), 
        .IN5(inq_dout[42]), .IN6(n1839), .Q(inq_in2[42]) );
  AO222X1 U2083 ( .IN1(n1737), .IN2(n1845), .IN3(fp_src2_in[43]), .IN4(n1841), 
        .IN5(inq_dout[43]), .IN6(n1840), .Q(inq_in2[43]) );
  AO222X1 U2084 ( .IN1(n1738), .IN2(n1846), .IN3(fp_src2_in[44]), .IN4(n1842), 
        .IN5(inq_dout[44]), .IN6(n1839), .Q(inq_in2[44]) );
  AO222X1 U2085 ( .IN1(n1739), .IN2(n1845), .IN3(fp_src2_in[45]), .IN4(n1841), 
        .IN5(inq_dout[45]), .IN6(n1839), .Q(inq_in2[45]) );
  AO222X1 U2086 ( .IN1(n1740), .IN2(n1847), .IN3(fp_src2_in[46]), .IN4(n1843), 
        .IN5(inq_dout[46]), .IN6(n1839), .Q(inq_in2[46]) );
  AO222X1 U2087 ( .IN1(n1741), .IN2(n1846), .IN3(fp_src2_in[47]), .IN4(n1843), 
        .IN5(inq_dout[47]), .IN6(n1839), .Q(inq_in2[47]) );
  AO222X1 U2088 ( .IN1(n1742), .IN2(n1846), .IN3(fp_src2_in[48]), .IN4(n1843), 
        .IN5(inq_dout[48]), .IN6(n1839), .Q(inq_in2[48]) );
  AO222X1 U2089 ( .IN1(n1743), .IN2(n1846), .IN3(fp_src2_in[49]), .IN4(n1843), 
        .IN5(inq_dout[49]), .IN6(n1839), .Q(inq_in2[49]) );
  AO222X1 U2090 ( .IN1(n1744), .IN2(n1847), .IN3(fp_src2_in[4]), .IN4(n1843), 
        .IN5(inq_dout[4]), .IN6(n1839), .Q(inq_in2[4]) );
  AO222X1 U2091 ( .IN1(n1745), .IN2(n1847), .IN3(fp_src2_in[50]), .IN4(n1843), 
        .IN5(inq_dout[50]), .IN6(n1839), .Q(inq_in2[50]) );
  AO222X1 U2092 ( .IN1(n1746), .IN2(n1847), .IN3(fp_src2_in[51]), .IN4(n1843), 
        .IN5(inq_dout[51]), .IN6(n1839), .Q(inq_in2[51]) );
  AO222X1 U2093 ( .IN1(n1747), .IN2(n1847), .IN3(fp_src2_in[52]), .IN4(n1841), 
        .IN5(inq_dout[52]), .IN6(n1839), .Q(inq_in2[52]) );
  AO222X1 U2094 ( .IN1(n1748), .IN2(n1845), .IN3(fp_src2_in[53]), .IN4(n1843), 
        .IN5(inq_dout[53]), .IN6(n1839), .Q(inq_in2[53]) );
  AO222X1 U2095 ( .IN1(n1749), .IN2(n1846), .IN3(fp_src2_in[54]), .IN4(n1843), 
        .IN5(inq_dout[54]), .IN6(n1839), .Q(inq_in2[54]) );
  AO222X1 U2096 ( .IN1(n1750), .IN2(n1847), .IN3(fp_src2_in[55]), .IN4(n1843), 
        .IN5(inq_dout[55]), .IN6(n1839), .Q(inq_in2[55]) );
  AO222X1 U2097 ( .IN1(n1751), .IN2(n1845), .IN3(fp_src2_in[56]), .IN4(n1843), 
        .IN5(inq_dout[56]), .IN6(n1839), .Q(inq_in2[56]) );
  AO222X1 U2098 ( .IN1(n1752), .IN2(n1846), .IN3(fp_src2_in[57]), .IN4(n1843), 
        .IN5(inq_dout[57]), .IN6(n1838), .Q(inq_in2[57]) );
  AO222X1 U2099 ( .IN1(n1753), .IN2(n1847), .IN3(fp_src2_in[58]), .IN4(n1843), 
        .IN5(inq_dout[58]), .IN6(n1840), .Q(inq_in2[58]) );
  AO222X1 U2100 ( .IN1(n1754), .IN2(n1846), .IN3(fp_src2_in[59]), .IN4(n1842), 
        .IN5(inq_dout[59]), .IN6(n1839), .Q(inq_in2[59]) );
  AO222X1 U2101 ( .IN1(n1755), .IN2(n1845), .IN3(fp_src2_in[5]), .IN4(n1843), 
        .IN5(inq_dout[5]), .IN6(n1839), .Q(inq_in2[5]) );
  AO222X1 U2102 ( .IN1(n1756), .IN2(n1845), .IN3(fp_src2_in[60]), .IN4(n1843), 
        .IN5(inq_dout[60]), .IN6(n1838), .Q(inq_in2[60]) );
  AO222X1 U2103 ( .IN1(n1757), .IN2(n1845), .IN3(fp_src2_in[61]), .IN4(n1841), 
        .IN5(inq_dout[61]), .IN6(n1840), .Q(inq_in2[61]) );
  AO222X1 U2104 ( .IN1(n1758), .IN2(n1846), .IN3(fp_src2_in[62]), .IN4(n1843), 
        .IN5(inq_dout[62]), .IN6(n1840), .Q(inq_in2[62]) );
  AO222X1 U2105 ( .IN1(n1759), .IN2(n1845), .IN3(fp_src2_in[63]), .IN4(n1843), 
        .IN5(inq_dout[63]), .IN6(n1839), .Q(inq_in2[63]) );
  AO222X1 U2106 ( .IN1(n1760), .IN2(n1846), .IN3(fp_src2_in[6]), .IN4(n1843), 
        .IN5(inq_dout[6]), .IN6(n1838), .Q(inq_in2[6]) );
  AO222X1 U2107 ( .IN1(n1761), .IN2(n1846), .IN3(fp_src2_in[7]), .IN4(n1842), 
        .IN5(inq_dout[7]), .IN6(n1840), .Q(inq_in2[7]) );
  AO222X1 U2108 ( .IN1(n1762), .IN2(n1847), .IN3(fp_src2_in[8]), .IN4(n1842), 
        .IN5(inq_dout[8]), .IN6(n1838), .Q(inq_in2[8]) );
  AO222X1 U2109 ( .IN1(n1763), .IN2(n1845), .IN3(fp_src2_in[9]), .IN4(n1841), 
        .IN5(inq_dout[9]), .IN6(n1839), .Q(inq_in2[9]) );
  AO222X1 U2110 ( .IN1(n1764), .IN2(n1845), .IN3(n1839), .IN4(inq_dout[65]), 
        .IN5(n1841), .IN6(fp_src2_in[65]), .Q(inq_in2_50_0_neq_0) );
  AO222X1 U2111 ( .IN1(n1765), .IN2(n1847), .IN3(n1839), .IN4(inq_dout[66]), 
        .IN5(n1841), .IN6(fp_src2_in[66]), .Q(inq_in2_53_0_neq_0) );
  AO222X1 U2112 ( .IN1(n1766), .IN2(n1845), .IN3(n1839), .IN4(inq_dout[64]), 
        .IN5(n1841), .IN6(fp_src2_in[64]), .Q(inq_in2_53_32_neq_0) );
  AO222X1 U2113 ( .IN1(n1767), .IN2(n1847), .IN3(fp_src2_in[67]), .IN4(n1843), 
        .IN5(inq_dout[67]), .IN6(n1838), .Q(inq_in2_exp_eq_0) );
  AO222X1 U2114 ( .IN1(n1768), .IN2(n1847), .IN3(n1838), .IN4(inq_dout[68]), 
        .IN5(n1841), .IN6(fp_src2_in[68]), .Q(inq_in2_exp_neq_ffs) );
  INVX0 U2115 ( .INP(inq_dout[138]), .ZN(n1919) );
  OAI222X1 U2116 ( .IN1(n1919), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n473 ), .IN5(n1697), .IN6(\fpu_in_dp/n32 ), .QN(inq_op[0])
         );
  INVX0 U2117 ( .INP(inq_dout[139]), .ZN(n1920) );
  OAI222X1 U2118 ( .IN1(n1920), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n458 ), .IN5(n1697), .IN6(\fpu_in_dp/n31 ), .QN(inq_op[1])
         );
  INVX0 U2119 ( .INP(inq_dout[140]), .ZN(n1921) );
  OAI222X1 U2120 ( .IN1(n1921), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n456 ), .IN5(n1697), .IN6(\fpu_in_dp/n29 ), .QN(inq_op[2])
         );
  INVX0 U2121 ( .INP(inq_dout[141]), .ZN(n1922) );
  OAI222X1 U2122 ( .IN1(n1922), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n454 ), .IN5(n1697), .IN6(\fpu_in_dp/n27 ), .QN(inq_op[3])
         );
  INVX0 U2123 ( .INP(inq_dout[142]), .ZN(n1923) );
  OAI222X1 U2124 ( .IN1(n1923), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n452 ), .IN5(n1697), .IN6(\fpu_in_dp/n25 ), .QN(inq_op[4])
         );
  INVX0 U2125 ( .INP(inq_dout[143]), .ZN(n1924) );
  OAI222X1 U2126 ( .IN1(n1924), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n450 ), .IN5(n1697), .IN6(\fpu_in_dp/n23 ), .QN(inq_op[5])
         );
  INVX0 U2127 ( .INP(inq_dout[144]), .ZN(n1925) );
  OAI222X1 U2128 ( .IN1(n1925), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n448 ), .IN5(n1697), .IN6(\fpu_in_dp/n21 ), .QN(inq_op[6])
         );
  AO222X1 U2129 ( .IN1(n1837), .IN2(n1845), .IN3(fp_op_in_7in), .IN4(n1842), 
        .IN5(inq_dout[145]), .IN6(n1838), .Q(inq_op[7]) );
  AO22X1 U2130 ( .IN1(n813), .IN2(n1930), .IN3(n257), .IN4(n1159), .Q(
        inq_rdaddr[0]) );
  AO22X1 U2131 ( .IN1(n755), .IN2(n1930), .IN3(n256), .IN4(n1159), .Q(
        inq_rdaddr[1]) );
  AO22X1 U2132 ( .IN1(n255), .IN2(n1159), .IN3(n1930), .IN4(n1671), .Q(
        inq_rdaddr[2]) );
  INVX0 U2133 ( .INP(inq_dout[148]), .ZN(n1933) );
  OAI222X1 U2134 ( .IN1(n1933), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n441 ), .IN5(n1697), .IN6(\fpu_in_dp/n14 ), .QN(
        inq_rnd_mode[0]) );
  INVX0 U2135 ( .INP(inq_dout[149]), .ZN(n1936) );
  OAI222X1 U2136 ( .IN1(n1936), .IN2(n1935), .IN3(n1934), .IN4(
        \fpu_in_dp/n439 ), .IN5(n1697), .IN6(\fpu_in_dp/n12 ), .QN(
        inq_rnd_mode[1]) );
  OR2X1 U2137 ( .IN1(n1938), .IN2(n1937), .Q(inq_we) );
  MUX21X1 U2138 ( .IN1(n1649), .IN2(n1670), .S(n1985), .Q(inq_wraddr[0]) );
  MUX21X1 U2139 ( .IN1(n754), .IN2(n1650), .S(n1985), .Q(inq_wraddr[1]) );
  MUX21X1 U2140 ( .IN1(n1651), .IN2(n1673), .S(n1985), .Q(inq_wraddr[2]) );
  OR2X1 U2141 ( .IN1(n1942), .IN2(n1967), .Q(n1963) );
  AND2X1 U2142 ( .IN1(n1966), .IN2(n1947), .Q(n1944) );
  AO22X1 U2143 ( .IN1(n899), .IN2(n1939), .IN3(n1967), .IN4(n1944), .Q(n322)
         );
  NOR3X0 U2144 ( .IN1(n1949), .IN2(n1961), .IN3(n1973), .QN(n1945) );
  AO22X1 U2145 ( .IN1(n898), .IN2(n1939), .IN3(n1967), .IN4(n1945), .Q(n323)
         );
  OR2X1 U2146 ( .IN1(n1942), .IN2(n1968), .Q(n1951) );
  AO22X1 U2147 ( .IN1(n907), .IN2(n1940), .IN3(n1944), .IN4(n1968), .Q(n325)
         );
  AO22X1 U2148 ( .IN1(n906), .IN2(n1940), .IN3(n1945), .IN4(n1968), .Q(n326)
         );
  OR2X1 U2149 ( .IN1(n1942), .IN2(n1969), .Q(n1953) );
  AO22X1 U2150 ( .IN1(n897), .IN2(n1941), .IN3(n1944), .IN4(n1969), .Q(n328)
         );
  AO22X1 U2151 ( .IN1(n896), .IN2(n1941), .IN3(n1945), .IN4(n1969), .Q(n329)
         );
  OR2X1 U2152 ( .IN1(n1942), .IN2(n1959), .Q(n1955) );
  AO22X1 U2153 ( .IN1(n905), .IN2(n1946), .IN3(n1944), .IN4(n1959), .Q(n331)
         );
  AO22X1 U2154 ( .IN1(n904), .IN2(n1946), .IN3(n1945), .IN4(n1959), .Q(n332)
         );
  NAND3X0 U2155 ( .IN1(n1961), .IN2(n1963), .IN3(n1962), .QN(n1950) );
  AND3X1 U2156 ( .IN1(n1972), .IN2(n1948), .IN3(n1947), .Q(n1957) );
  AO22X1 U2157 ( .IN1(n895), .IN2(n1950), .IN3(n1967), .IN4(n1957), .Q(n334)
         );
  AO22X1 U2158 ( .IN1(n894), .IN2(n1950), .IN3(n1967), .IN4(n1958), .Q(n335)
         );
  AO22X1 U2159 ( .IN1(n903), .IN2(n1952), .IN3(n1968), .IN4(n1957), .Q(n337)
         );
  AO22X1 U2160 ( .IN1(n902), .IN2(n1952), .IN3(n1968), .IN4(n1958), .Q(n338)
         );
  AO22X1 U2161 ( .IN1(n893), .IN2(n1954), .IN3(n1969), .IN4(n1957), .Q(n340)
         );
  AO22X1 U2162 ( .IN1(n892), .IN2(n1954), .IN3(n1969), .IN4(n1958), .Q(n341)
         );
  AO22X1 U2163 ( .IN1(n901), .IN2(n1960), .IN3(n1959), .IN4(n1957), .Q(n343)
         );
  AO22X1 U2164 ( .IN1(n900), .IN2(n1960), .IN3(n1959), .IN4(n1958), .Q(n344)
         );
  AO21X1 U2165 ( .IN1(n1972), .IN2(n1969), .IN3(n1968), .Q(n1971) );
  AO22X1 U2166 ( .IN1(n1848), .IN2(n1971), .IN3(n1970), .IN4(n1650), .Q(n348)
         );
  OA221X1 U2167 ( .IN1(n807), .IN2(n1973), .IN3(n1670), .IN4(n1972), .IN5(
        n1848), .Q(n349) );
  NAND3X0 U2168 ( .IN1(n1561), .IN2(inq_wraddr[3]), .IN3(n1848), .QN(n1974) );
  AO22X1 U2169 ( .IN1(n914), .IN2(n1848), .IN3(n1982), .IN4(n1975), .Q(n350)
         );
  AO22X1 U2170 ( .IN1(n912), .IN2(n1848), .IN3(n1982), .IN4(n1976), .Q(n353)
         );
  AO22X1 U2171 ( .IN1(n913), .IN2(n1848), .IN3(n1982), .IN4(n1978), .Q(n356)
         );
  AO21X1 U2172 ( .IN1(n1848), .IN2(n911), .IN3(n1983), .Q(n359) );
  NAND3X0 U2173 ( .IN1(inq_wraddr[3]), .IN2(n1848), .IN3(n1651), .QN(n1979) );
  AO22X1 U2174 ( .IN1(n1975), .IN2(n1977), .IN3(n1848), .IN4(n1695), .Q(n362)
         );
  AO22X1 U2175 ( .IN1(n1976), .IN2(n1977), .IN3(n1848), .IN4(n1669), .Q(n365)
         );
  AO22X1 U2176 ( .IN1(n1978), .IN2(n1977), .IN3(n1848), .IN4(n1696), .Q(n368)
         );
  AO21X1 U2177 ( .IN1(n1848), .IN2(n1557), .IN3(n1981), .Q(n371) );
  OA21X1 U2178 ( .IN1(n1985), .IN2(n1980), .IN3(n1848), .Q(n1984) );
  AO222X1 U2179 ( .IN1(n1652), .IN2(n1984), .IN3(n1652), .IN4(n1982), .IN5(
        n1981), .IN6(n1563), .Q(n374) );
  AO21X1 U2180 ( .IN1(n1984), .IN2(n1651), .IN3(n1983), .Q(n375) );
  OA221X1 U2181 ( .IN1(n754), .IN2(inq_wraddr[3]), .IN3(n754), .IN4(n1649), 
        .IN5(n1984), .Q(n376) );
  OA221X1 U2182 ( .IN1(n889), .IN2(n1985), .IN3(n1649), .IN4(inq_wraddr[3]), 
        .IN5(n1848), .Q(n377) );
  MUX21X1 U2183 ( .IN1(n891), .IN2(n917), .S(n1986), .Q(n1987) );
  INVX0 U2184 ( .INP(n1987), .ZN(n1161) );
endmodule

